* SPICE3 file created from 20bitCounter.ext - technology: sky130A
V1 VDD GND 1.8
V2 Vclk GND pulse(0V 1.8V clk_offset clk_risetime clk_falltime {clk_period/2} clk_period 0deg) 
V4 Vreset GND pwl(0.0us 1.8V, 0.090us 1.8V, 0.091us 0.0V, 0.100us 0.0V, 0.101us 1.8V)

.param clk_period=1us clk_offset={clk_period/2} clk_risetime=5ns clk_falltime={clk_risetime}
.func data_time(x) {clk_offset/2 + x*(clk_period/2)}

.tran 1us {32*clk_period}
.save Vclk Vreset 
.save sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_[15]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/Q
.lib ~/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D Q Q_N RESET_B VNB VPB
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPB a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VNB RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPB CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 Q_N a_1847_47# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_448_47# D VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VNB a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_761_289# a_543_47# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 Q a_1283_21# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# a_27_47# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPB a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPB a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_193_47# a_27_47# VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1283_21# RESET_B VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPB a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X25 VNB a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 Q_N a_1847_47# VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VNB CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_761_289# a_543_47# VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 a_651_413# RESET_B VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 Q a_1283_21# VPB VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
.ends


C0 Vreset sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.11fF
C1 Vreset sky130_fd_sc_hd__dfrbp_1_0[16]/D 1.55fF
C2 sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.12fF
C3 Vreset sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0.11fF
C4 sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.12fF
C5 Vreset sky130_fd_sc_hd__dfrbp_1_0[4]/D 1.45fF
C6 Vreset sky130_fd_sc_hd__dfrbp_1_0[11]/D 1.68fF
C7 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.08fF
C8 sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.12fF
C9 Vreset sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.11fF
C10 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.08fF
C11 sky130_fd_sc_hd__dfrbp_1_0[1]/D Vreset 1.15fF
C12 sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/D 0.12fF
C13 sky130_fd_sc_hd__dfrbp_1_0[1]/Q Vreset 0.11fF
C14 sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.12fF
C15 Vreset sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.11fF
C16 Vreset sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.11fF
C17 sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.12fF
C18 Vreset sky130_fd_sc_hd__dfrbp_1_0[18]/D 1.55fF
C19 sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.12fF
C20 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C21 Vreset sky130_fd_sc_hd__dfrbp_1_0[6]/D 1.55fF
C22 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.12fF
C23 Vreset sky130_fd_sc_hd__dfrbp_1_0[13]/D 1.51fF
C24 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C25 Vreset sky130_fd_sc_hd__dfrbp_1_0[19]/D 1.30fF
C26 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C27 Vreset sky130_fd_sc_hd__dfrbp_1_0[8]/D 1.55fF
C28 sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.08fF
C29 Vreset sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.11fF
C30 Vreset sky130_fd_sc_hd__dfrbp_1_0[12]/Q 0.11fF
C31 sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.12fF
C32 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.08fF
C33 Vreset sky130_fd_sc_hd__dfrbp_1_0[0]/D 1.04fF
C34 sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.12fF
C35 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.08fF
C36 sky130_fd_sc_hd__dfrbp_1_0[2]/Q Vreset 0.11fF
C37 Vreset sky130_fd_sc_hd__dfrbp_1_0[15]/D 1.68fF
C38 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.08fF
C39 Vreset sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.02fF
C40 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.08fF
C41 Vreset sky130_fd_sc_hd__dfrbp_1_0[3]/D 1.68fF
C42 Vreset sky130_fd_sc_hd__dfrbp_1_0[10]/D 1.55fF
C43 sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.12fF
C44 Vreset sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.11fF
C45 Vclk sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.04fF
C46 Vreset sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.11fF
C47 sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.12fF
C48 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.12fF
C49 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.08fF
C50 Vreset sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.11fF
C51 Vreset sky130_fd_sc_hd__dfrbp_1_0[17]/D 1.68fF
C52 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C53 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C54 Vreset sky130_fd_sc_hd__dfrbp_1_0[5]/D 1.68fF
C55 Vreset sky130_fd_sc_hd__dfrbp_1_0[12]/D 1.55fF
C56 sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.12fF
C57 Vreset sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.11fF
C58 sky130_fd_sc_hd__dfrbp_1_0[11]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.12fF
C59 Vreset sky130_fd_sc_hd__dfrbp_1_0[7]/D 1.68fF
C60 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.08fF
C61 Vreset sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.11fF
C62 Vreset sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.11fF
C63 sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.08fF
C64 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.08fF
C65 Vreset sky130_fd_sc_hd__dfrbp_1_0[14]/D 1.55fF
C66 sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.12fF
C67 Vreset sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.11fF
C68 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.12fF
C69 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.08fF
C70 Vreset sky130_fd_sc_hd__dfrbp_1_0[2]/D 1.45fF
C71 Vreset sky130_fd_sc_hd__dfrbp_1_0[9]/D 1.68fF
C72 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.08fF
C73 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.12fF
C74 Vreset sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.11fF
C75 Vreset sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.11fF
C76 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.08fF
R0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t4 350.253
R1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t5 189.586
R2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n1 97.205
R3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t2 89.119
R4 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n0 79.305
R5 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n2 66.705
R6 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t3 63.333
R7 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n3 41.041
R8 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_761_289.t1 31.979
R9 sky130_fd_sc_hd__dfrbp_1_0[0]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_639_47.t0 198.571
R10 sky130_fd_sc_hd__dfrbp_1_0[0]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_805_47.t1 60
R11 GND.n75 GND.t58 126.237
R12 GND.n154 GND.t110 126.237
R13 GND.n233 GND.t99 126.237
R14 GND.n312 GND.t105 126.237
R15 GND.n391 GND.t111 126.237
R16 GND.n470 GND.t45 126.237
R17 GND.n549 GND.t80 126.237
R18 GND.n628 GND.t181 126.237
R19 GND.n1519 GND.t17 126.237
R20 GND.n1440 GND.t78 126.237
R21 GND.n1361 GND.t124 126.237
R22 GND.n1282 GND.t75 126.237
R23 GND.n1203 GND.t66 126.237
R24 GND.n1124 GND.t51 126.237
R25 GND.n1045 GND.t1 126.237
R26 GND.n966 GND.t4 126.237
R27 GND.n887 GND.t197 126.237
R28 GND.n808 GND.t49 126.237
R29 GND.n729 GND.t40 126.237
R30 GND.n650 GND.t14 126.237
R31 GND.n38 GND.t141 100
R32 GND.n117 GND.t143 100
R33 GND.n196 GND.t145 100
R34 GND.n275 GND.t147 100
R35 GND.n354 GND.t149 100
R36 GND.n433 GND.t151 100
R37 GND.n512 GND.t153 100
R38 GND.n591 GND.t155 100
R39 GND.n1556 GND.t157 100
R40 GND.n1476 GND.t159 100
R41 GND.n1397 GND.t161 100
R42 GND.n1318 GND.t163 100
R43 GND.n1239 GND.t165 100
R44 GND.n1160 GND.t167 100
R45 GND.n1081 GND.t169 100
R46 GND.n1002 GND.t171 100
R47 GND.n923 GND.t173 100
R48 GND.n844 GND.t175 100
R49 GND.n765 GND.t177 100
R50 GND.n686 GND.t179 100
R51 GND.n52 GND.t142 72.857
R52 GND.n131 GND.t144 72.857
R53 GND.n210 GND.t146 72.857
R54 GND.n289 GND.t148 72.857
R55 GND.n368 GND.t150 72.857
R56 GND.n447 GND.t152 72.857
R57 GND.n526 GND.t154 72.857
R58 GND.n605 GND.t156 72.857
R59 GND.n1541 GND.t158 72.857
R60 GND.n1462 GND.t160 72.857
R61 GND.n1383 GND.t162 72.857
R62 GND.n1304 GND.t164 72.857
R63 GND.n1225 GND.t166 72.857
R64 GND.n1146 GND.t168 72.857
R65 GND.n1067 GND.t170 72.857
R66 GND.n988 GND.t172 72.857
R67 GND.n909 GND.t174 72.857
R68 GND.n830 GND.t176 72.857
R69 GND.n751 GND.t178 72.857
R70 GND.n672 GND.t180 72.857
R71 GND.n38 GND.t36 70
R72 GND.n117 GND.t123 70
R73 GND.n196 GND.t187 70
R74 GND.n275 GND.t95 70
R75 GND.n354 GND.t199 70
R76 GND.n433 GND.t112 70
R77 GND.n512 GND.t104 70
R78 GND.n591 GND.t72 70
R79 GND.n1556 GND.t82 70
R80 GND.n1476 GND.t41 70
R81 GND.n1397 GND.t115 70
R82 GND.n1318 GND.t35 70
R83 GND.n1239 GND.t198 70
R84 GND.n1160 GND.t97 70
R85 GND.n1081 GND.t34 70
R86 GND.n1002 GND.t20 70
R87 GND.n923 GND.t189 70
R88 GND.n844 GND.t39 70
R89 GND.n765 GND.t73 70
R90 GND.n686 GND.t46 70
R91 GND.n25 GND.t96 67.587
R92 GND.n104 GND.t107 67.587
R93 GND.n183 GND.t121 67.587
R94 GND.n262 GND.t84 67.587
R95 GND.n341 GND.t195 67.587
R96 GND.n420 GND.t85 67.587
R97 GND.n499 GND.t184 67.587
R98 GND.n578 GND.t23 67.587
R99 GND.n1490 GND.t10 67.587
R100 GND.n1411 GND.t83 67.587
R101 GND.n1332 GND.t136 67.587
R102 GND.n1253 GND.t5 67.587
R103 GND.n1174 GND.t7 67.587
R104 GND.n1095 GND.t16 67.587
R105 GND.n1016 GND.t25 67.587
R106 GND.n937 GND.t185 67.587
R107 GND.n858 GND.t43 67.587
R108 GND.n779 GND.t29 67.587
R109 GND.n700 GND.t192 67.587
R110 GND.t0 GND.n1572 67.587
R111 GND.n52 GND.t98 60.579
R112 GND.n131 GND.t113 60.579
R113 GND.n210 GND.t64 60.579
R114 GND.n289 GND.t118 60.579
R115 GND.n368 GND.t102 60.579
R116 GND.n447 GND.t18 60.579
R117 GND.n526 GND.t116 60.579
R118 GND.n605 GND.t9 60.579
R119 GND.n1541 GND.t69 60.579
R120 GND.n1462 GND.t129 60.579
R121 GND.n1383 GND.t131 60.579
R122 GND.n1304 GND.t94 60.579
R123 GND.n1225 GND.t57 60.579
R124 GND.n1146 GND.t15 60.579
R125 GND.n1067 GND.t81 60.579
R126 GND.n988 GND.t132 60.579
R127 GND.n909 GND.t193 60.579
R128 GND.n830 GND.t186 60.579
R129 GND.n751 GND.t21 60.579
R130 GND.n672 GND.t52 60.579
R131 GND.n16 GND.t24 57.142
R132 GND.n93 GND.t138 57.142
R133 GND.n172 GND.t109 57.142
R134 GND.n251 GND.t122 57.142
R135 GND.n330 GND.t91 57.142
R136 GND.n409 GND.t92 57.142
R137 GND.n488 GND.t127 57.142
R138 GND.n567 GND.t86 57.142
R139 GND.n0 GND.t126 57.142
R140 GND.n1500 GND.t63 57.142
R141 GND.n1421 GND.t120 57.142
R142 GND.n1342 GND.t26 57.142
R143 GND.n1263 GND.t42 57.142
R144 GND.n1184 GND.t77 57.142
R145 GND.n1105 GND.t2 57.142
R146 GND.n1026 GND.t135 57.142
R147 GND.n947 GND.t19 57.142
R148 GND.n868 GND.t47 57.142
R149 GND.n789 GND.t44 57.142
R150 GND.n710 GND.t194 57.142
R151 GND.n646 GND.n641 50.786
R152 GND.n646 GND.n645 50.667
R153 GND.n24 GND.n23 50.667
R154 GND.n28 GND.n27 50.667
R155 GND.n31 GND.n30 50.667
R156 GND.n34 GND.n33 50.667
R157 GND.n37 GND.n36 50.667
R158 GND.n42 GND.n41 50.667
R159 GND.n45 GND.n44 50.667
R160 GND.n48 GND.n47 50.667
R161 GND.n51 GND.n50 50.667
R162 GND.n56 GND.n55 50.667
R163 GND.n59 GND.n58 50.667
R164 GND.n62 GND.n61 50.667
R165 GND.n65 GND.n64 50.667
R166 GND.n68 GND.n67 50.667
R167 GND.n71 GND.n70 50.667
R168 GND.n74 GND.n73 50.667
R169 GND.n78 GND.n77 50.667
R170 GND.n81 GND.n80 50.667
R171 GND.n86 GND.n85 50.667
R172 GND.n89 GND.n88 50.667
R173 GND.n92 GND.n91 50.667
R174 GND.n97 GND.n96 50.667
R175 GND.n100 GND.n99 50.667
R176 GND.n103 GND.n102 50.667
R177 GND.n107 GND.n106 50.667
R178 GND.n110 GND.n109 50.667
R179 GND.n113 GND.n112 50.667
R180 GND.n116 GND.n115 50.667
R181 GND.n121 GND.n120 50.667
R182 GND.n124 GND.n123 50.667
R183 GND.n127 GND.n126 50.667
R184 GND.n130 GND.n129 50.667
R185 GND.n135 GND.n134 50.667
R186 GND.n138 GND.n137 50.667
R187 GND.n141 GND.n140 50.667
R188 GND.n144 GND.n143 50.667
R189 GND.n147 GND.n146 50.667
R190 GND.n150 GND.n149 50.667
R191 GND.n153 GND.n152 50.667
R192 GND.n157 GND.n156 50.667
R193 GND.n160 GND.n159 50.667
R194 GND.n165 GND.n164 50.667
R195 GND.n168 GND.n167 50.667
R196 GND.n171 GND.n170 50.667
R197 GND.n176 GND.n175 50.667
R198 GND.n179 GND.n178 50.667
R199 GND.n182 GND.n181 50.667
R200 GND.n186 GND.n185 50.667
R201 GND.n189 GND.n188 50.667
R202 GND.n192 GND.n191 50.667
R203 GND.n195 GND.n194 50.667
R204 GND.n200 GND.n199 50.667
R205 GND.n203 GND.n202 50.667
R206 GND.n206 GND.n205 50.667
R207 GND.n209 GND.n208 50.667
R208 GND.n214 GND.n213 50.667
R209 GND.n217 GND.n216 50.667
R210 GND.n220 GND.n219 50.667
R211 GND.n223 GND.n222 50.667
R212 GND.n226 GND.n225 50.667
R213 GND.n229 GND.n228 50.667
R214 GND.n232 GND.n231 50.667
R215 GND.n236 GND.n235 50.667
R216 GND.n239 GND.n238 50.667
R217 GND.n244 GND.n243 50.667
R218 GND.n247 GND.n246 50.667
R219 GND.n250 GND.n249 50.667
R220 GND.n255 GND.n254 50.667
R221 GND.n258 GND.n257 50.667
R222 GND.n261 GND.n260 50.667
R223 GND.n265 GND.n264 50.667
R224 GND.n268 GND.n267 50.667
R225 GND.n271 GND.n270 50.667
R226 GND.n274 GND.n273 50.667
R227 GND.n279 GND.n278 50.667
R228 GND.n282 GND.n281 50.667
R229 GND.n285 GND.n284 50.667
R230 GND.n288 GND.n287 50.667
R231 GND.n293 GND.n292 50.667
R232 GND.n296 GND.n295 50.667
R233 GND.n299 GND.n298 50.667
R234 GND.n302 GND.n301 50.667
R235 GND.n305 GND.n304 50.667
R236 GND.n308 GND.n307 50.667
R237 GND.n311 GND.n310 50.667
R238 GND.n315 GND.n314 50.667
R239 GND.n318 GND.n317 50.667
R240 GND.n323 GND.n322 50.667
R241 GND.n326 GND.n325 50.667
R242 GND.n329 GND.n328 50.667
R243 GND.n334 GND.n333 50.667
R244 GND.n337 GND.n336 50.667
R245 GND.n340 GND.n339 50.667
R246 GND.n344 GND.n343 50.667
R247 GND.n347 GND.n346 50.667
R248 GND.n350 GND.n349 50.667
R249 GND.n353 GND.n352 50.667
R250 GND.n358 GND.n357 50.667
R251 GND.n361 GND.n360 50.667
R252 GND.n364 GND.n363 50.667
R253 GND.n367 GND.n366 50.667
R254 GND.n372 GND.n371 50.667
R255 GND.n375 GND.n374 50.667
R256 GND.n378 GND.n377 50.667
R257 GND.n381 GND.n380 50.667
R258 GND.n384 GND.n383 50.667
R259 GND.n387 GND.n386 50.667
R260 GND.n390 GND.n389 50.667
R261 GND.n394 GND.n393 50.667
R262 GND.n397 GND.n396 50.667
R263 GND.n402 GND.n401 50.667
R264 GND.n405 GND.n404 50.667
R265 GND.n408 GND.n407 50.667
R266 GND.n413 GND.n412 50.667
R267 GND.n416 GND.n415 50.667
R268 GND.n419 GND.n418 50.667
R269 GND.n423 GND.n422 50.667
R270 GND.n426 GND.n425 50.667
R271 GND.n429 GND.n428 50.667
R272 GND.n432 GND.n431 50.667
R273 GND.n437 GND.n436 50.667
R274 GND.n440 GND.n439 50.667
R275 GND.n443 GND.n442 50.667
R276 GND.n446 GND.n445 50.667
R277 GND.n451 GND.n450 50.667
R278 GND.n454 GND.n453 50.667
R279 GND.n457 GND.n456 50.667
R280 GND.n460 GND.n459 50.667
R281 GND.n463 GND.n462 50.667
R282 GND.n466 GND.n465 50.667
R283 GND.n469 GND.n468 50.667
R284 GND.n473 GND.n472 50.667
R285 GND.n476 GND.n475 50.667
R286 GND.n481 GND.n480 50.667
R287 GND.n484 GND.n483 50.667
R288 GND.n487 GND.n486 50.667
R289 GND.n492 GND.n491 50.667
R290 GND.n495 GND.n494 50.667
R291 GND.n498 GND.n497 50.667
R292 GND.n502 GND.n501 50.667
R293 GND.n505 GND.n504 50.667
R294 GND.n508 GND.n507 50.667
R295 GND.n511 GND.n510 50.667
R296 GND.n516 GND.n515 50.667
R297 GND.n519 GND.n518 50.667
R298 GND.n522 GND.n521 50.667
R299 GND.n525 GND.n524 50.667
R300 GND.n530 GND.n529 50.667
R301 GND.n533 GND.n532 50.667
R302 GND.n536 GND.n535 50.667
R303 GND.n539 GND.n538 50.667
R304 GND.n542 GND.n541 50.667
R305 GND.n545 GND.n544 50.667
R306 GND.n548 GND.n547 50.667
R307 GND.n552 GND.n551 50.667
R308 GND.n555 GND.n554 50.667
R309 GND.n560 GND.n559 50.667
R310 GND.n563 GND.n562 50.667
R311 GND.n566 GND.n565 50.667
R312 GND.n571 GND.n570 50.667
R313 GND.n574 GND.n573 50.667
R314 GND.n577 GND.n576 50.667
R315 GND.n581 GND.n580 50.667
R316 GND.n584 GND.n583 50.667
R317 GND.n587 GND.n586 50.667
R318 GND.n590 GND.n589 50.667
R319 GND.n595 GND.n594 50.667
R320 GND.n598 GND.n597 50.667
R321 GND.n601 GND.n600 50.667
R322 GND.n604 GND.n603 50.667
R323 GND.n609 GND.n608 50.667
R324 GND.n612 GND.n611 50.667
R325 GND.n615 GND.n614 50.667
R326 GND.n618 GND.n617 50.667
R327 GND.n621 GND.n620 50.667
R328 GND.n624 GND.n623 50.667
R329 GND.n627 GND.n626 50.667
R330 GND.n631 GND.n630 50.667
R331 GND.n634 GND.n633 50.667
R332 GND.n1555 GND.n1553 50.667
R333 GND.n1545 GND.n1544 50.667
R334 GND.n1540 GND.n1539 50.667
R335 GND.n1537 GND.n1536 50.667
R336 GND.n1534 GND.n1533 50.667
R337 GND.n1531 GND.n1530 50.667
R338 GND.n1528 GND.n1527 50.667
R339 GND.n1525 GND.n1524 50.667
R340 GND.n1522 GND.n1521 50.667
R341 GND.n1518 GND.n1517 50.667
R342 GND.n1515 GND.n1514 50.667
R343 GND.n1510 GND.n1509 50.667
R344 GND.n1507 GND.n1506 50.667
R345 GND.n1504 GND.n1503 50.667
R346 GND.n1499 GND.n1498 50.667
R347 GND.n1496 GND.n1495 50.667
R348 GND.n1493 GND.n1492 50.667
R349 GND.n1489 GND.n1488 50.667
R350 GND.n1486 GND.n1485 50.667
R351 GND.n1483 GND.n1482 50.667
R352 GND.n1480 GND.n1479 50.667
R353 GND.n1475 GND.n1474 50.667
R354 GND.n1472 GND.n1471 50.667
R355 GND.n1469 GND.n1468 50.667
R356 GND.n1466 GND.n1465 50.667
R357 GND.n1461 GND.n1460 50.667
R358 GND.n1458 GND.n1457 50.667
R359 GND.n1455 GND.n1454 50.667
R360 GND.n1452 GND.n1451 50.667
R361 GND.n1449 GND.n1448 50.667
R362 GND.n1446 GND.n1445 50.667
R363 GND.n1443 GND.n1442 50.667
R364 GND.n1439 GND.n1438 50.667
R365 GND.n1436 GND.n1435 50.667
R366 GND.n1431 GND.n1430 50.667
R367 GND.n1428 GND.n1427 50.667
R368 GND.n1425 GND.n1424 50.667
R369 GND.n1420 GND.n1419 50.667
R370 GND.n1417 GND.n1416 50.667
R371 GND.n1414 GND.n1413 50.667
R372 GND.n1410 GND.n1409 50.667
R373 GND.n1407 GND.n1406 50.667
R374 GND.n1404 GND.n1403 50.667
R375 GND.n1401 GND.n1400 50.667
R376 GND.n1396 GND.n1395 50.667
R377 GND.n1393 GND.n1392 50.667
R378 GND.n1390 GND.n1389 50.667
R379 GND.n1387 GND.n1386 50.667
R380 GND.n1382 GND.n1381 50.667
R381 GND.n1379 GND.n1378 50.667
R382 GND.n1376 GND.n1375 50.667
R383 GND.n1373 GND.n1372 50.667
R384 GND.n1370 GND.n1369 50.667
R385 GND.n1367 GND.n1366 50.667
R386 GND.n1364 GND.n1363 50.667
R387 GND.n1360 GND.n1359 50.667
R388 GND.n1357 GND.n1356 50.667
R389 GND.n1352 GND.n1351 50.667
R390 GND.n1349 GND.n1348 50.667
R391 GND.n1346 GND.n1345 50.667
R392 GND.n1341 GND.n1340 50.667
R393 GND.n1338 GND.n1337 50.667
R394 GND.n1335 GND.n1334 50.667
R395 GND.n1331 GND.n1330 50.667
R396 GND.n1328 GND.n1327 50.667
R397 GND.n1325 GND.n1324 50.667
R398 GND.n1322 GND.n1321 50.667
R399 GND.n1317 GND.n1316 50.667
R400 GND.n1314 GND.n1313 50.667
R401 GND.n1311 GND.n1310 50.667
R402 GND.n1308 GND.n1307 50.667
R403 GND.n1303 GND.n1302 50.667
R404 GND.n1300 GND.n1299 50.667
R405 GND.n1297 GND.n1296 50.667
R406 GND.n1294 GND.n1293 50.667
R407 GND.n1291 GND.n1290 50.667
R408 GND.n1288 GND.n1287 50.667
R409 GND.n1285 GND.n1284 50.667
R410 GND.n1281 GND.n1280 50.667
R411 GND.n1278 GND.n1277 50.667
R412 GND.n1273 GND.n1272 50.667
R413 GND.n1270 GND.n1269 50.667
R414 GND.n1267 GND.n1266 50.667
R415 GND.n1262 GND.n1261 50.667
R416 GND.n1259 GND.n1258 50.667
R417 GND.n1256 GND.n1255 50.667
R418 GND.n1252 GND.n1251 50.667
R419 GND.n1249 GND.n1248 50.667
R420 GND.n1246 GND.n1245 50.667
R421 GND.n1243 GND.n1242 50.667
R422 GND.n1238 GND.n1237 50.667
R423 GND.n1235 GND.n1234 50.667
R424 GND.n1232 GND.n1231 50.667
R425 GND.n1229 GND.n1228 50.667
R426 GND.n1224 GND.n1223 50.667
R427 GND.n1221 GND.n1220 50.667
R428 GND.n1218 GND.n1217 50.667
R429 GND.n1215 GND.n1214 50.667
R430 GND.n1212 GND.n1211 50.667
R431 GND.n1209 GND.n1208 50.667
R432 GND.n1206 GND.n1205 50.667
R433 GND.n1202 GND.n1201 50.667
R434 GND.n1199 GND.n1198 50.667
R435 GND.n1194 GND.n1193 50.667
R436 GND.n1191 GND.n1190 50.667
R437 GND.n1188 GND.n1187 50.667
R438 GND.n1183 GND.n1182 50.667
R439 GND.n1180 GND.n1179 50.667
R440 GND.n1177 GND.n1176 50.667
R441 GND.n1173 GND.n1172 50.667
R442 GND.n1170 GND.n1169 50.667
R443 GND.n1167 GND.n1166 50.667
R444 GND.n1164 GND.n1163 50.667
R445 GND.n1159 GND.n1158 50.667
R446 GND.n1156 GND.n1155 50.667
R447 GND.n1153 GND.n1152 50.667
R448 GND.n1150 GND.n1149 50.667
R449 GND.n1145 GND.n1144 50.667
R450 GND.n1142 GND.n1141 50.667
R451 GND.n1139 GND.n1138 50.667
R452 GND.n1136 GND.n1135 50.667
R453 GND.n1133 GND.n1132 50.667
R454 GND.n1130 GND.n1129 50.667
R455 GND.n1127 GND.n1126 50.667
R456 GND.n1123 GND.n1122 50.667
R457 GND.n1120 GND.n1119 50.667
R458 GND.n1115 GND.n1114 50.667
R459 GND.n1112 GND.n1111 50.667
R460 GND.n1109 GND.n1108 50.667
R461 GND.n1104 GND.n1103 50.667
R462 GND.n1101 GND.n1100 50.667
R463 GND.n1098 GND.n1097 50.667
R464 GND.n1094 GND.n1093 50.667
R465 GND.n1091 GND.n1090 50.667
R466 GND.n1088 GND.n1087 50.667
R467 GND.n1085 GND.n1084 50.667
R468 GND.n1080 GND.n1079 50.667
R469 GND.n1077 GND.n1076 50.667
R470 GND.n1074 GND.n1073 50.667
R471 GND.n1071 GND.n1070 50.667
R472 GND.n1066 GND.n1065 50.667
R473 GND.n1063 GND.n1062 50.667
R474 GND.n1060 GND.n1059 50.667
R475 GND.n1057 GND.n1056 50.667
R476 GND.n1054 GND.n1053 50.667
R477 GND.n1051 GND.n1050 50.667
R478 GND.n1048 GND.n1047 50.667
R479 GND.n1044 GND.n1043 50.667
R480 GND.n1041 GND.n1040 50.667
R481 GND.n1036 GND.n1035 50.667
R482 GND.n1033 GND.n1032 50.667
R483 GND.n1030 GND.n1029 50.667
R484 GND.n1025 GND.n1024 50.667
R485 GND.n1022 GND.n1021 50.667
R486 GND.n1019 GND.n1018 50.667
R487 GND.n1015 GND.n1014 50.667
R488 GND.n1012 GND.n1011 50.667
R489 GND.n1009 GND.n1008 50.667
R490 GND.n1006 GND.n1005 50.667
R491 GND.n1001 GND.n1000 50.667
R492 GND.n998 GND.n997 50.667
R493 GND.n995 GND.n994 50.667
R494 GND.n992 GND.n991 50.667
R495 GND.n987 GND.n986 50.667
R496 GND.n984 GND.n983 50.667
R497 GND.n981 GND.n980 50.667
R498 GND.n978 GND.n977 50.667
R499 GND.n975 GND.n974 50.667
R500 GND.n972 GND.n971 50.667
R501 GND.n969 GND.n968 50.667
R502 GND.n965 GND.n964 50.667
R503 GND.n962 GND.n961 50.667
R504 GND.n957 GND.n956 50.667
R505 GND.n954 GND.n953 50.667
R506 GND.n951 GND.n950 50.667
R507 GND.n946 GND.n945 50.667
R508 GND.n943 GND.n942 50.667
R509 GND.n940 GND.n939 50.667
R510 GND.n936 GND.n935 50.667
R511 GND.n933 GND.n932 50.667
R512 GND.n930 GND.n929 50.667
R513 GND.n927 GND.n926 50.667
R514 GND.n922 GND.n921 50.667
R515 GND.n919 GND.n918 50.667
R516 GND.n916 GND.n915 50.667
R517 GND.n913 GND.n912 50.667
R518 GND.n908 GND.n907 50.667
R519 GND.n905 GND.n904 50.667
R520 GND.n902 GND.n901 50.667
R521 GND.n899 GND.n898 50.667
R522 GND.n896 GND.n895 50.667
R523 GND.n893 GND.n892 50.667
R524 GND.n890 GND.n889 50.667
R525 GND.n886 GND.n885 50.667
R526 GND.n883 GND.n882 50.667
R527 GND.n878 GND.n877 50.667
R528 GND.n875 GND.n874 50.667
R529 GND.n872 GND.n871 50.667
R530 GND.n867 GND.n866 50.667
R531 GND.n864 GND.n863 50.667
R532 GND.n861 GND.n860 50.667
R533 GND.n857 GND.n856 50.667
R534 GND.n854 GND.n853 50.667
R535 GND.n851 GND.n850 50.667
R536 GND.n848 GND.n847 50.667
R537 GND.n843 GND.n842 50.667
R538 GND.n840 GND.n839 50.667
R539 GND.n837 GND.n836 50.667
R540 GND.n834 GND.n833 50.667
R541 GND.n829 GND.n828 50.667
R542 GND.n826 GND.n825 50.667
R543 GND.n823 GND.n822 50.667
R544 GND.n820 GND.n819 50.667
R545 GND.n817 GND.n816 50.667
R546 GND.n814 GND.n813 50.667
R547 GND.n811 GND.n810 50.667
R548 GND.n807 GND.n806 50.667
R549 GND.n804 GND.n803 50.667
R550 GND.n799 GND.n798 50.667
R551 GND.n796 GND.n795 50.667
R552 GND.n793 GND.n792 50.667
R553 GND.n788 GND.n787 50.667
R554 GND.n785 GND.n784 50.667
R555 GND.n782 GND.n781 50.667
R556 GND.n778 GND.n777 50.667
R557 GND.n775 GND.n774 50.667
R558 GND.n772 GND.n771 50.667
R559 GND.n769 GND.n768 50.667
R560 GND.n764 GND.n763 50.667
R561 GND.n761 GND.n760 50.667
R562 GND.n758 GND.n757 50.667
R563 GND.n755 GND.n754 50.667
R564 GND.n750 GND.n749 50.667
R565 GND.n747 GND.n746 50.667
R566 GND.n744 GND.n743 50.667
R567 GND.n741 GND.n740 50.667
R568 GND.n738 GND.n737 50.667
R569 GND.n735 GND.n734 50.667
R570 GND.n732 GND.n731 50.667
R571 GND.n728 GND.n727 50.667
R572 GND.n725 GND.n724 50.667
R573 GND.n720 GND.n719 50.667
R574 GND.n717 GND.n716 50.667
R575 GND.n714 GND.n713 50.667
R576 GND.n709 GND.n708 50.667
R577 GND.n706 GND.n705 50.667
R578 GND.n703 GND.n702 50.667
R579 GND.n699 GND.n698 50.667
R580 GND.n696 GND.n695 50.667
R581 GND.n693 GND.n692 50.667
R582 GND.n690 GND.n689 50.667
R583 GND.n685 GND.n684 50.667
R584 GND.n682 GND.n681 50.667
R585 GND.n679 GND.n678 50.667
R586 GND.n676 GND.n675 50.667
R587 GND.n671 GND.n670 50.667
R588 GND.n668 GND.n667 50.667
R589 GND.n665 GND.n664 50.667
R590 GND.n662 GND.n661 50.667
R591 GND.n659 GND.n658 50.667
R592 GND.n656 GND.n655 50.667
R593 GND.n653 GND.n652 50.667
R594 GND.n649 GND.n648 50.667
R595 GND.n82 GND.t32 38.571
R596 GND.n82 GND.t100 38.571
R597 GND.n161 GND.t128 38.571
R598 GND.n161 GND.t68 38.571
R599 GND.n240 GND.t117 38.571
R600 GND.n240 GND.t134 38.571
R601 GND.n319 GND.t119 38.571
R602 GND.n319 GND.t133 38.571
R603 GND.n398 GND.t108 38.571
R604 GND.n398 GND.t60 38.571
R605 GND.n477 GND.t139 38.571
R606 GND.n477 GND.t88 38.571
R607 GND.n556 GND.t71 38.571
R608 GND.n556 GND.t190 38.571
R609 GND.n1 GND.t182 38.571
R610 GND.n1 GND.t28 38.571
R611 GND.n1511 GND.t125 38.571
R612 GND.n1511 GND.t79 38.571
R613 GND.n1432 GND.t59 38.571
R614 GND.n1432 GND.t183 38.571
R615 GND.n1353 GND.t74 38.571
R616 GND.n1353 GND.t76 38.571
R617 GND.n1274 GND.t137 38.571
R618 GND.n1274 GND.t87 38.571
R619 GND.n1195 GND.t114 38.571
R620 GND.n1195 GND.t53 38.571
R621 GND.n1116 GND.t90 38.571
R622 GND.n1116 GND.t3 38.571
R623 GND.n1037 GND.t27 38.571
R624 GND.n1037 GND.t196 38.571
R625 GND.n958 GND.t56 38.571
R626 GND.n958 GND.t55 38.571
R627 GND.n879 GND.t50 38.571
R628 GND.n879 GND.t12 38.571
R629 GND.n800 GND.t33 38.571
R630 GND.n800 GND.t11 38.571
R631 GND.n721 GND.t188 38.571
R632 GND.n721 GND.t37 38.571
R633 GND.n643 GND.t61 38.571
R634 GND.n643 GND.t103 38.571
R635 GND.n19 GND.n16 35.847
R636 GND.n94 GND.n93 35.847
R637 GND.n173 GND.n172 35.847
R638 GND.n252 GND.n251 35.847
R639 GND.n331 GND.n330 35.847
R640 GND.n410 GND.n409 35.847
R641 GND.n489 GND.n488 35.847
R642 GND.n568 GND.n567 35.847
R643 GND.n11 GND.n0 35.847
R644 GND.n1501 GND.n1500 35.847
R645 GND.n1422 GND.n1421 35.847
R646 GND.n1343 GND.n1342 35.847
R647 GND.n1264 GND.n1263 35.847
R648 GND.n1185 GND.n1184 35.847
R649 GND.n1106 GND.n1105 35.847
R650 GND.n1027 GND.n1026 35.847
R651 GND.n948 GND.n947 35.847
R652 GND.n869 GND.n868 35.847
R653 GND.n790 GND.n789 35.847
R654 GND.n711 GND.n710 35.847
R655 GND.n21 GND.n20 28.613
R656 GND.n16 GND.t130 25.428
R657 GND.n93 GND.t67 25.428
R658 GND.n172 GND.t89 25.428
R659 GND.n251 GND.t70 25.428
R660 GND.n330 GND.t106 25.428
R661 GND.n409 GND.t31 25.428
R662 GND.n488 GND.t65 25.428
R663 GND.n567 GND.t54 25.428
R664 GND.n0 GND.t93 25.428
R665 GND.n1500 GND.t101 25.428
R666 GND.n1421 GND.t38 25.428
R667 GND.n1342 GND.t22 25.428
R668 GND.n1263 GND.t8 25.428
R669 GND.n1184 GND.t140 25.428
R670 GND.n1105 GND.t6 25.428
R671 GND.n1026 GND.t62 25.428
R672 GND.n947 GND.t48 25.428
R673 GND.n868 GND.t13 25.428
R674 GND.n789 GND.t30 25.428
R675 GND.n710 GND.t191 25.428
R676 GND.n39 GND.n38 25.157
R677 GND.n118 GND.n117 25.157
R678 GND.n197 GND.n196 25.157
R679 GND.n276 GND.n275 25.157
R680 GND.n355 GND.n354 25.157
R681 GND.n434 GND.n433 25.157
R682 GND.n513 GND.n512 25.157
R683 GND.n592 GND.n591 25.157
R684 GND.n1565 GND.n1556 25.157
R685 GND.n1477 GND.n1476 25.157
R686 GND.n1398 GND.n1397 25.157
R687 GND.n1319 GND.n1318 25.157
R688 GND.n1240 GND.n1239 25.157
R689 GND.n1161 GND.n1160 25.157
R690 GND.n1082 GND.n1081 25.157
R691 GND.n1003 GND.n1002 25.157
R692 GND.n924 GND.n923 25.157
R693 GND.n845 GND.n844 25.157
R694 GND.n766 GND.n765 25.157
R695 GND.n687 GND.n686 25.157
R696 GND.n53 GND.n52 18.406
R697 GND.n83 GND.n82 18.406
R698 GND.n132 GND.n131 18.406
R699 GND.n162 GND.n161 18.406
R700 GND.n211 GND.n210 18.406
R701 GND.n241 GND.n240 18.406
R702 GND.n290 GND.n289 18.406
R703 GND.n320 GND.n319 18.406
R704 GND.n369 GND.n368 18.406
R705 GND.n399 GND.n398 18.406
R706 GND.n448 GND.n447 18.406
R707 GND.n478 GND.n477 18.406
R708 GND.n527 GND.n526 18.406
R709 GND.n557 GND.n556 18.406
R710 GND.n606 GND.n605 18.406
R711 GND.n4 GND.n1 18.406
R712 GND.n1542 GND.n1541 18.406
R713 GND.n1512 GND.n1511 18.406
R714 GND.n1463 GND.n1462 18.406
R715 GND.n1433 GND.n1432 18.406
R716 GND.n1384 GND.n1383 18.406
R717 GND.n1354 GND.n1353 18.406
R718 GND.n1305 GND.n1304 18.406
R719 GND.n1275 GND.n1274 18.406
R720 GND.n1226 GND.n1225 18.406
R721 GND.n1196 GND.n1195 18.406
R722 GND.n1147 GND.n1146 18.406
R723 GND.n1117 GND.n1116 18.406
R724 GND.n1068 GND.n1067 18.406
R725 GND.n1038 GND.n1037 18.406
R726 GND.n989 GND.n988 18.406
R727 GND.n959 GND.n958 18.406
R728 GND.n910 GND.n909 18.406
R729 GND.n880 GND.n879 18.406
R730 GND.n831 GND.n830 18.406
R731 GND.n801 GND.n800 18.406
R732 GND.n752 GND.n751 18.406
R733 GND.n722 GND.n721 18.406
R734 GND.n673 GND.n672 18.406
R735 GND.n644 GND.n643 18.406
R736 GND.n8 GND.n6 15.167
R737 GND.n10 GND.n8 15.167
R738 GND.n15 GND.n13 15.167
R739 GND.n1555 GND.n15 15.167
R740 GND.n1571 GND.n1569 15.167
R741 GND.n1569 GND.n1567 15.167
R742 GND.n1564 GND.n1562 15.167
R743 GND.n1562 GND.n1560 15.167
R744 GND.n1560 GND.n1558 15.167
R745 GND.n6 GND.n4 14.837
R746 GND.n19 GND.n18 13.683
R747 GND.n13 GND.n11 13.683
R748 GND.n1572 GND.n1571 12.2
R749 GND.n1567 GND.n1565 10.881
R750 GND.n645 GND.n642 7.147
R751 GND.n18 GND.n17 7.147
R752 GND.n23 GND.n22 7.147
R753 GND.n27 GND.n26 7.147
R754 GND.n30 GND.n29 7.147
R755 GND.n33 GND.n32 7.147
R756 GND.n36 GND.n35 7.147
R757 GND.n41 GND.n40 7.147
R758 GND.n44 GND.n43 7.147
R759 GND.n47 GND.n46 7.147
R760 GND.n50 GND.n49 7.147
R761 GND.n55 GND.n54 7.147
R762 GND.n58 GND.n57 7.147
R763 GND.n61 GND.n60 7.147
R764 GND.n64 GND.n63 7.147
R765 GND.n67 GND.n66 7.147
R766 GND.n70 GND.n69 7.147
R767 GND.n73 GND.n72 7.147
R768 GND.n77 GND.n76 7.147
R769 GND.n80 GND.n79 7.147
R770 GND.n85 GND.n84 7.147
R771 GND.n88 GND.n87 7.147
R772 GND.n91 GND.n90 7.147
R773 GND.n96 GND.n95 7.147
R774 GND.n99 GND.n98 7.147
R775 GND.n102 GND.n101 7.147
R776 GND.n106 GND.n105 7.147
R777 GND.n109 GND.n108 7.147
R778 GND.n112 GND.n111 7.147
R779 GND.n115 GND.n114 7.147
R780 GND.n120 GND.n119 7.147
R781 GND.n123 GND.n122 7.147
R782 GND.n126 GND.n125 7.147
R783 GND.n129 GND.n128 7.147
R784 GND.n134 GND.n133 7.147
R785 GND.n137 GND.n136 7.147
R786 GND.n140 GND.n139 7.147
R787 GND.n143 GND.n142 7.147
R788 GND.n146 GND.n145 7.147
R789 GND.n149 GND.n148 7.147
R790 GND.n152 GND.n151 7.147
R791 GND.n156 GND.n155 7.147
R792 GND.n159 GND.n158 7.147
R793 GND.n164 GND.n163 7.147
R794 GND.n167 GND.n166 7.147
R795 GND.n170 GND.n169 7.147
R796 GND.n175 GND.n174 7.147
R797 GND.n178 GND.n177 7.147
R798 GND.n181 GND.n180 7.147
R799 GND.n185 GND.n184 7.147
R800 GND.n188 GND.n187 7.147
R801 GND.n191 GND.n190 7.147
R802 GND.n194 GND.n193 7.147
R803 GND.n199 GND.n198 7.147
R804 GND.n202 GND.n201 7.147
R805 GND.n205 GND.n204 7.147
R806 GND.n208 GND.n207 7.147
R807 GND.n213 GND.n212 7.147
R808 GND.n216 GND.n215 7.147
R809 GND.n219 GND.n218 7.147
R810 GND.n222 GND.n221 7.147
R811 GND.n225 GND.n224 7.147
R812 GND.n228 GND.n227 7.147
R813 GND.n231 GND.n230 7.147
R814 GND.n235 GND.n234 7.147
R815 GND.n238 GND.n237 7.147
R816 GND.n243 GND.n242 7.147
R817 GND.n246 GND.n245 7.147
R818 GND.n249 GND.n248 7.147
R819 GND.n254 GND.n253 7.147
R820 GND.n257 GND.n256 7.147
R821 GND.n260 GND.n259 7.147
R822 GND.n264 GND.n263 7.147
R823 GND.n267 GND.n266 7.147
R824 GND.n270 GND.n269 7.147
R825 GND.n273 GND.n272 7.147
R826 GND.n278 GND.n277 7.147
R827 GND.n281 GND.n280 7.147
R828 GND.n284 GND.n283 7.147
R829 GND.n287 GND.n286 7.147
R830 GND.n292 GND.n291 7.147
R831 GND.n295 GND.n294 7.147
R832 GND.n298 GND.n297 7.147
R833 GND.n301 GND.n300 7.147
R834 GND.n304 GND.n303 7.147
R835 GND.n307 GND.n306 7.147
R836 GND.n310 GND.n309 7.147
R837 GND.n314 GND.n313 7.147
R838 GND.n317 GND.n316 7.147
R839 GND.n322 GND.n321 7.147
R840 GND.n325 GND.n324 7.147
R841 GND.n328 GND.n327 7.147
R842 GND.n333 GND.n332 7.147
R843 GND.n336 GND.n335 7.147
R844 GND.n339 GND.n338 7.147
R845 GND.n343 GND.n342 7.147
R846 GND.n346 GND.n345 7.147
R847 GND.n349 GND.n348 7.147
R848 GND.n352 GND.n351 7.147
R849 GND.n357 GND.n356 7.147
R850 GND.n360 GND.n359 7.147
R851 GND.n363 GND.n362 7.147
R852 GND.n366 GND.n365 7.147
R853 GND.n371 GND.n370 7.147
R854 GND.n374 GND.n373 7.147
R855 GND.n377 GND.n376 7.147
R856 GND.n380 GND.n379 7.147
R857 GND.n383 GND.n382 7.147
R858 GND.n386 GND.n385 7.147
R859 GND.n389 GND.n388 7.147
R860 GND.n393 GND.n392 7.147
R861 GND.n396 GND.n395 7.147
R862 GND.n401 GND.n400 7.147
R863 GND.n404 GND.n403 7.147
R864 GND.n407 GND.n406 7.147
R865 GND.n412 GND.n411 7.147
R866 GND.n415 GND.n414 7.147
R867 GND.n418 GND.n417 7.147
R868 GND.n422 GND.n421 7.147
R869 GND.n425 GND.n424 7.147
R870 GND.n428 GND.n427 7.147
R871 GND.n431 GND.n430 7.147
R872 GND.n436 GND.n435 7.147
R873 GND.n439 GND.n438 7.147
R874 GND.n442 GND.n441 7.147
R875 GND.n445 GND.n444 7.147
R876 GND.n450 GND.n449 7.147
R877 GND.n453 GND.n452 7.147
R878 GND.n456 GND.n455 7.147
R879 GND.n459 GND.n458 7.147
R880 GND.n462 GND.n461 7.147
R881 GND.n465 GND.n464 7.147
R882 GND.n468 GND.n467 7.147
R883 GND.n472 GND.n471 7.147
R884 GND.n475 GND.n474 7.147
R885 GND.n480 GND.n479 7.147
R886 GND.n483 GND.n482 7.147
R887 GND.n486 GND.n485 7.147
R888 GND.n491 GND.n490 7.147
R889 GND.n494 GND.n493 7.147
R890 GND.n497 GND.n496 7.147
R891 GND.n501 GND.n500 7.147
R892 GND.n504 GND.n503 7.147
R893 GND.n507 GND.n506 7.147
R894 GND.n510 GND.n509 7.147
R895 GND.n515 GND.n514 7.147
R896 GND.n518 GND.n517 7.147
R897 GND.n521 GND.n520 7.147
R898 GND.n524 GND.n523 7.147
R899 GND.n529 GND.n528 7.147
R900 GND.n532 GND.n531 7.147
R901 GND.n535 GND.n534 7.147
R902 GND.n538 GND.n537 7.147
R903 GND.n541 GND.n540 7.147
R904 GND.n544 GND.n543 7.147
R905 GND.n547 GND.n546 7.147
R906 GND.n551 GND.n550 7.147
R907 GND.n554 GND.n553 7.147
R908 GND.n559 GND.n558 7.147
R909 GND.n562 GND.n561 7.147
R910 GND.n565 GND.n564 7.147
R911 GND.n570 GND.n569 7.147
R912 GND.n573 GND.n572 7.147
R913 GND.n576 GND.n575 7.147
R914 GND.n580 GND.n579 7.147
R915 GND.n583 GND.n582 7.147
R916 GND.n586 GND.n585 7.147
R917 GND.n589 GND.n588 7.147
R918 GND.n594 GND.n593 7.147
R919 GND.n597 GND.n596 7.147
R920 GND.n600 GND.n599 7.147
R921 GND.n603 GND.n602 7.147
R922 GND.n608 GND.n607 7.147
R923 GND.n611 GND.n610 7.147
R924 GND.n614 GND.n613 7.147
R925 GND.n617 GND.n616 7.147
R926 GND.n620 GND.n619 7.147
R927 GND.n623 GND.n622 7.147
R928 GND.n626 GND.n625 7.147
R929 GND.n630 GND.n629 7.147
R930 GND.n633 GND.n632 7.147
R931 GND.n3 GND.n2 7.147
R932 GND.n6 GND.n5 7.147
R933 GND.n8 GND.n7 7.147
R934 GND.n10 GND.n9 7.147
R935 GND.n13 GND.n12 7.147
R936 GND.n15 GND.n14 7.147
R937 GND.n1555 GND.n1554 7.147
R938 GND.n1571 GND.n1570 7.147
R939 GND.n1569 GND.n1568 7.147
R940 GND.n1567 GND.n1566 7.147
R941 GND.n1564 GND.n1563 7.147
R942 GND.n1562 GND.n1561 7.147
R943 GND.n1560 GND.n1559 7.147
R944 GND.n1558 GND.n1557 7.147
R945 GND.n1544 GND.n1543 7.147
R946 GND.n1539 GND.n1538 7.147
R947 GND.n1536 GND.n1535 7.147
R948 GND.n1533 GND.n1532 7.147
R949 GND.n1530 GND.n1529 7.147
R950 GND.n1527 GND.n1526 7.147
R951 GND.n1524 GND.n1523 7.147
R952 GND.n1521 GND.n1520 7.147
R953 GND.n1517 GND.n1516 7.147
R954 GND.n1514 GND.n1513 7.147
R955 GND.n1509 GND.n1508 7.147
R956 GND.n1506 GND.n1505 7.147
R957 GND.n1503 GND.n1502 7.147
R958 GND.n1498 GND.n1497 7.147
R959 GND.n1495 GND.n1494 7.147
R960 GND.n1492 GND.n1491 7.147
R961 GND.n1488 GND.n1487 7.147
R962 GND.n1485 GND.n1484 7.147
R963 GND.n1482 GND.n1481 7.147
R964 GND.n1479 GND.n1478 7.147
R965 GND.n1474 GND.n1473 7.147
R966 GND.n1471 GND.n1470 7.147
R967 GND.n1468 GND.n1467 7.147
R968 GND.n1465 GND.n1464 7.147
R969 GND.n1460 GND.n1459 7.147
R970 GND.n1457 GND.n1456 7.147
R971 GND.n1454 GND.n1453 7.147
R972 GND.n1451 GND.n1450 7.147
R973 GND.n1448 GND.n1447 7.147
R974 GND.n1445 GND.n1444 7.147
R975 GND.n1442 GND.n1441 7.147
R976 GND.n1438 GND.n1437 7.147
R977 GND.n1435 GND.n1434 7.147
R978 GND.n1430 GND.n1429 7.147
R979 GND.n1427 GND.n1426 7.147
R980 GND.n1424 GND.n1423 7.147
R981 GND.n1419 GND.n1418 7.147
R982 GND.n1416 GND.n1415 7.147
R983 GND.n1413 GND.n1412 7.147
R984 GND.n1409 GND.n1408 7.147
R985 GND.n1406 GND.n1405 7.147
R986 GND.n1403 GND.n1402 7.147
R987 GND.n1400 GND.n1399 7.147
R988 GND.n1395 GND.n1394 7.147
R989 GND.n1392 GND.n1391 7.147
R990 GND.n1389 GND.n1388 7.147
R991 GND.n1386 GND.n1385 7.147
R992 GND.n1381 GND.n1380 7.147
R993 GND.n1378 GND.n1377 7.147
R994 GND.n1375 GND.n1374 7.147
R995 GND.n1372 GND.n1371 7.147
R996 GND.n1369 GND.n1368 7.147
R997 GND.n1366 GND.n1365 7.147
R998 GND.n1363 GND.n1362 7.147
R999 GND.n1359 GND.n1358 7.147
R1000 GND.n1356 GND.n1355 7.147
R1001 GND.n1351 GND.n1350 7.147
R1002 GND.n1348 GND.n1347 7.147
R1003 GND.n1345 GND.n1344 7.147
R1004 GND.n1340 GND.n1339 7.147
R1005 GND.n1337 GND.n1336 7.147
R1006 GND.n1334 GND.n1333 7.147
R1007 GND.n1330 GND.n1329 7.147
R1008 GND.n1327 GND.n1326 7.147
R1009 GND.n1324 GND.n1323 7.147
R1010 GND.n1321 GND.n1320 7.147
R1011 GND.n1316 GND.n1315 7.147
R1012 GND.n1313 GND.n1312 7.147
R1013 GND.n1310 GND.n1309 7.147
R1014 GND.n1307 GND.n1306 7.147
R1015 GND.n1302 GND.n1301 7.147
R1016 GND.n1299 GND.n1298 7.147
R1017 GND.n1296 GND.n1295 7.147
R1018 GND.n1293 GND.n1292 7.147
R1019 GND.n1290 GND.n1289 7.147
R1020 GND.n1287 GND.n1286 7.147
R1021 GND.n1284 GND.n1283 7.147
R1022 GND.n1280 GND.n1279 7.147
R1023 GND.n1277 GND.n1276 7.147
R1024 GND.n1272 GND.n1271 7.147
R1025 GND.n1269 GND.n1268 7.147
R1026 GND.n1266 GND.n1265 7.147
R1027 GND.n1261 GND.n1260 7.147
R1028 GND.n1258 GND.n1257 7.147
R1029 GND.n1255 GND.n1254 7.147
R1030 GND.n1251 GND.n1250 7.147
R1031 GND.n1248 GND.n1247 7.147
R1032 GND.n1245 GND.n1244 7.147
R1033 GND.n1242 GND.n1241 7.147
R1034 GND.n1237 GND.n1236 7.147
R1035 GND.n1234 GND.n1233 7.147
R1036 GND.n1231 GND.n1230 7.147
R1037 GND.n1228 GND.n1227 7.147
R1038 GND.n1223 GND.n1222 7.147
R1039 GND.n1220 GND.n1219 7.147
R1040 GND.n1217 GND.n1216 7.147
R1041 GND.n1214 GND.n1213 7.147
R1042 GND.n1211 GND.n1210 7.147
R1043 GND.n1208 GND.n1207 7.147
R1044 GND.n1205 GND.n1204 7.147
R1045 GND.n1201 GND.n1200 7.147
R1046 GND.n1198 GND.n1197 7.147
R1047 GND.n1193 GND.n1192 7.147
R1048 GND.n1190 GND.n1189 7.147
R1049 GND.n1187 GND.n1186 7.147
R1050 GND.n1182 GND.n1181 7.147
R1051 GND.n1179 GND.n1178 7.147
R1052 GND.n1176 GND.n1175 7.147
R1053 GND.n1172 GND.n1171 7.147
R1054 GND.n1169 GND.n1168 7.147
R1055 GND.n1166 GND.n1165 7.147
R1056 GND.n1163 GND.n1162 7.147
R1057 GND.n1158 GND.n1157 7.147
R1058 GND.n1155 GND.n1154 7.147
R1059 GND.n1152 GND.n1151 7.147
R1060 GND.n1149 GND.n1148 7.147
R1061 GND.n1144 GND.n1143 7.147
R1062 GND.n1141 GND.n1140 7.147
R1063 GND.n1138 GND.n1137 7.147
R1064 GND.n1135 GND.n1134 7.147
R1065 GND.n1132 GND.n1131 7.147
R1066 GND.n1129 GND.n1128 7.147
R1067 GND.n1126 GND.n1125 7.147
R1068 GND.n1122 GND.n1121 7.147
R1069 GND.n1119 GND.n1118 7.147
R1070 GND.n1114 GND.n1113 7.147
R1071 GND.n1111 GND.n1110 7.147
R1072 GND.n1108 GND.n1107 7.147
R1073 GND.n1103 GND.n1102 7.147
R1074 GND.n1100 GND.n1099 7.147
R1075 GND.n1097 GND.n1096 7.147
R1076 GND.n1093 GND.n1092 7.147
R1077 GND.n1090 GND.n1089 7.147
R1078 GND.n1087 GND.n1086 7.147
R1079 GND.n1084 GND.n1083 7.147
R1080 GND.n1079 GND.n1078 7.147
R1081 GND.n1076 GND.n1075 7.147
R1082 GND.n1073 GND.n1072 7.147
R1083 GND.n1070 GND.n1069 7.147
R1084 GND.n1065 GND.n1064 7.147
R1085 GND.n1062 GND.n1061 7.147
R1086 GND.n1059 GND.n1058 7.147
R1087 GND.n1056 GND.n1055 7.147
R1088 GND.n1053 GND.n1052 7.147
R1089 GND.n1050 GND.n1049 7.147
R1090 GND.n1047 GND.n1046 7.147
R1091 GND.n1043 GND.n1042 7.147
R1092 GND.n1040 GND.n1039 7.147
R1093 GND.n1035 GND.n1034 7.147
R1094 GND.n1032 GND.n1031 7.147
R1095 GND.n1029 GND.n1028 7.147
R1096 GND.n1024 GND.n1023 7.147
R1097 GND.n1021 GND.n1020 7.147
R1098 GND.n1018 GND.n1017 7.147
R1099 GND.n1014 GND.n1013 7.147
R1100 GND.n1011 GND.n1010 7.147
R1101 GND.n1008 GND.n1007 7.147
R1102 GND.n1005 GND.n1004 7.147
R1103 GND.n1000 GND.n999 7.147
R1104 GND.n997 GND.n996 7.147
R1105 GND.n994 GND.n993 7.147
R1106 GND.n991 GND.n990 7.147
R1107 GND.n986 GND.n985 7.147
R1108 GND.n983 GND.n982 7.147
R1109 GND.n980 GND.n979 7.147
R1110 GND.n977 GND.n976 7.147
R1111 GND.n974 GND.n973 7.147
R1112 GND.n971 GND.n970 7.147
R1113 GND.n968 GND.n967 7.147
R1114 GND.n964 GND.n963 7.147
R1115 GND.n961 GND.n960 7.147
R1116 GND.n956 GND.n955 7.147
R1117 GND.n953 GND.n952 7.147
R1118 GND.n950 GND.n949 7.147
R1119 GND.n945 GND.n944 7.147
R1120 GND.n942 GND.n941 7.147
R1121 GND.n939 GND.n938 7.147
R1122 GND.n935 GND.n934 7.147
R1123 GND.n932 GND.n931 7.147
R1124 GND.n929 GND.n928 7.147
R1125 GND.n926 GND.n925 7.147
R1126 GND.n921 GND.n920 7.147
R1127 GND.n918 GND.n917 7.147
R1128 GND.n915 GND.n914 7.147
R1129 GND.n912 GND.n911 7.147
R1130 GND.n907 GND.n906 7.147
R1131 GND.n904 GND.n903 7.147
R1132 GND.n901 GND.n900 7.147
R1133 GND.n898 GND.n897 7.147
R1134 GND.n895 GND.n894 7.147
R1135 GND.n892 GND.n891 7.147
R1136 GND.n889 GND.n888 7.147
R1137 GND.n885 GND.n884 7.147
R1138 GND.n882 GND.n881 7.147
R1139 GND.n877 GND.n876 7.147
R1140 GND.n874 GND.n873 7.147
R1141 GND.n871 GND.n870 7.147
R1142 GND.n866 GND.n865 7.147
R1143 GND.n863 GND.n862 7.147
R1144 GND.n860 GND.n859 7.147
R1145 GND.n856 GND.n855 7.147
R1146 GND.n853 GND.n852 7.147
R1147 GND.n850 GND.n849 7.147
R1148 GND.n847 GND.n846 7.147
R1149 GND.n842 GND.n841 7.147
R1150 GND.n839 GND.n838 7.147
R1151 GND.n836 GND.n835 7.147
R1152 GND.n833 GND.n832 7.147
R1153 GND.n828 GND.n827 7.147
R1154 GND.n825 GND.n824 7.147
R1155 GND.n822 GND.n821 7.147
R1156 GND.n819 GND.n818 7.147
R1157 GND.n816 GND.n815 7.147
R1158 GND.n813 GND.n812 7.147
R1159 GND.n810 GND.n809 7.147
R1160 GND.n806 GND.n805 7.147
R1161 GND.n803 GND.n802 7.147
R1162 GND.n798 GND.n797 7.147
R1163 GND.n795 GND.n794 7.147
R1164 GND.n792 GND.n791 7.147
R1165 GND.n787 GND.n786 7.147
R1166 GND.n784 GND.n783 7.147
R1167 GND.n781 GND.n780 7.147
R1168 GND.n777 GND.n776 7.147
R1169 GND.n774 GND.n773 7.147
R1170 GND.n771 GND.n770 7.147
R1171 GND.n768 GND.n767 7.147
R1172 GND.n763 GND.n762 7.147
R1173 GND.n760 GND.n759 7.147
R1174 GND.n757 GND.n756 7.147
R1175 GND.n754 GND.n753 7.147
R1176 GND.n749 GND.n748 7.147
R1177 GND.n746 GND.n745 7.147
R1178 GND.n743 GND.n742 7.147
R1179 GND.n740 GND.n739 7.147
R1180 GND.n737 GND.n736 7.147
R1181 GND.n734 GND.n733 7.147
R1182 GND.n731 GND.n730 7.147
R1183 GND.n727 GND.n726 7.147
R1184 GND.n724 GND.n723 7.147
R1185 GND.n719 GND.n718 7.147
R1186 GND.n716 GND.n715 7.147
R1187 GND.n713 GND.n712 7.147
R1188 GND.n708 GND.n707 7.147
R1189 GND.n705 GND.n704 7.147
R1190 GND.n702 GND.n701 7.147
R1191 GND.n698 GND.n697 7.147
R1192 GND.n695 GND.n694 7.147
R1193 GND.n692 GND.n691 7.147
R1194 GND.n689 GND.n688 7.147
R1195 GND.n684 GND.n683 7.147
R1196 GND.n681 GND.n680 7.147
R1197 GND.n678 GND.n677 7.147
R1198 GND.n675 GND.n674 7.147
R1199 GND.n670 GND.n669 7.147
R1200 GND.n667 GND.n666 7.147
R1201 GND.n664 GND.n663 7.147
R1202 GND.n661 GND.n660 7.147
R1203 GND.n658 GND.n657 7.147
R1204 GND.n655 GND.n654 7.147
R1205 GND.n652 GND.n651 7.147
R1206 GND.n648 GND.n647 7.147
R1207 GND.n55 GND.n53 6.264
R1208 GND.n134 GND.n132 6.264
R1209 GND.n213 GND.n211 6.264
R1210 GND.n292 GND.n290 6.264
R1211 GND.n371 GND.n369 6.264
R1212 GND.n450 GND.n448 6.264
R1213 GND.n529 GND.n527 6.264
R1214 GND.n608 GND.n606 6.264
R1215 GND.n1544 GND.n1542 6.264
R1216 GND.n1465 GND.n1463 6.264
R1217 GND.n1386 GND.n1384 6.264
R1218 GND.n1307 GND.n1305 6.264
R1219 GND.n1228 GND.n1226 6.264
R1220 GND.n1149 GND.n1147 6.264
R1221 GND.n1070 GND.n1068 6.264
R1222 GND.n991 GND.n989 6.264
R1223 GND.n912 GND.n910 6.264
R1224 GND.n833 GND.n831 6.264
R1225 GND.n754 GND.n752 6.264
R1226 GND.n675 GND.n673 6.264
R1227 GND.n41 GND.n39 4.286
R1228 GND.n120 GND.n118 4.286
R1229 GND.n199 GND.n197 4.286
R1230 GND.n278 GND.n276 4.286
R1231 GND.n357 GND.n355 4.286
R1232 GND.n436 GND.n434 4.286
R1233 GND.n515 GND.n513 4.286
R1234 GND.n594 GND.n592 4.286
R1235 GND.n1565 GND.n1564 4.286
R1236 GND.n1479 GND.n1477 4.286
R1237 GND.n1400 GND.n1398 4.286
R1238 GND.n1321 GND.n1319 4.286
R1239 GND.n1242 GND.n1240 4.286
R1240 GND.n1163 GND.n1161 4.286
R1241 GND.n1084 GND.n1082 4.286
R1242 GND.n1005 GND.n1003 4.286
R1243 GND.n926 GND.n924 4.286
R1244 GND.n847 GND.n845 4.286
R1245 GND.n768 GND.n766 4.286
R1246 GND.n689 GND.n687 4.286
R1247 GND.n77 GND.n75 3.297
R1248 GND.n156 GND.n154 3.297
R1249 GND.n235 GND.n233 3.297
R1250 GND.n314 GND.n312 3.297
R1251 GND.n393 GND.n391 3.297
R1252 GND.n472 GND.n470 3.297
R1253 GND.n551 GND.n549 3.297
R1254 GND.n630 GND.n628 3.297
R1255 GND.n1521 GND.n1519 3.297
R1256 GND.n1442 GND.n1440 3.297
R1257 GND.n1363 GND.n1361 3.297
R1258 GND.n1284 GND.n1282 3.297
R1259 GND.n1205 GND.n1203 3.297
R1260 GND.n1126 GND.n1124 3.297
R1261 GND.n1047 GND.n1045 3.297
R1262 GND.n968 GND.n966 3.297
R1263 GND.n889 GND.n887 3.297
R1264 GND.n810 GND.n808 3.297
R1265 GND.n731 GND.n729 3.297
R1266 GND.n652 GND.n650 3.297
R1267 GND.n27 GND.n25 2.967
R1268 GND.n106 GND.n104 2.967
R1269 GND.n185 GND.n183 2.967
R1270 GND.n264 GND.n262 2.967
R1271 GND.n343 GND.n341 2.967
R1272 GND.n422 GND.n420 2.967
R1273 GND.n501 GND.n499 2.967
R1274 GND.n580 GND.n578 2.967
R1275 GND.n1572 GND.n1555 2.967
R1276 GND.n1492 GND.n1490 2.967
R1277 GND.n1413 GND.n1411 2.967
R1278 GND.n1334 GND.n1332 2.967
R1279 GND.n1255 GND.n1253 2.967
R1280 GND.n1176 GND.n1174 2.967
R1281 GND.n1097 GND.n1095 2.967
R1282 GND.n1018 GND.n1016 2.967
R1283 GND.n939 GND.n937 2.967
R1284 GND.n860 GND.n858 2.967
R1285 GND.n781 GND.n779 2.967
R1286 GND.n702 GND.n700 2.967
R1287 GND.n20 GND.n19 1.568
R1288 GND.n96 GND.n94 1.483
R1289 GND.n175 GND.n173 1.483
R1290 GND.n254 GND.n252 1.483
R1291 GND.n333 GND.n331 1.483
R1292 GND.n412 GND.n410 1.483
R1293 GND.n491 GND.n489 1.483
R1294 GND.n570 GND.n568 1.483
R1295 GND.n11 GND.n10 1.483
R1296 GND.n1503 GND.n1501 1.483
R1297 GND.n1424 GND.n1422 1.483
R1298 GND.n1345 GND.n1343 1.483
R1299 GND.n1266 GND.n1264 1.483
R1300 GND.n1187 GND.n1185 1.483
R1301 GND.n1108 GND.n1106 1.483
R1302 GND.n1029 GND.n1027 1.483
R1303 GND.n950 GND.n948 1.483
R1304 GND.n871 GND.n869 1.483
R1305 GND.n792 GND.n790 1.483
R1306 GND.n713 GND.n711 1.483
R1307 GND.n85 GND.n83 0.329
R1308 GND.n164 GND.n162 0.329
R1309 GND.n243 GND.n241 0.329
R1310 GND.n322 GND.n320 0.329
R1311 GND.n401 GND.n399 0.329
R1312 GND.n480 GND.n478 0.329
R1313 GND.n559 GND.n557 0.329
R1314 GND.n4 GND.n3 0.329
R1315 GND.n1514 GND.n1512 0.329
R1316 GND.n1435 GND.n1433 0.329
R1317 GND.n1356 GND.n1354 0.329
R1318 GND.n1277 GND.n1275 0.329
R1319 GND.n1198 GND.n1196 0.329
R1320 GND.n1119 GND.n1117 0.329
R1321 GND.n1040 GND.n1038 0.329
R1322 GND.n961 GND.n959 0.329
R1323 GND.n882 GND.n880 0.329
R1324 GND.n803 GND.n801 0.329
R1325 GND.n724 GND.n722 0.329
R1326 GND.n645 GND.n644 0.329
R1327 GND.n24 GND.n21 0.119
R1328 GND.n28 GND.n24 0.119
R1329 GND.n31 GND.n28 0.119
R1330 GND.n34 GND.n31 0.119
R1331 GND.n37 GND.n34 0.119
R1332 GND.n42 GND.n37 0.119
R1333 GND.n45 GND.n42 0.119
R1334 GND.n48 GND.n45 0.119
R1335 GND.n51 GND.n48 0.119
R1336 GND.n56 GND.n51 0.119
R1337 GND.n59 GND.n56 0.119
R1338 GND.n62 GND.n59 0.119
R1339 GND.n65 GND.n62 0.119
R1340 GND.n68 GND.n65 0.119
R1341 GND.n71 GND.n68 0.119
R1342 GND.n74 GND.n71 0.119
R1343 GND.n78 GND.n74 0.119
R1344 GND.n81 GND.n78 0.119
R1345 GND.n86 GND.n81 0.119
R1346 GND.n89 GND.n86 0.119
R1347 GND.n92 GND.n89 0.119
R1348 GND.n97 GND.n92 0.119
R1349 GND.n100 GND.n97 0.119
R1350 GND.n103 GND.n100 0.119
R1351 GND.n107 GND.n103 0.119
R1352 GND.n110 GND.n107 0.119
R1353 GND.n113 GND.n110 0.119
R1354 GND.n116 GND.n113 0.119
R1355 GND.n121 GND.n116 0.119
R1356 GND.n124 GND.n121 0.119
R1357 GND.n127 GND.n124 0.119
R1358 GND.n130 GND.n127 0.119
R1359 GND.n135 GND.n130 0.119
R1360 GND.n138 GND.n135 0.119
R1361 GND.n141 GND.n138 0.119
R1362 GND.n144 GND.n141 0.119
R1363 GND.n147 GND.n144 0.119
R1364 GND.n150 GND.n147 0.119
R1365 GND.n153 GND.n150 0.119
R1366 GND.n157 GND.n153 0.119
R1367 GND.n160 GND.n157 0.119
R1368 GND.n165 GND.n160 0.119
R1369 GND.n168 GND.n165 0.119
R1370 GND.n171 GND.n168 0.119
R1371 GND.n176 GND.n171 0.119
R1372 GND.n179 GND.n176 0.119
R1373 GND.n182 GND.n179 0.119
R1374 GND.n186 GND.n182 0.119
R1375 GND.n189 GND.n186 0.119
R1376 GND.n192 GND.n189 0.119
R1377 GND.n195 GND.n192 0.119
R1378 GND.n200 GND.n195 0.119
R1379 GND.n203 GND.n200 0.119
R1380 GND.n206 GND.n203 0.119
R1381 GND.n209 GND.n206 0.119
R1382 GND.n214 GND.n209 0.119
R1383 GND.n217 GND.n214 0.119
R1384 GND.n220 GND.n217 0.119
R1385 GND.n223 GND.n220 0.119
R1386 GND.n226 GND.n223 0.119
R1387 GND.n229 GND.n226 0.119
R1388 GND.n232 GND.n229 0.119
R1389 GND.n236 GND.n232 0.119
R1390 GND.n239 GND.n236 0.119
R1391 GND.n244 GND.n239 0.119
R1392 GND.n247 GND.n244 0.119
R1393 GND.n250 GND.n247 0.119
R1394 GND.n255 GND.n250 0.119
R1395 GND.n258 GND.n255 0.119
R1396 GND.n261 GND.n258 0.119
R1397 GND.n265 GND.n261 0.119
R1398 GND.n268 GND.n265 0.119
R1399 GND.n271 GND.n268 0.119
R1400 GND.n274 GND.n271 0.119
R1401 GND.n279 GND.n274 0.119
R1402 GND.n282 GND.n279 0.119
R1403 GND.n285 GND.n282 0.119
R1404 GND.n288 GND.n285 0.119
R1405 GND.n293 GND.n288 0.119
R1406 GND.n296 GND.n293 0.119
R1407 GND.n299 GND.n296 0.119
R1408 GND.n302 GND.n299 0.119
R1409 GND.n305 GND.n302 0.119
R1410 GND.n308 GND.n305 0.119
R1411 GND.n311 GND.n308 0.119
R1412 GND.n315 GND.n311 0.119
R1413 GND.n318 GND.n315 0.119
R1414 GND.n323 GND.n318 0.119
R1415 GND.n326 GND.n323 0.119
R1416 GND.n329 GND.n326 0.119
R1417 GND.n334 GND.n329 0.119
R1418 GND.n337 GND.n334 0.119
R1419 GND.n340 GND.n337 0.119
R1420 GND.n344 GND.n340 0.119
R1421 GND.n347 GND.n344 0.119
R1422 GND.n350 GND.n347 0.119
R1423 GND.n353 GND.n350 0.119
R1424 GND.n358 GND.n353 0.119
R1425 GND.n361 GND.n358 0.119
R1426 GND.n364 GND.n361 0.119
R1427 GND.n367 GND.n364 0.119
R1428 GND.n372 GND.n367 0.119
R1429 GND.n375 GND.n372 0.119
R1430 GND.n378 GND.n375 0.119
R1431 GND.n381 GND.n378 0.119
R1432 GND.n384 GND.n381 0.119
R1433 GND.n387 GND.n384 0.119
R1434 GND.n390 GND.n387 0.119
R1435 GND.n394 GND.n390 0.119
R1436 GND.n397 GND.n394 0.119
R1437 GND.n402 GND.n397 0.119
R1438 GND.n405 GND.n402 0.119
R1439 GND.n408 GND.n405 0.119
R1440 GND.n413 GND.n408 0.119
R1441 GND.n416 GND.n413 0.119
R1442 GND.n419 GND.n416 0.119
R1443 GND.n423 GND.n419 0.119
R1444 GND.n426 GND.n423 0.119
R1445 GND.n429 GND.n426 0.119
R1446 GND.n432 GND.n429 0.119
R1447 GND.n437 GND.n432 0.119
R1448 GND.n440 GND.n437 0.119
R1449 GND.n443 GND.n440 0.119
R1450 GND.n446 GND.n443 0.119
R1451 GND.n451 GND.n446 0.119
R1452 GND.n454 GND.n451 0.119
R1453 GND.n457 GND.n454 0.119
R1454 GND.n460 GND.n457 0.119
R1455 GND.n463 GND.n460 0.119
R1456 GND.n466 GND.n463 0.119
R1457 GND.n469 GND.n466 0.119
R1458 GND.n473 GND.n469 0.119
R1459 GND.n476 GND.n473 0.119
R1460 GND.n481 GND.n476 0.119
R1461 GND.n484 GND.n481 0.119
R1462 GND.n487 GND.n484 0.119
R1463 GND.n492 GND.n487 0.119
R1464 GND.n495 GND.n492 0.119
R1465 GND.n498 GND.n495 0.119
R1466 GND.n502 GND.n498 0.119
R1467 GND.n505 GND.n502 0.119
R1468 GND.n508 GND.n505 0.119
R1469 GND.n511 GND.n508 0.119
R1470 GND.n516 GND.n511 0.119
R1471 GND.n519 GND.n516 0.119
R1472 GND.n522 GND.n519 0.119
R1473 GND.n525 GND.n522 0.119
R1474 GND.n530 GND.n525 0.119
R1475 GND.n533 GND.n530 0.119
R1476 GND.n536 GND.n533 0.119
R1477 GND.n539 GND.n536 0.119
R1478 GND.n542 GND.n539 0.119
R1479 GND.n545 GND.n542 0.119
R1480 GND.n548 GND.n545 0.119
R1481 GND.n552 GND.n548 0.119
R1482 GND.n555 GND.n552 0.119
R1483 GND.n560 GND.n555 0.119
R1484 GND.n563 GND.n560 0.119
R1485 GND.n566 GND.n563 0.119
R1486 GND.n571 GND.n566 0.119
R1487 GND.n574 GND.n571 0.119
R1488 GND.n577 GND.n574 0.119
R1489 GND.n581 GND.n577 0.119
R1490 GND.n584 GND.n581 0.119
R1491 GND.n587 GND.n584 0.119
R1492 GND.n590 GND.n587 0.119
R1493 GND.n595 GND.n590 0.119
R1494 GND.n598 GND.n595 0.119
R1495 GND.n601 GND.n598 0.119
R1496 GND.n604 GND.n601 0.119
R1497 GND.n609 GND.n604 0.119
R1498 GND.n612 GND.n609 0.119
R1499 GND.n615 GND.n612 0.119
R1500 GND.n618 GND.n615 0.119
R1501 GND.n621 GND.n618 0.119
R1502 GND.n624 GND.n621 0.119
R1503 GND.n627 GND.n624 0.119
R1504 GND.n631 GND.n627 0.119
R1505 GND.n634 GND.n631 0.119
R1506 GND.n635 GND.n634 0.119
R1507 GND.n636 GND.n635 0.119
R1508 GND.n637 GND.n636 0.119
R1509 GND.n638 GND.n637 0.119
R1510 GND.n639 GND.n638 0.119
R1511 GND.n640 GND.n639 0.119
R1512 GND.n1553 GND.n640 0.119
R1513 GND.n1553 GND.n1552 0.119
R1514 GND.n1552 GND.n1551 0.119
R1515 GND.n1551 GND.n1550 0.119
R1516 GND.n1550 GND.n1549 0.119
R1517 GND.n1549 GND.n1548 0.119
R1518 GND.n1548 GND.n1547 0.119
R1519 GND.n1547 GND.n1546 0.119
R1520 GND.n1546 GND.n1545 0.119
R1521 GND.n1545 GND.n1540 0.119
R1522 GND.n1540 GND.n1537 0.119
R1523 GND.n1537 GND.n1534 0.119
R1524 GND.n1534 GND.n1531 0.119
R1525 GND.n1531 GND.n1528 0.119
R1526 GND.n1528 GND.n1525 0.119
R1527 GND.n1525 GND.n1522 0.119
R1528 GND.n1522 GND.n1518 0.119
R1529 GND.n1518 GND.n1515 0.119
R1530 GND.n1515 GND.n1510 0.119
R1531 GND.n1510 GND.n1507 0.119
R1532 GND.n1507 GND.n1504 0.119
R1533 GND.n1504 GND.n1499 0.119
R1534 GND.n1499 GND.n1496 0.119
R1535 GND.n1496 GND.n1493 0.119
R1536 GND.n1493 GND.n1489 0.119
R1537 GND.n1489 GND.n1486 0.119
R1538 GND.n1486 GND.n1483 0.119
R1539 GND.n1483 GND.n1480 0.119
R1540 GND.n1480 GND.n1475 0.119
R1541 GND.n1475 GND.n1472 0.119
R1542 GND.n1472 GND.n1469 0.119
R1543 GND.n1469 GND.n1466 0.119
R1544 GND.n1466 GND.n1461 0.119
R1545 GND.n1461 GND.n1458 0.119
R1546 GND.n1458 GND.n1455 0.119
R1547 GND.n1455 GND.n1452 0.119
R1548 GND.n1452 GND.n1449 0.119
R1549 GND.n1449 GND.n1446 0.119
R1550 GND.n1446 GND.n1443 0.119
R1551 GND.n1443 GND.n1439 0.119
R1552 GND.n1439 GND.n1436 0.119
R1553 GND.n1436 GND.n1431 0.119
R1554 GND.n1431 GND.n1428 0.119
R1555 GND.n1428 GND.n1425 0.119
R1556 GND.n1425 GND.n1420 0.119
R1557 GND.n1420 GND.n1417 0.119
R1558 GND.n1417 GND.n1414 0.119
R1559 GND.n1414 GND.n1410 0.119
R1560 GND.n1410 GND.n1407 0.119
R1561 GND.n1407 GND.n1404 0.119
R1562 GND.n1404 GND.n1401 0.119
R1563 GND.n1401 GND.n1396 0.119
R1564 GND.n1396 GND.n1393 0.119
R1565 GND.n1393 GND.n1390 0.119
R1566 GND.n1390 GND.n1387 0.119
R1567 GND.n1387 GND.n1382 0.119
R1568 GND.n1382 GND.n1379 0.119
R1569 GND.n1379 GND.n1376 0.119
R1570 GND.n1376 GND.n1373 0.119
R1571 GND.n1373 GND.n1370 0.119
R1572 GND.n1370 GND.n1367 0.119
R1573 GND.n1367 GND.n1364 0.119
R1574 GND.n1364 GND.n1360 0.119
R1575 GND.n1360 GND.n1357 0.119
R1576 GND.n1357 GND.n1352 0.119
R1577 GND.n1352 GND.n1349 0.119
R1578 GND.n1349 GND.n1346 0.119
R1579 GND.n1346 GND.n1341 0.119
R1580 GND.n1341 GND.n1338 0.119
R1581 GND.n1338 GND.n1335 0.119
R1582 GND.n1335 GND.n1331 0.119
R1583 GND.n1331 GND.n1328 0.119
R1584 GND.n1328 GND.n1325 0.119
R1585 GND.n1325 GND.n1322 0.119
R1586 GND.n1322 GND.n1317 0.119
R1587 GND.n1317 GND.n1314 0.119
R1588 GND.n1314 GND.n1311 0.119
R1589 GND.n1311 GND.n1308 0.119
R1590 GND.n1308 GND.n1303 0.119
R1591 GND.n1303 GND.n1300 0.119
R1592 GND.n1300 GND.n1297 0.119
R1593 GND.n1297 GND.n1294 0.119
R1594 GND.n1294 GND.n1291 0.119
R1595 GND.n1291 GND.n1288 0.119
R1596 GND.n1288 GND.n1285 0.119
R1597 GND.n1285 GND.n1281 0.119
R1598 GND.n1281 GND.n1278 0.119
R1599 GND.n1278 GND.n1273 0.119
R1600 GND.n1273 GND.n1270 0.119
R1601 GND.n1270 GND.n1267 0.119
R1602 GND.n1267 GND.n1262 0.119
R1603 GND.n1262 GND.n1259 0.119
R1604 GND.n1259 GND.n1256 0.119
R1605 GND.n1256 GND.n1252 0.119
R1606 GND.n1252 GND.n1249 0.119
R1607 GND.n1249 GND.n1246 0.119
R1608 GND.n1246 GND.n1243 0.119
R1609 GND.n1243 GND.n1238 0.119
R1610 GND.n1238 GND.n1235 0.119
R1611 GND.n1235 GND.n1232 0.119
R1612 GND.n1232 GND.n1229 0.119
R1613 GND.n1229 GND.n1224 0.119
R1614 GND.n1224 GND.n1221 0.119
R1615 GND.n1221 GND.n1218 0.119
R1616 GND.n1218 GND.n1215 0.119
R1617 GND.n1215 GND.n1212 0.119
R1618 GND.n1212 GND.n1209 0.119
R1619 GND.n1209 GND.n1206 0.119
R1620 GND.n1206 GND.n1202 0.119
R1621 GND.n1202 GND.n1199 0.119
R1622 GND.n1199 GND.n1194 0.119
R1623 GND.n1194 GND.n1191 0.119
R1624 GND.n1191 GND.n1188 0.119
R1625 GND.n1188 GND.n1183 0.119
R1626 GND.n1183 GND.n1180 0.119
R1627 GND.n1180 GND.n1177 0.119
R1628 GND.n1177 GND.n1173 0.119
R1629 GND.n1173 GND.n1170 0.119
R1630 GND.n1170 GND.n1167 0.119
R1631 GND.n1167 GND.n1164 0.119
R1632 GND.n1164 GND.n1159 0.119
R1633 GND.n1159 GND.n1156 0.119
R1634 GND.n1156 GND.n1153 0.119
R1635 GND.n1153 GND.n1150 0.119
R1636 GND.n1150 GND.n1145 0.119
R1637 GND.n1145 GND.n1142 0.119
R1638 GND.n1142 GND.n1139 0.119
R1639 GND.n1139 GND.n1136 0.119
R1640 GND.n1136 GND.n1133 0.119
R1641 GND.n1133 GND.n1130 0.119
R1642 GND.n1130 GND.n1127 0.119
R1643 GND.n1127 GND.n1123 0.119
R1644 GND.n1123 GND.n1120 0.119
R1645 GND.n1120 GND.n1115 0.119
R1646 GND.n1115 GND.n1112 0.119
R1647 GND.n1112 GND.n1109 0.119
R1648 GND.n1109 GND.n1104 0.119
R1649 GND.n1104 GND.n1101 0.119
R1650 GND.n1101 GND.n1098 0.119
R1651 GND.n1098 GND.n1094 0.119
R1652 GND.n1094 GND.n1091 0.119
R1653 GND.n1091 GND.n1088 0.119
R1654 GND.n1088 GND.n1085 0.119
R1655 GND.n1085 GND.n1080 0.119
R1656 GND.n1080 GND.n1077 0.119
R1657 GND.n1077 GND.n1074 0.119
R1658 GND.n1074 GND.n1071 0.119
R1659 GND.n1071 GND.n1066 0.119
R1660 GND.n1066 GND.n1063 0.119
R1661 GND.n1063 GND.n1060 0.119
R1662 GND.n1060 GND.n1057 0.119
R1663 GND.n1057 GND.n1054 0.119
R1664 GND.n1054 GND.n1051 0.119
R1665 GND.n1051 GND.n1048 0.119
R1666 GND.n1048 GND.n1044 0.119
R1667 GND.n1044 GND.n1041 0.119
R1668 GND.n1041 GND.n1036 0.119
R1669 GND.n1036 GND.n1033 0.119
R1670 GND.n1033 GND.n1030 0.119
R1671 GND.n1030 GND.n1025 0.119
R1672 GND.n1025 GND.n1022 0.119
R1673 GND.n1022 GND.n1019 0.119
R1674 GND.n1019 GND.n1015 0.119
R1675 GND.n1015 GND.n1012 0.119
R1676 GND.n1012 GND.n1009 0.119
R1677 GND.n1009 GND.n1006 0.119
R1678 GND.n1006 GND.n1001 0.119
R1679 GND.n1001 GND.n998 0.119
R1680 GND.n998 GND.n995 0.119
R1681 GND.n995 GND.n992 0.119
R1682 GND.n992 GND.n987 0.119
R1683 GND.n987 GND.n984 0.119
R1684 GND.n984 GND.n981 0.119
R1685 GND.n981 GND.n978 0.119
R1686 GND.n978 GND.n975 0.119
R1687 GND.n975 GND.n972 0.119
R1688 GND.n972 GND.n969 0.119
R1689 GND.n969 GND.n965 0.119
R1690 GND.n965 GND.n962 0.119
R1691 GND.n962 GND.n957 0.119
R1692 GND.n957 GND.n954 0.119
R1693 GND.n954 GND.n951 0.119
R1694 GND.n951 GND.n946 0.119
R1695 GND.n946 GND.n943 0.119
R1696 GND.n943 GND.n940 0.119
R1697 GND.n940 GND.n936 0.119
R1698 GND.n936 GND.n933 0.119
R1699 GND.n933 GND.n930 0.119
R1700 GND.n930 GND.n927 0.119
R1701 GND.n927 GND.n922 0.119
R1702 GND.n922 GND.n919 0.119
R1703 GND.n919 GND.n916 0.119
R1704 GND.n916 GND.n913 0.119
R1705 GND.n913 GND.n908 0.119
R1706 GND.n908 GND.n905 0.119
R1707 GND.n905 GND.n902 0.119
R1708 GND.n902 GND.n899 0.119
R1709 GND.n899 GND.n896 0.119
R1710 GND.n896 GND.n893 0.119
R1711 GND.n893 GND.n890 0.119
R1712 GND.n890 GND.n886 0.119
R1713 GND.n886 GND.n883 0.119
R1714 GND.n883 GND.n878 0.119
R1715 GND.n878 GND.n875 0.119
R1716 GND.n875 GND.n872 0.119
R1717 GND.n872 GND.n867 0.119
R1718 GND.n867 GND.n864 0.119
R1719 GND.n864 GND.n861 0.119
R1720 GND.n861 GND.n857 0.119
R1721 GND.n857 GND.n854 0.119
R1722 GND.n854 GND.n851 0.119
R1723 GND.n851 GND.n848 0.119
R1724 GND.n848 GND.n843 0.119
R1725 GND.n843 GND.n840 0.119
R1726 GND.n840 GND.n837 0.119
R1727 GND.n837 GND.n834 0.119
R1728 GND.n834 GND.n829 0.119
R1729 GND.n829 GND.n826 0.119
R1730 GND.n826 GND.n823 0.119
R1731 GND.n823 GND.n820 0.119
R1732 GND.n820 GND.n817 0.119
R1733 GND.n817 GND.n814 0.119
R1734 GND.n814 GND.n811 0.119
R1735 GND.n811 GND.n807 0.119
R1736 GND.n807 GND.n804 0.119
R1737 GND.n804 GND.n799 0.119
R1738 GND.n799 GND.n796 0.119
R1739 GND.n796 GND.n793 0.119
R1740 GND.n793 GND.n788 0.119
R1741 GND.n788 GND.n785 0.119
R1742 GND.n785 GND.n782 0.119
R1743 GND.n782 GND.n778 0.119
R1744 GND.n778 GND.n775 0.119
R1745 GND.n775 GND.n772 0.119
R1746 GND.n772 GND.n769 0.119
R1747 GND.n769 GND.n764 0.119
R1748 GND.n764 GND.n761 0.119
R1749 GND.n761 GND.n758 0.119
R1750 GND.n758 GND.n755 0.119
R1751 GND.n755 GND.n750 0.119
R1752 GND.n750 GND.n747 0.119
R1753 GND.n747 GND.n744 0.119
R1754 GND.n744 GND.n741 0.119
R1755 GND.n741 GND.n738 0.119
R1756 GND.n738 GND.n735 0.119
R1757 GND.n735 GND.n732 0.119
R1758 GND.n732 GND.n728 0.119
R1759 GND.n728 GND.n725 0.119
R1760 GND.n725 GND.n720 0.119
R1761 GND.n720 GND.n717 0.119
R1762 GND.n717 GND.n714 0.119
R1763 GND.n714 GND.n709 0.119
R1764 GND.n709 GND.n706 0.119
R1765 GND.n706 GND.n703 0.119
R1766 GND.n703 GND.n699 0.119
R1767 GND.n699 GND.n696 0.119
R1768 GND.n696 GND.n693 0.119
R1769 GND.n693 GND.n690 0.119
R1770 GND.n690 GND.n685 0.119
R1771 GND.n685 GND.n682 0.119
R1772 GND.n682 GND.n679 0.119
R1773 GND.n679 GND.n676 0.119
R1774 GND.n676 GND.n671 0.119
R1775 GND.n671 GND.n668 0.119
R1776 GND.n668 GND.n665 0.119
R1777 GND.n665 GND.n662 0.119
R1778 GND.n662 GND.n659 0.119
R1779 GND.n659 GND.n656 0.119
R1780 GND.n656 GND.n653 0.119
R1781 GND.n653 GND.n649 0.119
R1782 GND.n649 GND.n646 0.119
R1783 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t6 389.181
R1784 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t3 256.987
R1785 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t8 212.079
R1786 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t7 174.888
R1787 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t4 163.801
R1788 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n0 161.578
R1789 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t5 139.779
R1790 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n1 129.263
R1791 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n5 102.015
R1792 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t1 63.321
R1793 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t2 63.321
R1794 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n6 46.071
R1795 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n3 37.442
R1796 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n4 23.54
R1797 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1283_21.n2 22.639
R1798 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.t3 239.038
R1799 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.t2 166.738
R1800 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n1 95.895
R1801 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.t1 71.217
R1802 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1847_47.n0 30.051
R1803 VDD.n1612 VDD.t239 225.592
R1804 VDD.n1529 VDD.t8 225.592
R1805 VDD.n1446 VDD.t52 225.592
R1806 VDD.n1363 VDD.t86 225.592
R1807 VDD.n1280 VDD.t63 225.592
R1808 VDD.n1197 VDD.t33 225.592
R1809 VDD.n52 VDD.t109 225.592
R1810 VDD.n135 VDD.t128 225.592
R1811 VDD.n218 VDD.t168 225.592
R1812 VDD.n301 VDD.t18 225.592
R1813 VDD.n384 VDD.t140 225.592
R1814 VDD.n467 VDD.t51 225.592
R1815 VDD.n550 VDD.t66 225.592
R1816 VDD.n633 VDD.t112 225.592
R1817 VDD.n716 VDD.t101 225.592
R1818 VDD.n799 VDD.t164 225.592
R1819 VDD.n882 VDD.t49 225.592
R1820 VDD.n965 VDD.t178 225.592
R1821 VDD.n1048 VDD.t100 225.592
R1822 VDD.n1131 VDD.t65 225.592
R1823 VDD.n1632 VDD.t26 119.607
R1824 VDD.n1542 VDD.t38 119.607
R1825 VDD.n1459 VDD.t80 119.607
R1826 VDD.n1376 VDD.t234 119.607
R1827 VDD.n1293 VDD.t34 119.607
R1828 VDD.n1210 VDD.t132 119.607
R1829 VDD.n38 VDD.t96 119.607
R1830 VDD.n121 VDD.t114 119.607
R1831 VDD.n204 VDD.t185 119.607
R1832 VDD.n287 VDD.t122 119.607
R1833 VDD.n370 VDD.t6 119.607
R1834 VDD.n453 VDD.t154 119.607
R1835 VDD.n536 VDD.t88 119.607
R1836 VDD.n619 VDD.t58 119.607
R1837 VDD.n702 VDD.t87 119.607
R1838 VDD.n785 VDD.t69 119.607
R1839 VDD.n868 VDD.t146 119.607
R1840 VDD.n951 VDD.t78 119.607
R1841 VDD.n1034 VDD.t236 119.607
R1842 VDD.n1117 VDD.t139 119.607
R1843 VDD.n1604 VDD.t53 93.809
R1844 VDD.n1521 VDD.t77 93.809
R1845 VDD.n1438 VDD.t20 93.809
R1846 VDD.n1355 VDD.t23 93.809
R1847 VDD.n1272 VDD.t30 93.809
R1848 VDD.n1189 VDD.t70 93.809
R1849 VDD.n59 VDD.t163 93.809
R1850 VDD.n142 VDD.t169 93.809
R1851 VDD.n225 VDD.t45 93.809
R1852 VDD.n308 VDD.t91 93.809
R1853 VDD.n391 VDD.t124 93.809
R1854 VDD.n474 VDD.t107 93.809
R1855 VDD.n557 VDD.t105 93.809
R1856 VDD.n640 VDD.t186 93.809
R1857 VDD.n723 VDD.t40 93.809
R1858 VDD.n806 VDD.t32 93.809
R1859 VDD.n889 VDD.t93 93.809
R1860 VDD.n972 VDD.t44 93.809
R1861 VDD.n1055 VDD.t85 93.809
R1862 VDD.n1138 VDD.t156 93.809
R1863 VDD.n1588 VDD.t0 85.217
R1864 VDD.n1505 VDD.t56 85.217
R1865 VDD.n1422 VDD.t98 85.217
R1866 VDD.n1339 VDD.t67 85.217
R1867 VDD.n1256 VDD.t59 85.217
R1868 VDD.n1173 VDD.t25 85.217
R1869 VDD.n76 VDD.t116 85.217
R1870 VDD.n159 VDD.t151 85.217
R1871 VDD.n242 VDD.t43 85.217
R1872 VDD.n325 VDD.t147 85.217
R1873 VDD.n408 VDD.t228 85.217
R1874 VDD.n491 VDD.t31 85.217
R1875 VDD.n574 VDD.t11 85.217
R1876 VDD.n657 VDD.t94 85.217
R1877 VDD.n740 VDD.t81 85.217
R1878 VDD.n823 VDD.t111 85.217
R1879 VDD.n906 VDD.t176 85.217
R1880 VDD.n989 VDD.t102 85.217
R1881 VDD.n1072 VDD.t159 85.217
R1882 VDD.n3 VDD.t84 85.217
R1883 VDD.n1109 VDD.t103 68.011
R1884 VDD.n1026 VDD.t113 68.011
R1885 VDD.n943 VDD.t184 68.011
R1886 VDD.n860 VDD.t142 68.011
R1887 VDD.n777 VDD.t15 68.011
R1888 VDD.n694 VDD.t173 68.011
R1889 VDD.n611 VDD.t55 68.011
R1890 VDD.n528 VDD.t76 68.011
R1891 VDD.n445 VDD.t36 68.011
R1892 VDD.n362 VDD.t137 68.011
R1893 VDD.n279 VDD.t129 68.011
R1894 VDD.n196 VDD.t134 68.011
R1895 VDD.n113 VDD.t177 68.011
R1896 VDD.n30 VDD.t180 68.011
R1897 VDD.n1220 VDD.t83 68.011
R1898 VDD.n1303 VDD.t74 68.011
R1899 VDD.n1386 VDD.t82 68.011
R1900 VDD.n1469 VDD.t41 68.011
R1901 VDD.n1552 VDD.t9 68.011
R1902 VDD.n1631 VDD.t175 68.011
R1903 VDD.n1604 VDD.t215 63.321
R1904 VDD.n1632 VDD.t216 63.321
R1905 VDD.n1521 VDD.t217 63.321
R1906 VDD.n1542 VDD.t218 63.321
R1907 VDD.n1438 VDD.t219 63.321
R1908 VDD.n1459 VDD.t220 63.321
R1909 VDD.n1355 VDD.t221 63.321
R1910 VDD.n1376 VDD.t222 63.321
R1911 VDD.n1272 VDD.t223 63.321
R1912 VDD.n1293 VDD.t224 63.321
R1913 VDD.n1189 VDD.t225 63.321
R1914 VDD.n1210 VDD.t226 63.321
R1915 VDD.n59 VDD.t187 63.321
R1916 VDD.n38 VDD.t188 63.321
R1917 VDD.n142 VDD.t189 63.321
R1918 VDD.n121 VDD.t190 63.321
R1919 VDD.n225 VDD.t191 63.321
R1920 VDD.n204 VDD.t192 63.321
R1921 VDD.n308 VDD.t193 63.321
R1922 VDD.n287 VDD.t194 63.321
R1923 VDD.n391 VDD.t195 63.321
R1924 VDD.n370 VDD.t196 63.321
R1925 VDD.n474 VDD.t197 63.321
R1926 VDD.n453 VDD.t198 63.321
R1927 VDD.n557 VDD.t199 63.321
R1928 VDD.n536 VDD.t200 63.321
R1929 VDD.n640 VDD.t201 63.321
R1930 VDD.n619 VDD.t202 63.321
R1931 VDD.n723 VDD.t203 63.321
R1932 VDD.n702 VDD.t204 63.321
R1933 VDD.n806 VDD.t205 63.321
R1934 VDD.n785 VDD.t206 63.321
R1935 VDD.n889 VDD.t207 63.321
R1936 VDD.n868 VDD.t208 63.321
R1937 VDD.n972 VDD.t209 63.321
R1938 VDD.n951 VDD.t210 63.321
R1939 VDD.n1055 VDD.t211 63.321
R1940 VDD.n1034 VDD.t212 63.321
R1941 VDD.n1138 VDD.t213 63.321
R1942 VDD.n1117 VDD.t214 63.321
R1943 VDD.n1566 VDD.t3 61.575
R1944 VDD.n1483 VDD.t64 61.575
R1945 VDD.n1400 VDD.t62 61.575
R1946 VDD.n1317 VDD.t60 61.575
R1947 VDD.n1234 VDD.t133 61.575
R1948 VDD.n16 VDD.t135 61.575
R1949 VDD.n97 VDD.t126 61.575
R1950 VDD.n180 VDD.t181 61.575
R1951 VDD.n263 VDD.t167 61.575
R1952 VDD.n346 VDD.t235 61.575
R1953 VDD.n429 VDD.t183 61.575
R1954 VDD.n512 VDD.t179 61.575
R1955 VDD.n595 VDD.t89 61.575
R1956 VDD.n678 VDD.t170 61.575
R1957 VDD.n761 VDD.t73 61.575
R1958 VDD.n844 VDD.t171 61.575
R1959 VDD.n927 VDD.t230 61.575
R1960 VDD.n1010 VDD.t13 61.575
R1961 VDD.n1093 VDD.t14 61.575
R1962 VDD.n1653 VDD.t237 61.562
R1963 VDD.n1166 VDD.n1161 50.786
R1964 VDD.n1621 VDD.n1620 50.667
R1965 VDD.n1618 VDD.n1617 50.667
R1966 VDD.n1615 VDD.n1614 50.667
R1967 VDD.n1611 VDD.n1610 50.667
R1968 VDD.n1608 VDD.n1607 50.667
R1969 VDD.n1603 VDD.n1602 50.667
R1970 VDD.n1600 VDD.n1599 50.667
R1971 VDD.n1597 VDD.n1596 50.667
R1972 VDD.n1594 VDD.n1593 50.667
R1973 VDD.n1591 VDD.n1590 50.667
R1974 VDD.n1587 VDD.n1586 50.667
R1975 VDD.n1584 VDD.n1583 50.667
R1976 VDD.n1581 VDD.n1580 50.667
R1977 VDD.n1576 VDD.n1575 50.667
R1978 VDD.n1573 VDD.n1572 50.667
R1979 VDD.n1570 VDD.n1569 50.667
R1980 VDD.n1565 VDD.n1564 50.667
R1981 VDD.n1562 VDD.n1561 50.667
R1982 VDD.n1559 VDD.n1558 50.667
R1983 VDD.n1556 VDD.n1555 50.667
R1984 VDD.n1549 VDD.n1548 50.667
R1985 VDD.n1546 VDD.n1545 50.667
R1986 VDD.n1541 VDD.n1540 50.667
R1987 VDD.n1538 VDD.n1537 50.667
R1988 VDD.n1535 VDD.n1534 50.667
R1989 VDD.n1532 VDD.n1531 50.667
R1990 VDD.n1528 VDD.n1527 50.667
R1991 VDD.n1525 VDD.n1524 50.667
R1992 VDD.n1520 VDD.n1519 50.667
R1993 VDD.n1517 VDD.n1516 50.667
R1994 VDD.n1514 VDD.n1513 50.667
R1995 VDD.n1511 VDD.n1510 50.667
R1996 VDD.n1508 VDD.n1507 50.667
R1997 VDD.n1504 VDD.n1503 50.667
R1998 VDD.n1501 VDD.n1500 50.667
R1999 VDD.n1498 VDD.n1497 50.667
R2000 VDD.n1493 VDD.n1492 50.667
R2001 VDD.n1490 VDD.n1489 50.667
R2002 VDD.n1487 VDD.n1486 50.667
R2003 VDD.n1482 VDD.n1481 50.667
R2004 VDD.n1479 VDD.n1478 50.667
R2005 VDD.n1476 VDD.n1475 50.667
R2006 VDD.n1473 VDD.n1472 50.667
R2007 VDD.n1466 VDD.n1465 50.667
R2008 VDD.n1463 VDD.n1462 50.667
R2009 VDD.n1458 VDD.n1457 50.667
R2010 VDD.n1455 VDD.n1454 50.667
R2011 VDD.n1452 VDD.n1451 50.667
R2012 VDD.n1449 VDD.n1448 50.667
R2013 VDD.n1445 VDD.n1444 50.667
R2014 VDD.n1442 VDD.n1441 50.667
R2015 VDD.n1437 VDD.n1436 50.667
R2016 VDD.n1434 VDD.n1433 50.667
R2017 VDD.n1431 VDD.n1430 50.667
R2018 VDD.n1428 VDD.n1427 50.667
R2019 VDD.n1425 VDD.n1424 50.667
R2020 VDD.n1421 VDD.n1420 50.667
R2021 VDD.n1418 VDD.n1417 50.667
R2022 VDD.n1415 VDD.n1414 50.667
R2023 VDD.n1410 VDD.n1409 50.667
R2024 VDD.n1407 VDD.n1406 50.667
R2025 VDD.n1404 VDD.n1403 50.667
R2026 VDD.n1399 VDD.n1398 50.667
R2027 VDD.n1396 VDD.n1395 50.667
R2028 VDD.n1393 VDD.n1392 50.667
R2029 VDD.n1390 VDD.n1389 50.667
R2030 VDD.n1383 VDD.n1382 50.667
R2031 VDD.n1380 VDD.n1379 50.667
R2032 VDD.n1375 VDD.n1374 50.667
R2033 VDD.n1372 VDD.n1371 50.667
R2034 VDD.n1369 VDD.n1368 50.667
R2035 VDD.n1366 VDD.n1365 50.667
R2036 VDD.n1362 VDD.n1361 50.667
R2037 VDD.n1359 VDD.n1358 50.667
R2038 VDD.n1354 VDD.n1353 50.667
R2039 VDD.n1351 VDD.n1350 50.667
R2040 VDD.n1348 VDD.n1347 50.667
R2041 VDD.n1345 VDD.n1344 50.667
R2042 VDD.n1342 VDD.n1341 50.667
R2043 VDD.n1338 VDD.n1337 50.667
R2044 VDD.n1335 VDD.n1334 50.667
R2045 VDD.n1332 VDD.n1331 50.667
R2046 VDD.n1327 VDD.n1326 50.667
R2047 VDD.n1324 VDD.n1323 50.667
R2048 VDD.n1321 VDD.n1320 50.667
R2049 VDD.n1316 VDD.n1315 50.667
R2050 VDD.n1313 VDD.n1312 50.667
R2051 VDD.n1310 VDD.n1309 50.667
R2052 VDD.n1307 VDD.n1306 50.667
R2053 VDD.n1300 VDD.n1299 50.667
R2054 VDD.n1297 VDD.n1296 50.667
R2055 VDD.n1292 VDD.n1291 50.667
R2056 VDD.n1289 VDD.n1288 50.667
R2057 VDD.n1286 VDD.n1285 50.667
R2058 VDD.n1283 VDD.n1282 50.667
R2059 VDD.n1279 VDD.n1278 50.667
R2060 VDD.n1276 VDD.n1275 50.667
R2061 VDD.n1271 VDD.n1270 50.667
R2062 VDD.n1268 VDD.n1267 50.667
R2063 VDD.n1265 VDD.n1264 50.667
R2064 VDD.n1262 VDD.n1261 50.667
R2065 VDD.n1259 VDD.n1258 50.667
R2066 VDD.n1255 VDD.n1254 50.667
R2067 VDD.n1252 VDD.n1251 50.667
R2068 VDD.n1249 VDD.n1248 50.667
R2069 VDD.n1244 VDD.n1243 50.667
R2070 VDD.n1241 VDD.n1240 50.667
R2071 VDD.n1238 VDD.n1237 50.667
R2072 VDD.n1233 VDD.n1232 50.667
R2073 VDD.n1230 VDD.n1229 50.667
R2074 VDD.n1227 VDD.n1226 50.667
R2075 VDD.n1224 VDD.n1223 50.667
R2076 VDD.n1217 VDD.n1216 50.667
R2077 VDD.n1214 VDD.n1213 50.667
R2078 VDD.n1209 VDD.n1208 50.667
R2079 VDD.n1206 VDD.n1205 50.667
R2080 VDD.n1203 VDD.n1202 50.667
R2081 VDD.n1200 VDD.n1199 50.667
R2082 VDD.n1196 VDD.n1195 50.667
R2083 VDD.n1193 VDD.n1192 50.667
R2084 VDD.n1188 VDD.n1187 50.667
R2085 VDD.n1185 VDD.n1184 50.667
R2086 VDD.n1182 VDD.n1181 50.667
R2087 VDD.n1179 VDD.n1178 50.667
R2088 VDD.n1176 VDD.n1175 50.667
R2089 VDD.n1172 VDD.n1171 50.667
R2090 VDD.n1169 VDD.n1168 50.667
R2091 VDD.n1166 VDD.n1165 50.667
R2092 VDD.n27 VDD.n26 50.667
R2093 VDD.n24 VDD.n23 50.667
R2094 VDD.n34 VDD.n33 50.667
R2095 VDD.n37 VDD.n36 50.667
R2096 VDD.n42 VDD.n41 50.667
R2097 VDD.n45 VDD.n44 50.667
R2098 VDD.n48 VDD.n47 50.667
R2099 VDD.n51 VDD.n50 50.667
R2100 VDD.n55 VDD.n54 50.667
R2101 VDD.n58 VDD.n57 50.667
R2102 VDD.n63 VDD.n62 50.667
R2103 VDD.n66 VDD.n65 50.667
R2104 VDD.n69 VDD.n68 50.667
R2105 VDD.n72 VDD.n71 50.667
R2106 VDD.n75 VDD.n74 50.667
R2107 VDD.n79 VDD.n78 50.667
R2108 VDD.n82 VDD.n81 50.667
R2109 VDD.n85 VDD.n84 50.667
R2110 VDD.n90 VDD.n89 50.667
R2111 VDD.n93 VDD.n92 50.667
R2112 VDD.n96 VDD.n95 50.667
R2113 VDD.n101 VDD.n100 50.667
R2114 VDD.n104 VDD.n103 50.667
R2115 VDD.n107 VDD.n106 50.667
R2116 VDD.n110 VDD.n109 50.667
R2117 VDD.n117 VDD.n116 50.667
R2118 VDD.n120 VDD.n119 50.667
R2119 VDD.n125 VDD.n124 50.667
R2120 VDD.n128 VDD.n127 50.667
R2121 VDD.n131 VDD.n130 50.667
R2122 VDD.n134 VDD.n133 50.667
R2123 VDD.n138 VDD.n137 50.667
R2124 VDD.n141 VDD.n140 50.667
R2125 VDD.n146 VDD.n145 50.667
R2126 VDD.n149 VDD.n148 50.667
R2127 VDD.n152 VDD.n151 50.667
R2128 VDD.n155 VDD.n154 50.667
R2129 VDD.n158 VDD.n157 50.667
R2130 VDD.n162 VDD.n161 50.667
R2131 VDD.n165 VDD.n164 50.667
R2132 VDD.n168 VDD.n167 50.667
R2133 VDD.n173 VDD.n172 50.667
R2134 VDD.n176 VDD.n175 50.667
R2135 VDD.n179 VDD.n178 50.667
R2136 VDD.n184 VDD.n183 50.667
R2137 VDD.n187 VDD.n186 50.667
R2138 VDD.n190 VDD.n189 50.667
R2139 VDD.n193 VDD.n192 50.667
R2140 VDD.n200 VDD.n199 50.667
R2141 VDD.n203 VDD.n202 50.667
R2142 VDD.n208 VDD.n207 50.667
R2143 VDD.n211 VDD.n210 50.667
R2144 VDD.n214 VDD.n213 50.667
R2145 VDD.n217 VDD.n216 50.667
R2146 VDD.n221 VDD.n220 50.667
R2147 VDD.n224 VDD.n223 50.667
R2148 VDD.n229 VDD.n228 50.667
R2149 VDD.n232 VDD.n231 50.667
R2150 VDD.n235 VDD.n234 50.667
R2151 VDD.n238 VDD.n237 50.667
R2152 VDD.n241 VDD.n240 50.667
R2153 VDD.n245 VDD.n244 50.667
R2154 VDD.n248 VDD.n247 50.667
R2155 VDD.n251 VDD.n250 50.667
R2156 VDD.n256 VDD.n255 50.667
R2157 VDD.n259 VDD.n258 50.667
R2158 VDD.n262 VDD.n261 50.667
R2159 VDD.n267 VDD.n266 50.667
R2160 VDD.n270 VDD.n269 50.667
R2161 VDD.n273 VDD.n272 50.667
R2162 VDD.n276 VDD.n275 50.667
R2163 VDD.n283 VDD.n282 50.667
R2164 VDD.n286 VDD.n285 50.667
R2165 VDD.n291 VDD.n290 50.667
R2166 VDD.n294 VDD.n293 50.667
R2167 VDD.n297 VDD.n296 50.667
R2168 VDD.n300 VDD.n299 50.667
R2169 VDD.n304 VDD.n303 50.667
R2170 VDD.n307 VDD.n306 50.667
R2171 VDD.n312 VDD.n311 50.667
R2172 VDD.n315 VDD.n314 50.667
R2173 VDD.n318 VDD.n317 50.667
R2174 VDD.n321 VDD.n320 50.667
R2175 VDD.n324 VDD.n323 50.667
R2176 VDD.n328 VDD.n327 50.667
R2177 VDD.n331 VDD.n330 50.667
R2178 VDD.n334 VDD.n333 50.667
R2179 VDD.n339 VDD.n338 50.667
R2180 VDD.n342 VDD.n341 50.667
R2181 VDD.n345 VDD.n344 50.667
R2182 VDD.n350 VDD.n349 50.667
R2183 VDD.n353 VDD.n352 50.667
R2184 VDD.n356 VDD.n355 50.667
R2185 VDD.n359 VDD.n358 50.667
R2186 VDD.n366 VDD.n365 50.667
R2187 VDD.n369 VDD.n368 50.667
R2188 VDD.n374 VDD.n373 50.667
R2189 VDD.n377 VDD.n376 50.667
R2190 VDD.n380 VDD.n379 50.667
R2191 VDD.n383 VDD.n382 50.667
R2192 VDD.n387 VDD.n386 50.667
R2193 VDD.n390 VDD.n389 50.667
R2194 VDD.n395 VDD.n394 50.667
R2195 VDD.n398 VDD.n397 50.667
R2196 VDD.n401 VDD.n400 50.667
R2197 VDD.n404 VDD.n403 50.667
R2198 VDD.n407 VDD.n406 50.667
R2199 VDD.n411 VDD.n410 50.667
R2200 VDD.n414 VDD.n413 50.667
R2201 VDD.n417 VDD.n416 50.667
R2202 VDD.n422 VDD.n421 50.667
R2203 VDD.n425 VDD.n424 50.667
R2204 VDD.n428 VDD.n427 50.667
R2205 VDD.n433 VDD.n432 50.667
R2206 VDD.n436 VDD.n435 50.667
R2207 VDD.n439 VDD.n438 50.667
R2208 VDD.n442 VDD.n441 50.667
R2209 VDD.n449 VDD.n448 50.667
R2210 VDD.n452 VDD.n451 50.667
R2211 VDD.n457 VDD.n456 50.667
R2212 VDD.n460 VDD.n459 50.667
R2213 VDD.n463 VDD.n462 50.667
R2214 VDD.n466 VDD.n465 50.667
R2215 VDD.n470 VDD.n469 50.667
R2216 VDD.n473 VDD.n472 50.667
R2217 VDD.n478 VDD.n477 50.667
R2218 VDD.n481 VDD.n480 50.667
R2219 VDD.n484 VDD.n483 50.667
R2220 VDD.n487 VDD.n486 50.667
R2221 VDD.n490 VDD.n489 50.667
R2222 VDD.n494 VDD.n493 50.667
R2223 VDD.n497 VDD.n496 50.667
R2224 VDD.n500 VDD.n499 50.667
R2225 VDD.n505 VDD.n504 50.667
R2226 VDD.n508 VDD.n507 50.667
R2227 VDD.n511 VDD.n510 50.667
R2228 VDD.n516 VDD.n515 50.667
R2229 VDD.n519 VDD.n518 50.667
R2230 VDD.n522 VDD.n521 50.667
R2231 VDD.n525 VDD.n524 50.667
R2232 VDD.n532 VDD.n531 50.667
R2233 VDD.n535 VDD.n534 50.667
R2234 VDD.n540 VDD.n539 50.667
R2235 VDD.n543 VDD.n542 50.667
R2236 VDD.n546 VDD.n545 50.667
R2237 VDD.n549 VDD.n548 50.667
R2238 VDD.n553 VDD.n552 50.667
R2239 VDD.n556 VDD.n555 50.667
R2240 VDD.n561 VDD.n560 50.667
R2241 VDD.n564 VDD.n563 50.667
R2242 VDD.n567 VDD.n566 50.667
R2243 VDD.n570 VDD.n569 50.667
R2244 VDD.n573 VDD.n572 50.667
R2245 VDD.n577 VDD.n576 50.667
R2246 VDD.n580 VDD.n579 50.667
R2247 VDD.n583 VDD.n582 50.667
R2248 VDD.n588 VDD.n587 50.667
R2249 VDD.n591 VDD.n590 50.667
R2250 VDD.n594 VDD.n593 50.667
R2251 VDD.n599 VDD.n598 50.667
R2252 VDD.n602 VDD.n601 50.667
R2253 VDD.n605 VDD.n604 50.667
R2254 VDD.n608 VDD.n607 50.667
R2255 VDD.n615 VDD.n614 50.667
R2256 VDD.n618 VDD.n617 50.667
R2257 VDD.n623 VDD.n622 50.667
R2258 VDD.n626 VDD.n625 50.667
R2259 VDD.n629 VDD.n628 50.667
R2260 VDD.n632 VDD.n631 50.667
R2261 VDD.n636 VDD.n635 50.667
R2262 VDD.n639 VDD.n638 50.667
R2263 VDD.n644 VDD.n643 50.667
R2264 VDD.n647 VDD.n646 50.667
R2265 VDD.n650 VDD.n649 50.667
R2266 VDD.n653 VDD.n652 50.667
R2267 VDD.n656 VDD.n655 50.667
R2268 VDD.n660 VDD.n659 50.667
R2269 VDD.n663 VDD.n662 50.667
R2270 VDD.n666 VDD.n665 50.667
R2271 VDD.n671 VDD.n670 50.667
R2272 VDD.n674 VDD.n673 50.667
R2273 VDD.n677 VDD.n676 50.667
R2274 VDD.n682 VDD.n681 50.667
R2275 VDD.n685 VDD.n684 50.667
R2276 VDD.n688 VDD.n687 50.667
R2277 VDD.n691 VDD.n690 50.667
R2278 VDD.n698 VDD.n697 50.667
R2279 VDD.n701 VDD.n700 50.667
R2280 VDD.n706 VDD.n705 50.667
R2281 VDD.n709 VDD.n708 50.667
R2282 VDD.n712 VDD.n711 50.667
R2283 VDD.n715 VDD.n714 50.667
R2284 VDD.n719 VDD.n718 50.667
R2285 VDD.n722 VDD.n721 50.667
R2286 VDD.n727 VDD.n726 50.667
R2287 VDD.n730 VDD.n729 50.667
R2288 VDD.n733 VDD.n732 50.667
R2289 VDD.n736 VDD.n735 50.667
R2290 VDD.n739 VDD.n738 50.667
R2291 VDD.n743 VDD.n742 50.667
R2292 VDD.n746 VDD.n745 50.667
R2293 VDD.n749 VDD.n748 50.667
R2294 VDD.n754 VDD.n753 50.667
R2295 VDD.n757 VDD.n756 50.667
R2296 VDD.n760 VDD.n759 50.667
R2297 VDD.n765 VDD.n764 50.667
R2298 VDD.n768 VDD.n767 50.667
R2299 VDD.n771 VDD.n770 50.667
R2300 VDD.n774 VDD.n773 50.667
R2301 VDD.n781 VDD.n780 50.667
R2302 VDD.n784 VDD.n783 50.667
R2303 VDD.n789 VDD.n788 50.667
R2304 VDD.n792 VDD.n791 50.667
R2305 VDD.n795 VDD.n794 50.667
R2306 VDD.n798 VDD.n797 50.667
R2307 VDD.n802 VDD.n801 50.667
R2308 VDD.n805 VDD.n804 50.667
R2309 VDD.n810 VDD.n809 50.667
R2310 VDD.n813 VDD.n812 50.667
R2311 VDD.n816 VDD.n815 50.667
R2312 VDD.n819 VDD.n818 50.667
R2313 VDD.n822 VDD.n821 50.667
R2314 VDD.n826 VDD.n825 50.667
R2315 VDD.n829 VDD.n828 50.667
R2316 VDD.n832 VDD.n831 50.667
R2317 VDD.n837 VDD.n836 50.667
R2318 VDD.n840 VDD.n839 50.667
R2319 VDD.n843 VDD.n842 50.667
R2320 VDD.n848 VDD.n847 50.667
R2321 VDD.n851 VDD.n850 50.667
R2322 VDD.n854 VDD.n853 50.667
R2323 VDD.n857 VDD.n856 50.667
R2324 VDD.n864 VDD.n863 50.667
R2325 VDD.n867 VDD.n866 50.667
R2326 VDD.n872 VDD.n871 50.667
R2327 VDD.n875 VDD.n874 50.667
R2328 VDD.n878 VDD.n877 50.667
R2329 VDD.n881 VDD.n880 50.667
R2330 VDD.n885 VDD.n884 50.667
R2331 VDD.n888 VDD.n887 50.667
R2332 VDD.n893 VDD.n892 50.667
R2333 VDD.n896 VDD.n895 50.667
R2334 VDD.n899 VDD.n898 50.667
R2335 VDD.n902 VDD.n901 50.667
R2336 VDD.n905 VDD.n904 50.667
R2337 VDD.n909 VDD.n908 50.667
R2338 VDD.n912 VDD.n911 50.667
R2339 VDD.n915 VDD.n914 50.667
R2340 VDD.n920 VDD.n919 50.667
R2341 VDD.n923 VDD.n922 50.667
R2342 VDD.n926 VDD.n925 50.667
R2343 VDD.n931 VDD.n930 50.667
R2344 VDD.n934 VDD.n933 50.667
R2345 VDD.n937 VDD.n936 50.667
R2346 VDD.n940 VDD.n939 50.667
R2347 VDD.n947 VDD.n946 50.667
R2348 VDD.n950 VDD.n949 50.667
R2349 VDD.n955 VDD.n954 50.667
R2350 VDD.n958 VDD.n957 50.667
R2351 VDD.n961 VDD.n960 50.667
R2352 VDD.n964 VDD.n963 50.667
R2353 VDD.n968 VDD.n967 50.667
R2354 VDD.n971 VDD.n970 50.667
R2355 VDD.n976 VDD.n975 50.667
R2356 VDD.n979 VDD.n978 50.667
R2357 VDD.n982 VDD.n981 50.667
R2358 VDD.n985 VDD.n984 50.667
R2359 VDD.n988 VDD.n987 50.667
R2360 VDD.n992 VDD.n991 50.667
R2361 VDD.n995 VDD.n994 50.667
R2362 VDD.n998 VDD.n997 50.667
R2363 VDD.n1003 VDD.n1002 50.667
R2364 VDD.n1006 VDD.n1005 50.667
R2365 VDD.n1009 VDD.n1008 50.667
R2366 VDD.n1014 VDD.n1013 50.667
R2367 VDD.n1017 VDD.n1016 50.667
R2368 VDD.n1020 VDD.n1019 50.667
R2369 VDD.n1023 VDD.n1022 50.667
R2370 VDD.n1030 VDD.n1029 50.667
R2371 VDD.n1033 VDD.n1032 50.667
R2372 VDD.n1038 VDD.n1037 50.667
R2373 VDD.n1041 VDD.n1040 50.667
R2374 VDD.n1044 VDD.n1043 50.667
R2375 VDD.n1047 VDD.n1046 50.667
R2376 VDD.n1051 VDD.n1050 50.667
R2377 VDD.n1054 VDD.n1053 50.667
R2378 VDD.n1059 VDD.n1058 50.667
R2379 VDD.n1062 VDD.n1061 50.667
R2380 VDD.n1065 VDD.n1064 50.667
R2381 VDD.n1068 VDD.n1067 50.667
R2382 VDD.n1071 VDD.n1070 50.667
R2383 VDD.n1075 VDD.n1074 50.667
R2384 VDD.n1078 VDD.n1077 50.667
R2385 VDD.n1081 VDD.n1080 50.667
R2386 VDD.n1086 VDD.n1085 50.667
R2387 VDD.n1089 VDD.n1088 50.667
R2388 VDD.n1092 VDD.n1091 50.667
R2389 VDD.n1097 VDD.n1096 50.667
R2390 VDD.n1100 VDD.n1099 50.667
R2391 VDD.n1103 VDD.n1102 50.667
R2392 VDD.n1106 VDD.n1105 50.667
R2393 VDD.n1113 VDD.n1112 50.667
R2394 VDD.n1116 VDD.n1115 50.667
R2395 VDD.n1121 VDD.n1120 50.667
R2396 VDD.n1124 VDD.n1123 50.667
R2397 VDD.n1127 VDD.n1126 50.667
R2398 VDD.n1130 VDD.n1129 50.667
R2399 VDD.n1134 VDD.n1133 50.667
R2400 VDD.n1137 VDD.n1136 50.667
R2401 VDD.n1142 VDD.n1141 50.667
R2402 VDD.n1145 VDD.n1144 50.667
R2403 VDD.n1148 VDD.n1147 50.667
R2404 VDD.n1151 VDD.n1150 50.667
R2405 VDD.n1154 VDD.n1153 50.667
R2406 VDD.n1630 VDD.n1629 50.667
R2407 VDD.n1577 VDD.t10 41.554
R2408 VDD.n1577 VDD.t12 41.554
R2409 VDD.n1494 VDD.t144 41.554
R2410 VDD.n1494 VDD.t238 41.554
R2411 VDD.n1411 VDD.t29 41.554
R2412 VDD.n1411 VDD.t21 41.554
R2413 VDD.n1328 VDD.t75 41.554
R2414 VDD.n1328 VDD.t17 41.554
R2415 VDD.n1245 VDD.t42 41.554
R2416 VDD.n1245 VDD.t57 41.554
R2417 VDD.n1162 VDD.t37 41.554
R2418 VDD.n1162 VDD.t123 41.554
R2419 VDD.n86 VDD.t127 41.554
R2420 VDD.n86 VDD.t136 41.554
R2421 VDD.n169 VDD.t99 41.554
R2422 VDD.n169 VDD.t118 41.554
R2423 VDD.n252 VDD.t130 41.554
R2424 VDD.n252 VDD.t50 41.554
R2425 VDD.n335 VDD.t143 41.554
R2426 VDD.n335 VDD.t97 41.554
R2427 VDD.n418 VDD.t141 41.554
R2428 VDD.n418 VDD.t46 41.554
R2429 VDD.n501 VDD.t166 41.554
R2430 VDD.n501 VDD.t172 41.554
R2431 VDD.n584 VDD.t148 41.554
R2432 VDD.n584 VDD.t35 41.554
R2433 VDD.n667 VDD.t233 41.554
R2434 VDD.n667 VDD.t72 41.554
R2435 VDD.n750 VDD.t120 41.554
R2436 VDD.n750 VDD.t61 41.554
R2437 VDD.n833 VDD.t1 41.554
R2438 VDD.n833 VDD.t229 41.554
R2439 VDD.n916 VDD.t153 41.554
R2440 VDD.n916 VDD.t161 41.554
R2441 VDD.n999 VDD.t182 41.554
R2442 VDD.n999 VDD.t231 41.554
R2443 VDD.n1082 VDD.t104 41.554
R2444 VDD.n1082 VDD.t54 41.554
R2445 VDD.n0 VDD.t110 41.554
R2446 VDD.n0 VDD.t2 41.554
R2447 VDD.n1655 VDD.n1654 40.334
R2448 VDD.n1566 VDD.t71 30.569
R2449 VDD.n1483 VDD.t7 30.569
R2450 VDD.n1400 VDD.t24 30.569
R2451 VDD.n1317 VDD.t28 30.569
R2452 VDD.n1234 VDD.t165 30.569
R2453 VDD.n16 VDD.t119 30.569
R2454 VDD.n97 VDD.t155 30.569
R2455 VDD.n180 VDD.t138 30.569
R2456 VDD.n263 VDD.t227 30.569
R2457 VDD.n346 VDD.t150 30.569
R2458 VDD.n429 VDD.t39 30.569
R2459 VDD.n512 VDD.t125 30.569
R2460 VDD.n595 VDD.t145 30.569
R2461 VDD.n678 VDD.t152 30.569
R2462 VDD.n761 VDD.t95 30.569
R2463 VDD.n844 VDD.t48 30.569
R2464 VDD.n927 VDD.t162 30.569
R2465 VDD.n1010 VDD.t68 30.569
R2466 VDD.n1093 VDD.t160 30.569
R2467 VDD.n1107 VDD.t157 29.315
R2468 VDD.n1024 VDD.t22 29.315
R2469 VDD.n941 VDD.t5 29.315
R2470 VDD.n858 VDD.t149 29.315
R2471 VDD.n775 VDD.t108 29.315
R2472 VDD.n692 VDD.t16 29.315
R2473 VDD.n609 VDD.t79 29.315
R2474 VDD.n526 VDD.t121 29.315
R2475 VDD.n443 VDD.t115 29.315
R2476 VDD.n360 VDD.t106 29.315
R2477 VDD.n277 VDD.t92 29.315
R2478 VDD.n194 VDD.t174 29.315
R2479 VDD.n111 VDD.t90 29.315
R2480 VDD.n28 VDD.t117 29.315
R2481 VDD.n1218 VDD.t131 29.315
R2482 VDD.n1301 VDD.t158 29.315
R2483 VDD.n1384 VDD.t27 29.315
R2484 VDD.n1467 VDD.t19 29.315
R2485 VDD.n1550 VDD.t232 29.315
R2486 VDD.n1643 VDD.t47 29.315
R2487 VDD.n1652 VDD.t4 29.055
R2488 VDD.n21 VDD.n20 28.517
R2489 VDD.n1567 VDD.n1566 27.22
R2490 VDD.n1484 VDD.n1483 27.22
R2491 VDD.n1401 VDD.n1400 27.22
R2492 VDD.n1318 VDD.n1317 27.22
R2493 VDD.n1235 VDD.n1234 27.22
R2494 VDD.n19 VDD.n16 27.22
R2495 VDD.n98 VDD.n97 27.22
R2496 VDD.n181 VDD.n180 27.22
R2497 VDD.n264 VDD.n263 27.22
R2498 VDD.n347 VDD.n346 27.22
R2499 VDD.n430 VDD.n429 27.22
R2500 VDD.n513 VDD.n512 27.22
R2501 VDD.n596 VDD.n595 27.22
R2502 VDD.n679 VDD.n678 27.22
R2503 VDD.n762 VDD.n761 27.22
R2504 VDD.n845 VDD.n844 27.22
R2505 VDD.n928 VDD.n927 27.22
R2506 VDD.n1011 VDD.n1010 27.22
R2507 VDD.n1094 VDD.n1093 27.22
R2508 VDD.n1654 VDD.n1651 25.815
R2509 VDD.n1578 VDD.n1577 22.842
R2510 VDD.n1495 VDD.n1494 22.842
R2511 VDD.n1412 VDD.n1411 22.842
R2512 VDD.n1329 VDD.n1328 22.842
R2513 VDD.n1246 VDD.n1245 22.842
R2514 VDD.n1163 VDD.n1162 22.842
R2515 VDD.n87 VDD.n86 22.842
R2516 VDD.n170 VDD.n169 22.842
R2517 VDD.n253 VDD.n252 22.842
R2518 VDD.n336 VDD.n335 22.842
R2519 VDD.n419 VDD.n418 22.842
R2520 VDD.n502 VDD.n501 22.842
R2521 VDD.n585 VDD.n584 22.842
R2522 VDD.n668 VDD.n667 22.842
R2523 VDD.n751 VDD.n750 22.842
R2524 VDD.n834 VDD.n833 22.842
R2525 VDD.n917 VDD.n916 22.842
R2526 VDD.n1000 VDD.n999 22.842
R2527 VDD.n1083 VDD.n1082 22.842
R2528 VDD.n10 VDD.n0 22.842
R2529 VDD.n1635 VDD.n1632 21.896
R2530 VDD.n1543 VDD.n1542 21.896
R2531 VDD.n1460 VDD.n1459 21.896
R2532 VDD.n1377 VDD.n1376 21.896
R2533 VDD.n1294 VDD.n1293 21.896
R2534 VDD.n1211 VDD.n1210 21.896
R2535 VDD.n39 VDD.n38 21.896
R2536 VDD.n122 VDD.n121 21.896
R2537 VDD.n205 VDD.n204 21.896
R2538 VDD.n288 VDD.n287 21.896
R2539 VDD.n371 VDD.n370 21.896
R2540 VDD.n454 VDD.n453 21.896
R2541 VDD.n537 VDD.n536 21.896
R2542 VDD.n620 VDD.n619 21.896
R2543 VDD.n703 VDD.n702 21.896
R2544 VDD.n786 VDD.n785 21.896
R2545 VDD.n869 VDD.n868 21.896
R2546 VDD.n952 VDD.n951 21.896
R2547 VDD.n1035 VDD.n1034 21.896
R2548 VDD.n1118 VDD.n1117 21.896
R2549 VDD.n1605 VDD.n1604 20.254
R2550 VDD.n1522 VDD.n1521 20.254
R2551 VDD.n1439 VDD.n1438 20.254
R2552 VDD.n1356 VDD.n1355 20.254
R2553 VDD.n1273 VDD.n1272 20.254
R2554 VDD.n1190 VDD.n1189 20.254
R2555 VDD.n60 VDD.n59 20.254
R2556 VDD.n143 VDD.n142 20.254
R2557 VDD.n226 VDD.n225 20.254
R2558 VDD.n309 VDD.n308 20.254
R2559 VDD.n392 VDD.n391 20.254
R2560 VDD.n475 VDD.n474 20.254
R2561 VDD.n558 VDD.n557 20.254
R2562 VDD.n641 VDD.n640 20.254
R2563 VDD.n724 VDD.n723 20.254
R2564 VDD.n807 VDD.n806 20.254
R2565 VDD.n890 VDD.n889 20.254
R2566 VDD.n973 VDD.n972 20.254
R2567 VDD.n1056 VDD.n1055 20.254
R2568 VDD.n1139 VDD.n1138 20.254
R2569 VDD.n1639 VDD.n1637 15.167
R2570 VDD.n7 VDD.n5 15.167
R2571 VDD.n9 VDD.n7 15.167
R2572 VDD.n14 VDD.n12 15.167
R2573 VDD.n1630 VDD.n14 15.167
R2574 VDD.n1650 VDD.n1648 15.167
R2575 VDD.n1648 VDD.n1646 15.167
R2576 VDD.n12 VDD.n10 14.837
R2577 VDD.n19 VDD.n18 13.683
R2578 VDD.n1651 VDD.n1650 13.683
R2579 VDD.n1635 VDD.n1634 13.024
R2580 VDD.n5 VDD.n3 12.035
R2581 VDD.n1640 VDD.n1631 7.5
R2582 VDD.n1644 VDD.n1643 7.5
R2583 VDD.n1553 VDD.n1552 7.5
R2584 VDD.n1551 VDD.n1550 7.5
R2585 VDD.n1470 VDD.n1469 7.5
R2586 VDD.n1468 VDD.n1467 7.5
R2587 VDD.n1387 VDD.n1386 7.5
R2588 VDD.n1385 VDD.n1384 7.5
R2589 VDD.n1304 VDD.n1303 7.5
R2590 VDD.n1302 VDD.n1301 7.5
R2591 VDD.n1221 VDD.n1220 7.5
R2592 VDD.n1219 VDD.n1218 7.5
R2593 VDD.n31 VDD.n30 7.5
R2594 VDD.n29 VDD.n28 7.5
R2595 VDD.n114 VDD.n113 7.5
R2596 VDD.n112 VDD.n111 7.5
R2597 VDD.n197 VDD.n196 7.5
R2598 VDD.n195 VDD.n194 7.5
R2599 VDD.n280 VDD.n279 7.5
R2600 VDD.n278 VDD.n277 7.5
R2601 VDD.n363 VDD.n362 7.5
R2602 VDD.n361 VDD.n360 7.5
R2603 VDD.n446 VDD.n445 7.5
R2604 VDD.n444 VDD.n443 7.5
R2605 VDD.n529 VDD.n528 7.5
R2606 VDD.n527 VDD.n526 7.5
R2607 VDD.n612 VDD.n611 7.5
R2608 VDD.n610 VDD.n609 7.5
R2609 VDD.n695 VDD.n694 7.5
R2610 VDD.n693 VDD.n692 7.5
R2611 VDD.n778 VDD.n777 7.5
R2612 VDD.n776 VDD.n775 7.5
R2613 VDD.n861 VDD.n860 7.5
R2614 VDD.n859 VDD.n858 7.5
R2615 VDD.n944 VDD.n943 7.5
R2616 VDD.n942 VDD.n941 7.5
R2617 VDD.n1027 VDD.n1026 7.5
R2618 VDD.n1025 VDD.n1024 7.5
R2619 VDD.n1110 VDD.n1109 7.5
R2620 VDD.n1108 VDD.n1107 7.5
R2621 VDD.n1165 VDD.n1164 7.147
R2622 VDD.n1168 VDD.n1167 7.147
R2623 VDD.n1171 VDD.n1170 7.147
R2624 VDD.n1175 VDD.n1174 7.147
R2625 VDD.n1178 VDD.n1177 7.147
R2626 VDD.n1181 VDD.n1180 7.147
R2627 VDD.n1184 VDD.n1183 7.147
R2628 VDD.n1187 VDD.n1186 7.147
R2629 VDD.n1192 VDD.n1191 7.147
R2630 VDD.n1195 VDD.n1194 7.147
R2631 VDD.n1199 VDD.n1198 7.147
R2632 VDD.n1202 VDD.n1201 7.147
R2633 VDD.n1205 VDD.n1204 7.147
R2634 VDD.n1208 VDD.n1207 7.147
R2635 VDD.n1213 VDD.n1212 7.147
R2636 VDD.n1216 VDD.n1215 7.147
R2637 VDD.n1223 VDD.n1222 7.147
R2638 VDD.n1226 VDD.n1225 7.147
R2639 VDD.n1229 VDD.n1228 7.147
R2640 VDD.n1232 VDD.n1231 7.147
R2641 VDD.n1237 VDD.n1236 7.147
R2642 VDD.n1240 VDD.n1239 7.147
R2643 VDD.n1243 VDD.n1242 7.147
R2644 VDD.n1248 VDD.n1247 7.147
R2645 VDD.n1251 VDD.n1250 7.147
R2646 VDD.n1254 VDD.n1253 7.147
R2647 VDD.n1258 VDD.n1257 7.147
R2648 VDD.n1261 VDD.n1260 7.147
R2649 VDD.n1264 VDD.n1263 7.147
R2650 VDD.n1267 VDD.n1266 7.147
R2651 VDD.n1270 VDD.n1269 7.147
R2652 VDD.n1275 VDD.n1274 7.147
R2653 VDD.n1278 VDD.n1277 7.147
R2654 VDD.n1282 VDD.n1281 7.147
R2655 VDD.n1285 VDD.n1284 7.147
R2656 VDD.n1288 VDD.n1287 7.147
R2657 VDD.n1291 VDD.n1290 7.147
R2658 VDD.n1296 VDD.n1295 7.147
R2659 VDD.n1299 VDD.n1298 7.147
R2660 VDD.n1306 VDD.n1305 7.147
R2661 VDD.n1309 VDD.n1308 7.147
R2662 VDD.n1312 VDD.n1311 7.147
R2663 VDD.n1315 VDD.n1314 7.147
R2664 VDD.n1320 VDD.n1319 7.147
R2665 VDD.n1323 VDD.n1322 7.147
R2666 VDD.n1326 VDD.n1325 7.147
R2667 VDD.n1331 VDD.n1330 7.147
R2668 VDD.n1334 VDD.n1333 7.147
R2669 VDD.n1337 VDD.n1336 7.147
R2670 VDD.n1341 VDD.n1340 7.147
R2671 VDD.n1344 VDD.n1343 7.147
R2672 VDD.n1347 VDD.n1346 7.147
R2673 VDD.n1350 VDD.n1349 7.147
R2674 VDD.n1353 VDD.n1352 7.147
R2675 VDD.n1358 VDD.n1357 7.147
R2676 VDD.n1361 VDD.n1360 7.147
R2677 VDD.n1365 VDD.n1364 7.147
R2678 VDD.n1368 VDD.n1367 7.147
R2679 VDD.n1371 VDD.n1370 7.147
R2680 VDD.n1374 VDD.n1373 7.147
R2681 VDD.n1379 VDD.n1378 7.147
R2682 VDD.n1382 VDD.n1381 7.147
R2683 VDD.n1389 VDD.n1388 7.147
R2684 VDD.n1392 VDD.n1391 7.147
R2685 VDD.n1395 VDD.n1394 7.147
R2686 VDD.n1398 VDD.n1397 7.147
R2687 VDD.n1403 VDD.n1402 7.147
R2688 VDD.n1406 VDD.n1405 7.147
R2689 VDD.n1409 VDD.n1408 7.147
R2690 VDD.n1414 VDD.n1413 7.147
R2691 VDD.n1417 VDD.n1416 7.147
R2692 VDD.n1420 VDD.n1419 7.147
R2693 VDD.n1424 VDD.n1423 7.147
R2694 VDD.n1427 VDD.n1426 7.147
R2695 VDD.n1430 VDD.n1429 7.147
R2696 VDD.n1433 VDD.n1432 7.147
R2697 VDD.n1436 VDD.n1435 7.147
R2698 VDD.n1441 VDD.n1440 7.147
R2699 VDD.n1444 VDD.n1443 7.147
R2700 VDD.n1448 VDD.n1447 7.147
R2701 VDD.n1451 VDD.n1450 7.147
R2702 VDD.n1454 VDD.n1453 7.147
R2703 VDD.n1457 VDD.n1456 7.147
R2704 VDD.n1462 VDD.n1461 7.147
R2705 VDD.n1465 VDD.n1464 7.147
R2706 VDD.n1472 VDD.n1471 7.147
R2707 VDD.n1475 VDD.n1474 7.147
R2708 VDD.n1478 VDD.n1477 7.147
R2709 VDD.n1481 VDD.n1480 7.147
R2710 VDD.n1486 VDD.n1485 7.147
R2711 VDD.n1489 VDD.n1488 7.147
R2712 VDD.n1492 VDD.n1491 7.147
R2713 VDD.n1497 VDD.n1496 7.147
R2714 VDD.n1500 VDD.n1499 7.147
R2715 VDD.n1503 VDD.n1502 7.147
R2716 VDD.n1507 VDD.n1506 7.147
R2717 VDD.n1510 VDD.n1509 7.147
R2718 VDD.n1513 VDD.n1512 7.147
R2719 VDD.n1516 VDD.n1515 7.147
R2720 VDD.n1519 VDD.n1518 7.147
R2721 VDD.n1524 VDD.n1523 7.147
R2722 VDD.n1527 VDD.n1526 7.147
R2723 VDD.n1531 VDD.n1530 7.147
R2724 VDD.n1534 VDD.n1533 7.147
R2725 VDD.n1537 VDD.n1536 7.147
R2726 VDD.n1540 VDD.n1539 7.147
R2727 VDD.n1545 VDD.n1544 7.147
R2728 VDD.n1548 VDD.n1547 7.147
R2729 VDD.n1555 VDD.n1554 7.147
R2730 VDD.n1558 VDD.n1557 7.147
R2731 VDD.n1561 VDD.n1560 7.147
R2732 VDD.n1564 VDD.n1563 7.147
R2733 VDD.n1569 VDD.n1568 7.147
R2734 VDD.n1572 VDD.n1571 7.147
R2735 VDD.n1575 VDD.n1574 7.147
R2736 VDD.n1580 VDD.n1579 7.147
R2737 VDD.n1583 VDD.n1582 7.147
R2738 VDD.n1586 VDD.n1585 7.147
R2739 VDD.n1590 VDD.n1589 7.147
R2740 VDD.n1593 VDD.n1592 7.147
R2741 VDD.n1596 VDD.n1595 7.147
R2742 VDD.n1599 VDD.n1598 7.147
R2743 VDD.n1602 VDD.n1601 7.147
R2744 VDD.n1607 VDD.n1606 7.147
R2745 VDD.n1610 VDD.n1609 7.147
R2746 VDD.n1614 VDD.n1613 7.147
R2747 VDD.n1617 VDD.n1616 7.147
R2748 VDD.n1620 VDD.n1619 7.147
R2749 VDD.n1634 VDD.n1633 7.147
R2750 VDD.n1637 VDD.n1636 7.147
R2751 VDD.n1639 VDD.n1638 7.147
R2752 VDD.n1642 VDD.n1641 7.147
R2753 VDD.n26 VDD.n25 7.147
R2754 VDD.n23 VDD.n22 7.147
R2755 VDD.n18 VDD.n17 7.147
R2756 VDD.n33 VDD.n32 7.147
R2757 VDD.n109 VDD.n108 7.147
R2758 VDD.n106 VDD.n105 7.147
R2759 VDD.n103 VDD.n102 7.147
R2760 VDD.n100 VDD.n99 7.147
R2761 VDD.n95 VDD.n94 7.147
R2762 VDD.n92 VDD.n91 7.147
R2763 VDD.n89 VDD.n88 7.147
R2764 VDD.n84 VDD.n83 7.147
R2765 VDD.n81 VDD.n80 7.147
R2766 VDD.n78 VDD.n77 7.147
R2767 VDD.n74 VDD.n73 7.147
R2768 VDD.n71 VDD.n70 7.147
R2769 VDD.n68 VDD.n67 7.147
R2770 VDD.n65 VDD.n64 7.147
R2771 VDD.n62 VDD.n61 7.147
R2772 VDD.n57 VDD.n56 7.147
R2773 VDD.n54 VDD.n53 7.147
R2774 VDD.n50 VDD.n49 7.147
R2775 VDD.n47 VDD.n46 7.147
R2776 VDD.n44 VDD.n43 7.147
R2777 VDD.n41 VDD.n40 7.147
R2778 VDD.n36 VDD.n35 7.147
R2779 VDD.n116 VDD.n115 7.147
R2780 VDD.n192 VDD.n191 7.147
R2781 VDD.n189 VDD.n188 7.147
R2782 VDD.n186 VDD.n185 7.147
R2783 VDD.n183 VDD.n182 7.147
R2784 VDD.n178 VDD.n177 7.147
R2785 VDD.n175 VDD.n174 7.147
R2786 VDD.n172 VDD.n171 7.147
R2787 VDD.n167 VDD.n166 7.147
R2788 VDD.n164 VDD.n163 7.147
R2789 VDD.n161 VDD.n160 7.147
R2790 VDD.n157 VDD.n156 7.147
R2791 VDD.n154 VDD.n153 7.147
R2792 VDD.n151 VDD.n150 7.147
R2793 VDD.n148 VDD.n147 7.147
R2794 VDD.n145 VDD.n144 7.147
R2795 VDD.n140 VDD.n139 7.147
R2796 VDD.n137 VDD.n136 7.147
R2797 VDD.n133 VDD.n132 7.147
R2798 VDD.n130 VDD.n129 7.147
R2799 VDD.n127 VDD.n126 7.147
R2800 VDD.n124 VDD.n123 7.147
R2801 VDD.n119 VDD.n118 7.147
R2802 VDD.n199 VDD.n198 7.147
R2803 VDD.n275 VDD.n274 7.147
R2804 VDD.n272 VDD.n271 7.147
R2805 VDD.n269 VDD.n268 7.147
R2806 VDD.n266 VDD.n265 7.147
R2807 VDD.n261 VDD.n260 7.147
R2808 VDD.n258 VDD.n257 7.147
R2809 VDD.n255 VDD.n254 7.147
R2810 VDD.n250 VDD.n249 7.147
R2811 VDD.n247 VDD.n246 7.147
R2812 VDD.n244 VDD.n243 7.147
R2813 VDD.n240 VDD.n239 7.147
R2814 VDD.n237 VDD.n236 7.147
R2815 VDD.n234 VDD.n233 7.147
R2816 VDD.n231 VDD.n230 7.147
R2817 VDD.n228 VDD.n227 7.147
R2818 VDD.n223 VDD.n222 7.147
R2819 VDD.n220 VDD.n219 7.147
R2820 VDD.n216 VDD.n215 7.147
R2821 VDD.n213 VDD.n212 7.147
R2822 VDD.n210 VDD.n209 7.147
R2823 VDD.n207 VDD.n206 7.147
R2824 VDD.n202 VDD.n201 7.147
R2825 VDD.n282 VDD.n281 7.147
R2826 VDD.n358 VDD.n357 7.147
R2827 VDD.n355 VDD.n354 7.147
R2828 VDD.n352 VDD.n351 7.147
R2829 VDD.n349 VDD.n348 7.147
R2830 VDD.n344 VDD.n343 7.147
R2831 VDD.n341 VDD.n340 7.147
R2832 VDD.n338 VDD.n337 7.147
R2833 VDD.n333 VDD.n332 7.147
R2834 VDD.n330 VDD.n329 7.147
R2835 VDD.n327 VDD.n326 7.147
R2836 VDD.n323 VDD.n322 7.147
R2837 VDD.n320 VDD.n319 7.147
R2838 VDD.n317 VDD.n316 7.147
R2839 VDD.n314 VDD.n313 7.147
R2840 VDD.n311 VDD.n310 7.147
R2841 VDD.n306 VDD.n305 7.147
R2842 VDD.n303 VDD.n302 7.147
R2843 VDD.n299 VDD.n298 7.147
R2844 VDD.n296 VDD.n295 7.147
R2845 VDD.n293 VDD.n292 7.147
R2846 VDD.n290 VDD.n289 7.147
R2847 VDD.n285 VDD.n284 7.147
R2848 VDD.n365 VDD.n364 7.147
R2849 VDD.n441 VDD.n440 7.147
R2850 VDD.n438 VDD.n437 7.147
R2851 VDD.n435 VDD.n434 7.147
R2852 VDD.n432 VDD.n431 7.147
R2853 VDD.n427 VDD.n426 7.147
R2854 VDD.n424 VDD.n423 7.147
R2855 VDD.n421 VDD.n420 7.147
R2856 VDD.n416 VDD.n415 7.147
R2857 VDD.n413 VDD.n412 7.147
R2858 VDD.n410 VDD.n409 7.147
R2859 VDD.n406 VDD.n405 7.147
R2860 VDD.n403 VDD.n402 7.147
R2861 VDD.n400 VDD.n399 7.147
R2862 VDD.n397 VDD.n396 7.147
R2863 VDD.n394 VDD.n393 7.147
R2864 VDD.n389 VDD.n388 7.147
R2865 VDD.n386 VDD.n385 7.147
R2866 VDD.n382 VDD.n381 7.147
R2867 VDD.n379 VDD.n378 7.147
R2868 VDD.n376 VDD.n375 7.147
R2869 VDD.n373 VDD.n372 7.147
R2870 VDD.n368 VDD.n367 7.147
R2871 VDD.n448 VDD.n447 7.147
R2872 VDD.n524 VDD.n523 7.147
R2873 VDD.n521 VDD.n520 7.147
R2874 VDD.n518 VDD.n517 7.147
R2875 VDD.n515 VDD.n514 7.147
R2876 VDD.n510 VDD.n509 7.147
R2877 VDD.n507 VDD.n506 7.147
R2878 VDD.n504 VDD.n503 7.147
R2879 VDD.n499 VDD.n498 7.147
R2880 VDD.n496 VDD.n495 7.147
R2881 VDD.n493 VDD.n492 7.147
R2882 VDD.n489 VDD.n488 7.147
R2883 VDD.n486 VDD.n485 7.147
R2884 VDD.n483 VDD.n482 7.147
R2885 VDD.n480 VDD.n479 7.147
R2886 VDD.n477 VDD.n476 7.147
R2887 VDD.n472 VDD.n471 7.147
R2888 VDD.n469 VDD.n468 7.147
R2889 VDD.n465 VDD.n464 7.147
R2890 VDD.n462 VDD.n461 7.147
R2891 VDD.n459 VDD.n458 7.147
R2892 VDD.n456 VDD.n455 7.147
R2893 VDD.n451 VDD.n450 7.147
R2894 VDD.n531 VDD.n530 7.147
R2895 VDD.n607 VDD.n606 7.147
R2896 VDD.n604 VDD.n603 7.147
R2897 VDD.n601 VDD.n600 7.147
R2898 VDD.n598 VDD.n597 7.147
R2899 VDD.n593 VDD.n592 7.147
R2900 VDD.n590 VDD.n589 7.147
R2901 VDD.n587 VDD.n586 7.147
R2902 VDD.n582 VDD.n581 7.147
R2903 VDD.n579 VDD.n578 7.147
R2904 VDD.n576 VDD.n575 7.147
R2905 VDD.n572 VDD.n571 7.147
R2906 VDD.n569 VDD.n568 7.147
R2907 VDD.n566 VDD.n565 7.147
R2908 VDD.n563 VDD.n562 7.147
R2909 VDD.n560 VDD.n559 7.147
R2910 VDD.n555 VDD.n554 7.147
R2911 VDD.n552 VDD.n551 7.147
R2912 VDD.n548 VDD.n547 7.147
R2913 VDD.n545 VDD.n544 7.147
R2914 VDD.n542 VDD.n541 7.147
R2915 VDD.n539 VDD.n538 7.147
R2916 VDD.n534 VDD.n533 7.147
R2917 VDD.n614 VDD.n613 7.147
R2918 VDD.n690 VDD.n689 7.147
R2919 VDD.n687 VDD.n686 7.147
R2920 VDD.n684 VDD.n683 7.147
R2921 VDD.n681 VDD.n680 7.147
R2922 VDD.n676 VDD.n675 7.147
R2923 VDD.n673 VDD.n672 7.147
R2924 VDD.n670 VDD.n669 7.147
R2925 VDD.n665 VDD.n664 7.147
R2926 VDD.n662 VDD.n661 7.147
R2927 VDD.n659 VDD.n658 7.147
R2928 VDD.n655 VDD.n654 7.147
R2929 VDD.n652 VDD.n651 7.147
R2930 VDD.n649 VDD.n648 7.147
R2931 VDD.n646 VDD.n645 7.147
R2932 VDD.n643 VDD.n642 7.147
R2933 VDD.n638 VDD.n637 7.147
R2934 VDD.n635 VDD.n634 7.147
R2935 VDD.n631 VDD.n630 7.147
R2936 VDD.n628 VDD.n627 7.147
R2937 VDD.n625 VDD.n624 7.147
R2938 VDD.n622 VDD.n621 7.147
R2939 VDD.n617 VDD.n616 7.147
R2940 VDD.n697 VDD.n696 7.147
R2941 VDD.n773 VDD.n772 7.147
R2942 VDD.n770 VDD.n769 7.147
R2943 VDD.n767 VDD.n766 7.147
R2944 VDD.n764 VDD.n763 7.147
R2945 VDD.n759 VDD.n758 7.147
R2946 VDD.n756 VDD.n755 7.147
R2947 VDD.n753 VDD.n752 7.147
R2948 VDD.n748 VDD.n747 7.147
R2949 VDD.n745 VDD.n744 7.147
R2950 VDD.n742 VDD.n741 7.147
R2951 VDD.n738 VDD.n737 7.147
R2952 VDD.n735 VDD.n734 7.147
R2953 VDD.n732 VDD.n731 7.147
R2954 VDD.n729 VDD.n728 7.147
R2955 VDD.n726 VDD.n725 7.147
R2956 VDD.n721 VDD.n720 7.147
R2957 VDD.n718 VDD.n717 7.147
R2958 VDD.n714 VDD.n713 7.147
R2959 VDD.n711 VDD.n710 7.147
R2960 VDD.n708 VDD.n707 7.147
R2961 VDD.n705 VDD.n704 7.147
R2962 VDD.n700 VDD.n699 7.147
R2963 VDD.n780 VDD.n779 7.147
R2964 VDD.n856 VDD.n855 7.147
R2965 VDD.n853 VDD.n852 7.147
R2966 VDD.n850 VDD.n849 7.147
R2967 VDD.n847 VDD.n846 7.147
R2968 VDD.n842 VDD.n841 7.147
R2969 VDD.n839 VDD.n838 7.147
R2970 VDD.n836 VDD.n835 7.147
R2971 VDD.n831 VDD.n830 7.147
R2972 VDD.n828 VDD.n827 7.147
R2973 VDD.n825 VDD.n824 7.147
R2974 VDD.n821 VDD.n820 7.147
R2975 VDD.n818 VDD.n817 7.147
R2976 VDD.n815 VDD.n814 7.147
R2977 VDD.n812 VDD.n811 7.147
R2978 VDD.n809 VDD.n808 7.147
R2979 VDD.n804 VDD.n803 7.147
R2980 VDD.n801 VDD.n800 7.147
R2981 VDD.n797 VDD.n796 7.147
R2982 VDD.n794 VDD.n793 7.147
R2983 VDD.n791 VDD.n790 7.147
R2984 VDD.n788 VDD.n787 7.147
R2985 VDD.n783 VDD.n782 7.147
R2986 VDD.n863 VDD.n862 7.147
R2987 VDD.n939 VDD.n938 7.147
R2988 VDD.n936 VDD.n935 7.147
R2989 VDD.n933 VDD.n932 7.147
R2990 VDD.n930 VDD.n929 7.147
R2991 VDD.n925 VDD.n924 7.147
R2992 VDD.n922 VDD.n921 7.147
R2993 VDD.n919 VDD.n918 7.147
R2994 VDD.n914 VDD.n913 7.147
R2995 VDD.n911 VDD.n910 7.147
R2996 VDD.n908 VDD.n907 7.147
R2997 VDD.n904 VDD.n903 7.147
R2998 VDD.n901 VDD.n900 7.147
R2999 VDD.n898 VDD.n897 7.147
R3000 VDD.n895 VDD.n894 7.147
R3001 VDD.n892 VDD.n891 7.147
R3002 VDD.n887 VDD.n886 7.147
R3003 VDD.n884 VDD.n883 7.147
R3004 VDD.n880 VDD.n879 7.147
R3005 VDD.n877 VDD.n876 7.147
R3006 VDD.n874 VDD.n873 7.147
R3007 VDD.n871 VDD.n870 7.147
R3008 VDD.n866 VDD.n865 7.147
R3009 VDD.n946 VDD.n945 7.147
R3010 VDD.n1022 VDD.n1021 7.147
R3011 VDD.n1019 VDD.n1018 7.147
R3012 VDD.n1016 VDD.n1015 7.147
R3013 VDD.n1013 VDD.n1012 7.147
R3014 VDD.n1008 VDD.n1007 7.147
R3015 VDD.n1005 VDD.n1004 7.147
R3016 VDD.n1002 VDD.n1001 7.147
R3017 VDD.n997 VDD.n996 7.147
R3018 VDD.n994 VDD.n993 7.147
R3019 VDD.n991 VDD.n990 7.147
R3020 VDD.n987 VDD.n986 7.147
R3021 VDD.n984 VDD.n983 7.147
R3022 VDD.n981 VDD.n980 7.147
R3023 VDD.n978 VDD.n977 7.147
R3024 VDD.n975 VDD.n974 7.147
R3025 VDD.n970 VDD.n969 7.147
R3026 VDD.n967 VDD.n966 7.147
R3027 VDD.n963 VDD.n962 7.147
R3028 VDD.n960 VDD.n959 7.147
R3029 VDD.n957 VDD.n956 7.147
R3030 VDD.n954 VDD.n953 7.147
R3031 VDD.n949 VDD.n948 7.147
R3032 VDD.n1029 VDD.n1028 7.147
R3033 VDD.n1105 VDD.n1104 7.147
R3034 VDD.n1102 VDD.n1101 7.147
R3035 VDD.n1099 VDD.n1098 7.147
R3036 VDD.n1096 VDD.n1095 7.147
R3037 VDD.n1091 VDD.n1090 7.147
R3038 VDD.n1088 VDD.n1087 7.147
R3039 VDD.n1085 VDD.n1084 7.147
R3040 VDD.n1080 VDD.n1079 7.147
R3041 VDD.n1077 VDD.n1076 7.147
R3042 VDD.n1074 VDD.n1073 7.147
R3043 VDD.n1070 VDD.n1069 7.147
R3044 VDD.n1067 VDD.n1066 7.147
R3045 VDD.n1064 VDD.n1063 7.147
R3046 VDD.n1061 VDD.n1060 7.147
R3047 VDD.n1058 VDD.n1057 7.147
R3048 VDD.n1053 VDD.n1052 7.147
R3049 VDD.n1050 VDD.n1049 7.147
R3050 VDD.n1046 VDD.n1045 7.147
R3051 VDD.n1043 VDD.n1042 7.147
R3052 VDD.n1040 VDD.n1039 7.147
R3053 VDD.n1037 VDD.n1036 7.147
R3054 VDD.n1032 VDD.n1031 7.147
R3055 VDD.n1112 VDD.n1111 7.147
R3056 VDD.n1646 VDD.n1645 7.147
R3057 VDD.n1648 VDD.n1647 7.147
R3058 VDD.n1650 VDD.n1649 7.147
R3059 VDD.n1630 VDD.n15 7.147
R3060 VDD.n14 VDD.n13 7.147
R3061 VDD.n12 VDD.n11 7.147
R3062 VDD.n9 VDD.n8 7.147
R3063 VDD.n7 VDD.n6 7.147
R3064 VDD.n5 VDD.n4 7.147
R3065 VDD.n2 VDD.n1 7.147
R3066 VDD.n1153 VDD.n1152 7.147
R3067 VDD.n1150 VDD.n1149 7.147
R3068 VDD.n1147 VDD.n1146 7.147
R3069 VDD.n1144 VDD.n1143 7.147
R3070 VDD.n1141 VDD.n1140 7.147
R3071 VDD.n1136 VDD.n1135 7.147
R3072 VDD.n1133 VDD.n1132 7.147
R3073 VDD.n1129 VDD.n1128 7.147
R3074 VDD.n1126 VDD.n1125 7.147
R3075 VDD.n1123 VDD.n1122 7.147
R3076 VDD.n1120 VDD.n1119 7.147
R3077 VDD.n1115 VDD.n1114 7.147
R3078 VDD.n1607 VDD.n1605 7.089
R3079 VDD.n1524 VDD.n1522 7.089
R3080 VDD.n1441 VDD.n1439 7.089
R3081 VDD.n1358 VDD.n1356 7.089
R3082 VDD.n1275 VDD.n1273 7.089
R3083 VDD.n1192 VDD.n1190 7.089
R3084 VDD.n62 VDD.n60 7.089
R3085 VDD.n145 VDD.n143 7.089
R3086 VDD.n228 VDD.n226 7.089
R3087 VDD.n311 VDD.n309 7.089
R3088 VDD.n394 VDD.n392 7.089
R3089 VDD.n477 VDD.n475 7.089
R3090 VDD.n560 VDD.n558 7.089
R3091 VDD.n643 VDD.n641 7.089
R3092 VDD.n726 VDD.n724 7.089
R3093 VDD.n809 VDD.n807 7.089
R3094 VDD.n892 VDD.n890 7.089
R3095 VDD.n975 VDD.n973 7.089
R3096 VDD.n1058 VDD.n1056 7.089
R3097 VDD.n1141 VDD.n1139 7.089
R3098 VDD.n1640 VDD.n1639 6.64
R3099 VDD.n1646 VDD.n1644 5.321
R3100 VDD.n1614 VDD.n1612 4.945
R3101 VDD.n1531 VDD.n1529 4.945
R3102 VDD.n1448 VDD.n1446 4.945
R3103 VDD.n1365 VDD.n1363 4.945
R3104 VDD.n1282 VDD.n1280 4.945
R3105 VDD.n1199 VDD.n1197 4.945
R3106 VDD.n54 VDD.n52 4.945
R3107 VDD.n137 VDD.n135 4.945
R3108 VDD.n220 VDD.n218 4.945
R3109 VDD.n303 VDD.n301 4.945
R3110 VDD.n386 VDD.n384 4.945
R3111 VDD.n469 VDD.n467 4.945
R3112 VDD.n552 VDD.n550 4.945
R3113 VDD.n635 VDD.n633 4.945
R3114 VDD.n718 VDD.n716 4.945
R3115 VDD.n801 VDD.n799 4.945
R3116 VDD.n884 VDD.n882 4.945
R3117 VDD.n967 VDD.n965 4.945
R3118 VDD.n1050 VDD.n1048 4.945
R3119 VDD.n1133 VDD.n1131 4.945
R3120 VDD.n1644 VDD.n1642 3.497
R3121 VDD.n1555 VDD.n1551 3.497
R3122 VDD.n1472 VDD.n1468 3.497
R3123 VDD.n1389 VDD.n1385 3.497
R3124 VDD.n1306 VDD.n1302 3.497
R3125 VDD.n1223 VDD.n1219 3.497
R3126 VDD.n33 VDD.n29 3.497
R3127 VDD.n116 VDD.n112 3.497
R3128 VDD.n199 VDD.n195 3.497
R3129 VDD.n282 VDD.n278 3.497
R3130 VDD.n365 VDD.n361 3.497
R3131 VDD.n448 VDD.n444 3.497
R3132 VDD.n531 VDD.n527 3.497
R3133 VDD.n614 VDD.n610 3.497
R3134 VDD.n697 VDD.n693 3.497
R3135 VDD.n780 VDD.n776 3.497
R3136 VDD.n863 VDD.n859 3.497
R3137 VDD.n946 VDD.n942 3.497
R3138 VDD.n1029 VDD.n1025 3.497
R3139 VDD.n1112 VDD.n1108 3.497
R3140 VDD.n1590 VDD.n1588 3.132
R3141 VDD.n1507 VDD.n1505 3.132
R3142 VDD.n1424 VDD.n1422 3.132
R3143 VDD.n1341 VDD.n1339 3.132
R3144 VDD.n1258 VDD.n1256 3.132
R3145 VDD.n1175 VDD.n1173 3.132
R3146 VDD.n78 VDD.n76 3.132
R3147 VDD.n161 VDD.n159 3.132
R3148 VDD.n244 VDD.n242 3.132
R3149 VDD.n327 VDD.n325 3.132
R3150 VDD.n410 VDD.n408 3.132
R3151 VDD.n493 VDD.n491 3.132
R3152 VDD.n576 VDD.n574 3.132
R3153 VDD.n659 VDD.n657 3.132
R3154 VDD.n742 VDD.n740 3.132
R3155 VDD.n825 VDD.n823 3.132
R3156 VDD.n908 VDD.n906 3.132
R3157 VDD.n991 VDD.n989 3.132
R3158 VDD.n1074 VDD.n1072 3.132
R3159 VDD.n3 VDD.n2 3.132
R3160 VDD.n1642 VDD.n1640 2.846
R3161 VDD.n1555 VDD.n1553 2.846
R3162 VDD.n1472 VDD.n1470 2.846
R3163 VDD.n1389 VDD.n1387 2.846
R3164 VDD.n1306 VDD.n1304 2.846
R3165 VDD.n1223 VDD.n1221 2.846
R3166 VDD.n33 VDD.n31 2.846
R3167 VDD.n116 VDD.n114 2.846
R3168 VDD.n199 VDD.n197 2.846
R3169 VDD.n282 VDD.n280 2.846
R3170 VDD.n365 VDD.n363 2.846
R3171 VDD.n448 VDD.n446 2.846
R3172 VDD.n531 VDD.n529 2.846
R3173 VDD.n614 VDD.n612 2.846
R3174 VDD.n697 VDD.n695 2.846
R3175 VDD.n780 VDD.n778 2.846
R3176 VDD.n863 VDD.n861 2.846
R3177 VDD.n946 VDD.n944 2.846
R3178 VDD.n1029 VDD.n1027 2.846
R3179 VDD.n1112 VDD.n1110 2.846
R3180 VDD.n1637 VDD.n1635 2.143
R3181 VDD.n1545 VDD.n1543 2.143
R3182 VDD.n1462 VDD.n1460 2.143
R3183 VDD.n1379 VDD.n1377 2.143
R3184 VDD.n1296 VDD.n1294 2.143
R3185 VDD.n1213 VDD.n1211 2.143
R3186 VDD.n41 VDD.n39 2.143
R3187 VDD.n124 VDD.n122 2.143
R3188 VDD.n207 VDD.n205 2.143
R3189 VDD.n290 VDD.n288 2.143
R3190 VDD.n373 VDD.n371 2.143
R3191 VDD.n456 VDD.n454 2.143
R3192 VDD.n539 VDD.n537 2.143
R3193 VDD.n622 VDD.n620 2.143
R3194 VDD.n705 VDD.n703 2.143
R3195 VDD.n788 VDD.n786 2.143
R3196 VDD.n871 VDD.n869 2.143
R3197 VDD.n954 VDD.n952 2.143
R3198 VDD.n1037 VDD.n1035 2.143
R3199 VDD.n1120 VDD.n1118 2.143
R3200 VDD.n20 VDD.n19 1.618
R3201 VDD.n1653 VDD.n1652 1.539
R3202 VDD.n1569 VDD.n1567 1.483
R3203 VDD.n1486 VDD.n1484 1.483
R3204 VDD.n1403 VDD.n1401 1.483
R3205 VDD.n1320 VDD.n1318 1.483
R3206 VDD.n1237 VDD.n1235 1.483
R3207 VDD.n100 VDD.n98 1.483
R3208 VDD.n183 VDD.n181 1.483
R3209 VDD.n266 VDD.n264 1.483
R3210 VDD.n349 VDD.n347 1.483
R3211 VDD.n432 VDD.n430 1.483
R3212 VDD.n515 VDD.n513 1.483
R3213 VDD.n598 VDD.n596 1.483
R3214 VDD.n681 VDD.n679 1.483
R3215 VDD.n764 VDD.n762 1.483
R3216 VDD.n847 VDD.n845 1.483
R3217 VDD.n930 VDD.n928 1.483
R3218 VDD.n1013 VDD.n1011 1.483
R3219 VDD.n1096 VDD.n1094 1.483
R3220 VDD.n1651 VDD.n1630 1.483
R3221 VDD.n1654 VDD.n1653 1.428
R3222 VDD.n1580 VDD.n1578 0.329
R3223 VDD.n1497 VDD.n1495 0.329
R3224 VDD.n1414 VDD.n1412 0.329
R3225 VDD.n1331 VDD.n1329 0.329
R3226 VDD.n1248 VDD.n1246 0.329
R3227 VDD.n1165 VDD.n1163 0.329
R3228 VDD.n89 VDD.n87 0.329
R3229 VDD.n172 VDD.n170 0.329
R3230 VDD.n255 VDD.n253 0.329
R3231 VDD.n338 VDD.n336 0.329
R3232 VDD.n421 VDD.n419 0.329
R3233 VDD.n504 VDD.n502 0.329
R3234 VDD.n587 VDD.n585 0.329
R3235 VDD.n670 VDD.n668 0.329
R3236 VDD.n753 VDD.n751 0.329
R3237 VDD.n836 VDD.n834 0.329
R3238 VDD.n919 VDD.n917 0.329
R3239 VDD.n1002 VDD.n1000 0.329
R3240 VDD.n1085 VDD.n1083 0.329
R3241 VDD.n10 VDD.n9 0.329
R3242 VDD.n24 VDD.n21 0.119
R3243 VDD.n27 VDD.n24 0.119
R3244 VDD.n34 VDD.n27 0.119
R3245 VDD.n37 VDD.n34 0.119
R3246 VDD.n42 VDD.n37 0.119
R3247 VDD.n45 VDD.n42 0.119
R3248 VDD.n48 VDD.n45 0.119
R3249 VDD.n51 VDD.n48 0.119
R3250 VDD.n55 VDD.n51 0.119
R3251 VDD.n58 VDD.n55 0.119
R3252 VDD.n63 VDD.n58 0.119
R3253 VDD.n66 VDD.n63 0.119
R3254 VDD.n69 VDD.n66 0.119
R3255 VDD.n72 VDD.n69 0.119
R3256 VDD.n75 VDD.n72 0.119
R3257 VDD.n79 VDD.n75 0.119
R3258 VDD.n82 VDD.n79 0.119
R3259 VDD.n85 VDD.n82 0.119
R3260 VDD.n90 VDD.n85 0.119
R3261 VDD.n93 VDD.n90 0.119
R3262 VDD.n96 VDD.n93 0.119
R3263 VDD.n101 VDD.n96 0.119
R3264 VDD.n104 VDD.n101 0.119
R3265 VDD.n107 VDD.n104 0.119
R3266 VDD.n110 VDD.n107 0.119
R3267 VDD.n117 VDD.n110 0.119
R3268 VDD.n120 VDD.n117 0.119
R3269 VDD.n125 VDD.n120 0.119
R3270 VDD.n128 VDD.n125 0.119
R3271 VDD.n131 VDD.n128 0.119
R3272 VDD.n134 VDD.n131 0.119
R3273 VDD.n138 VDD.n134 0.119
R3274 VDD.n141 VDD.n138 0.119
R3275 VDD.n146 VDD.n141 0.119
R3276 VDD.n149 VDD.n146 0.119
R3277 VDD.n152 VDD.n149 0.119
R3278 VDD.n155 VDD.n152 0.119
R3279 VDD.n158 VDD.n155 0.119
R3280 VDD.n162 VDD.n158 0.119
R3281 VDD.n165 VDD.n162 0.119
R3282 VDD.n168 VDD.n165 0.119
R3283 VDD.n173 VDD.n168 0.119
R3284 VDD.n176 VDD.n173 0.119
R3285 VDD.n179 VDD.n176 0.119
R3286 VDD.n184 VDD.n179 0.119
R3287 VDD.n187 VDD.n184 0.119
R3288 VDD.n190 VDD.n187 0.119
R3289 VDD.n193 VDD.n190 0.119
R3290 VDD.n200 VDD.n193 0.119
R3291 VDD.n203 VDD.n200 0.119
R3292 VDD.n208 VDD.n203 0.119
R3293 VDD.n211 VDD.n208 0.119
R3294 VDD.n214 VDD.n211 0.119
R3295 VDD.n217 VDD.n214 0.119
R3296 VDD.n221 VDD.n217 0.119
R3297 VDD.n224 VDD.n221 0.119
R3298 VDD.n229 VDD.n224 0.119
R3299 VDD.n232 VDD.n229 0.119
R3300 VDD.n235 VDD.n232 0.119
R3301 VDD.n238 VDD.n235 0.119
R3302 VDD.n241 VDD.n238 0.119
R3303 VDD.n245 VDD.n241 0.119
R3304 VDD.n248 VDD.n245 0.119
R3305 VDD.n251 VDD.n248 0.119
R3306 VDD.n256 VDD.n251 0.119
R3307 VDD.n259 VDD.n256 0.119
R3308 VDD.n262 VDD.n259 0.119
R3309 VDD.n267 VDD.n262 0.119
R3310 VDD.n270 VDD.n267 0.119
R3311 VDD.n273 VDD.n270 0.119
R3312 VDD.n276 VDD.n273 0.119
R3313 VDD.n283 VDD.n276 0.119
R3314 VDD.n286 VDD.n283 0.119
R3315 VDD.n291 VDD.n286 0.119
R3316 VDD.n294 VDD.n291 0.119
R3317 VDD.n297 VDD.n294 0.119
R3318 VDD.n300 VDD.n297 0.119
R3319 VDD.n304 VDD.n300 0.119
R3320 VDD.n307 VDD.n304 0.119
R3321 VDD.n312 VDD.n307 0.119
R3322 VDD.n315 VDD.n312 0.119
R3323 VDD.n318 VDD.n315 0.119
R3324 VDD.n321 VDD.n318 0.119
R3325 VDD.n324 VDD.n321 0.119
R3326 VDD.n328 VDD.n324 0.119
R3327 VDD.n331 VDD.n328 0.119
R3328 VDD.n334 VDD.n331 0.119
R3329 VDD.n339 VDD.n334 0.119
R3330 VDD.n342 VDD.n339 0.119
R3331 VDD.n345 VDD.n342 0.119
R3332 VDD.n350 VDD.n345 0.119
R3333 VDD.n353 VDD.n350 0.119
R3334 VDD.n356 VDD.n353 0.119
R3335 VDD.n359 VDD.n356 0.119
R3336 VDD.n366 VDD.n359 0.119
R3337 VDD.n369 VDD.n366 0.119
R3338 VDD.n374 VDD.n369 0.119
R3339 VDD.n377 VDD.n374 0.119
R3340 VDD.n380 VDD.n377 0.119
R3341 VDD.n383 VDD.n380 0.119
R3342 VDD.n387 VDD.n383 0.119
R3343 VDD.n390 VDD.n387 0.119
R3344 VDD.n395 VDD.n390 0.119
R3345 VDD.n398 VDD.n395 0.119
R3346 VDD.n401 VDD.n398 0.119
R3347 VDD.n404 VDD.n401 0.119
R3348 VDD.n407 VDD.n404 0.119
R3349 VDD.n411 VDD.n407 0.119
R3350 VDD.n414 VDD.n411 0.119
R3351 VDD.n417 VDD.n414 0.119
R3352 VDD.n422 VDD.n417 0.119
R3353 VDD.n425 VDD.n422 0.119
R3354 VDD.n428 VDD.n425 0.119
R3355 VDD.n433 VDD.n428 0.119
R3356 VDD.n436 VDD.n433 0.119
R3357 VDD.n439 VDD.n436 0.119
R3358 VDD.n442 VDD.n439 0.119
R3359 VDD.n449 VDD.n442 0.119
R3360 VDD.n452 VDD.n449 0.119
R3361 VDD.n457 VDD.n452 0.119
R3362 VDD.n460 VDD.n457 0.119
R3363 VDD.n463 VDD.n460 0.119
R3364 VDD.n466 VDD.n463 0.119
R3365 VDD.n470 VDD.n466 0.119
R3366 VDD.n473 VDD.n470 0.119
R3367 VDD.n478 VDD.n473 0.119
R3368 VDD.n481 VDD.n478 0.119
R3369 VDD.n484 VDD.n481 0.119
R3370 VDD.n487 VDD.n484 0.119
R3371 VDD.n490 VDD.n487 0.119
R3372 VDD.n494 VDD.n490 0.119
R3373 VDD.n497 VDD.n494 0.119
R3374 VDD.n500 VDD.n497 0.119
R3375 VDD.n505 VDD.n500 0.119
R3376 VDD.n508 VDD.n505 0.119
R3377 VDD.n511 VDD.n508 0.119
R3378 VDD.n516 VDD.n511 0.119
R3379 VDD.n519 VDD.n516 0.119
R3380 VDD.n522 VDD.n519 0.119
R3381 VDD.n525 VDD.n522 0.119
R3382 VDD.n532 VDD.n525 0.119
R3383 VDD.n535 VDD.n532 0.119
R3384 VDD.n540 VDD.n535 0.119
R3385 VDD.n543 VDD.n540 0.119
R3386 VDD.n546 VDD.n543 0.119
R3387 VDD.n549 VDD.n546 0.119
R3388 VDD.n553 VDD.n549 0.119
R3389 VDD.n556 VDD.n553 0.119
R3390 VDD.n561 VDD.n556 0.119
R3391 VDD.n564 VDD.n561 0.119
R3392 VDD.n567 VDD.n564 0.119
R3393 VDD.n570 VDD.n567 0.119
R3394 VDD.n573 VDD.n570 0.119
R3395 VDD.n577 VDD.n573 0.119
R3396 VDD.n580 VDD.n577 0.119
R3397 VDD.n583 VDD.n580 0.119
R3398 VDD.n588 VDD.n583 0.119
R3399 VDD.n591 VDD.n588 0.119
R3400 VDD.n594 VDD.n591 0.119
R3401 VDD.n599 VDD.n594 0.119
R3402 VDD.n602 VDD.n599 0.119
R3403 VDD.n605 VDD.n602 0.119
R3404 VDD.n608 VDD.n605 0.119
R3405 VDD.n615 VDD.n608 0.119
R3406 VDD.n618 VDD.n615 0.119
R3407 VDD.n623 VDD.n618 0.119
R3408 VDD.n626 VDD.n623 0.119
R3409 VDD.n629 VDD.n626 0.119
R3410 VDD.n632 VDD.n629 0.119
R3411 VDD.n636 VDD.n632 0.119
R3412 VDD.n639 VDD.n636 0.119
R3413 VDD.n644 VDD.n639 0.119
R3414 VDD.n647 VDD.n644 0.119
R3415 VDD.n650 VDD.n647 0.119
R3416 VDD.n653 VDD.n650 0.119
R3417 VDD.n656 VDD.n653 0.119
R3418 VDD.n660 VDD.n656 0.119
R3419 VDD.n663 VDD.n660 0.119
R3420 VDD.n666 VDD.n663 0.119
R3421 VDD.n671 VDD.n666 0.119
R3422 VDD.n674 VDD.n671 0.119
R3423 VDD.n677 VDD.n674 0.119
R3424 VDD.n682 VDD.n677 0.119
R3425 VDD.n685 VDD.n682 0.119
R3426 VDD.n688 VDD.n685 0.119
R3427 VDD.n691 VDD.n688 0.119
R3428 VDD.n698 VDD.n691 0.119
R3429 VDD.n701 VDD.n698 0.119
R3430 VDD.n706 VDD.n701 0.119
R3431 VDD.n709 VDD.n706 0.119
R3432 VDD.n712 VDD.n709 0.119
R3433 VDD.n715 VDD.n712 0.119
R3434 VDD.n719 VDD.n715 0.119
R3435 VDD.n722 VDD.n719 0.119
R3436 VDD.n727 VDD.n722 0.119
R3437 VDD.n730 VDD.n727 0.119
R3438 VDD.n733 VDD.n730 0.119
R3439 VDD.n736 VDD.n733 0.119
R3440 VDD.n739 VDD.n736 0.119
R3441 VDD.n743 VDD.n739 0.119
R3442 VDD.n746 VDD.n743 0.119
R3443 VDD.n749 VDD.n746 0.119
R3444 VDD.n754 VDD.n749 0.119
R3445 VDD.n757 VDD.n754 0.119
R3446 VDD.n760 VDD.n757 0.119
R3447 VDD.n765 VDD.n760 0.119
R3448 VDD.n768 VDD.n765 0.119
R3449 VDD.n771 VDD.n768 0.119
R3450 VDD.n774 VDD.n771 0.119
R3451 VDD.n781 VDD.n774 0.119
R3452 VDD.n784 VDD.n781 0.119
R3453 VDD.n789 VDD.n784 0.119
R3454 VDD.n792 VDD.n789 0.119
R3455 VDD.n795 VDD.n792 0.119
R3456 VDD.n798 VDD.n795 0.119
R3457 VDD.n802 VDD.n798 0.119
R3458 VDD.n805 VDD.n802 0.119
R3459 VDD.n810 VDD.n805 0.119
R3460 VDD.n813 VDD.n810 0.119
R3461 VDD.n816 VDD.n813 0.119
R3462 VDD.n819 VDD.n816 0.119
R3463 VDD.n822 VDD.n819 0.119
R3464 VDD.n826 VDD.n822 0.119
R3465 VDD.n829 VDD.n826 0.119
R3466 VDD.n832 VDD.n829 0.119
R3467 VDD.n837 VDD.n832 0.119
R3468 VDD.n840 VDD.n837 0.119
R3469 VDD.n843 VDD.n840 0.119
R3470 VDD.n848 VDD.n843 0.119
R3471 VDD.n851 VDD.n848 0.119
R3472 VDD.n854 VDD.n851 0.119
R3473 VDD.n857 VDD.n854 0.119
R3474 VDD.n864 VDD.n857 0.119
R3475 VDD.n867 VDD.n864 0.119
R3476 VDD.n872 VDD.n867 0.119
R3477 VDD.n875 VDD.n872 0.119
R3478 VDD.n878 VDD.n875 0.119
R3479 VDD.n881 VDD.n878 0.119
R3480 VDD.n885 VDD.n881 0.119
R3481 VDD.n888 VDD.n885 0.119
R3482 VDD.n893 VDD.n888 0.119
R3483 VDD.n896 VDD.n893 0.119
R3484 VDD.n899 VDD.n896 0.119
R3485 VDD.n902 VDD.n899 0.119
R3486 VDD.n905 VDD.n902 0.119
R3487 VDD.n909 VDD.n905 0.119
R3488 VDD.n912 VDD.n909 0.119
R3489 VDD.n915 VDD.n912 0.119
R3490 VDD.n920 VDD.n915 0.119
R3491 VDD.n923 VDD.n920 0.119
R3492 VDD.n926 VDD.n923 0.119
R3493 VDD.n931 VDD.n926 0.119
R3494 VDD.n934 VDD.n931 0.119
R3495 VDD.n937 VDD.n934 0.119
R3496 VDD.n940 VDD.n937 0.119
R3497 VDD.n947 VDD.n940 0.119
R3498 VDD.n950 VDD.n947 0.119
R3499 VDD.n955 VDD.n950 0.119
R3500 VDD.n958 VDD.n955 0.119
R3501 VDD.n961 VDD.n958 0.119
R3502 VDD.n964 VDD.n961 0.119
R3503 VDD.n968 VDD.n964 0.119
R3504 VDD.n971 VDD.n968 0.119
R3505 VDD.n976 VDD.n971 0.119
R3506 VDD.n979 VDD.n976 0.119
R3507 VDD.n982 VDD.n979 0.119
R3508 VDD.n985 VDD.n982 0.119
R3509 VDD.n988 VDD.n985 0.119
R3510 VDD.n992 VDD.n988 0.119
R3511 VDD.n995 VDD.n992 0.119
R3512 VDD.n998 VDD.n995 0.119
R3513 VDD.n1003 VDD.n998 0.119
R3514 VDD.n1006 VDD.n1003 0.119
R3515 VDD.n1009 VDD.n1006 0.119
R3516 VDD.n1014 VDD.n1009 0.119
R3517 VDD.n1017 VDD.n1014 0.119
R3518 VDD.n1020 VDD.n1017 0.119
R3519 VDD.n1023 VDD.n1020 0.119
R3520 VDD.n1030 VDD.n1023 0.119
R3521 VDD.n1033 VDD.n1030 0.119
R3522 VDD.n1038 VDD.n1033 0.119
R3523 VDD.n1041 VDD.n1038 0.119
R3524 VDD.n1044 VDD.n1041 0.119
R3525 VDD.n1047 VDD.n1044 0.119
R3526 VDD.n1051 VDD.n1047 0.119
R3527 VDD.n1054 VDD.n1051 0.119
R3528 VDD.n1059 VDD.n1054 0.119
R3529 VDD.n1062 VDD.n1059 0.119
R3530 VDD.n1065 VDD.n1062 0.119
R3531 VDD.n1068 VDD.n1065 0.119
R3532 VDD.n1071 VDD.n1068 0.119
R3533 VDD.n1075 VDD.n1071 0.119
R3534 VDD.n1078 VDD.n1075 0.119
R3535 VDD.n1081 VDD.n1078 0.119
R3536 VDD.n1086 VDD.n1081 0.119
R3537 VDD.n1089 VDD.n1086 0.119
R3538 VDD.n1092 VDD.n1089 0.119
R3539 VDD.n1097 VDD.n1092 0.119
R3540 VDD.n1100 VDD.n1097 0.119
R3541 VDD.n1103 VDD.n1100 0.119
R3542 VDD.n1106 VDD.n1103 0.119
R3543 VDD.n1113 VDD.n1106 0.119
R3544 VDD.n1116 VDD.n1113 0.119
R3545 VDD.n1121 VDD.n1116 0.119
R3546 VDD.n1124 VDD.n1121 0.119
R3547 VDD.n1127 VDD.n1124 0.119
R3548 VDD.n1130 VDD.n1127 0.119
R3549 VDD.n1134 VDD.n1130 0.119
R3550 VDD.n1137 VDD.n1134 0.119
R3551 VDD.n1142 VDD.n1137 0.119
R3552 VDD.n1145 VDD.n1142 0.119
R3553 VDD.n1148 VDD.n1145 0.119
R3554 VDD.n1151 VDD.n1148 0.119
R3555 VDD.n1154 VDD.n1151 0.119
R3556 VDD.n1155 VDD.n1154 0.119
R3557 VDD.n1156 VDD.n1155 0.119
R3558 VDD.n1157 VDD.n1156 0.119
R3559 VDD.n1158 VDD.n1157 0.119
R3560 VDD.n1159 VDD.n1158 0.119
R3561 VDD.n1160 VDD.n1159 0.119
R3562 VDD.n1629 VDD.n1160 0.119
R3563 VDD.n1629 VDD.n1628 0.119
R3564 VDD.n1628 VDD.n1627 0.119
R3565 VDD.n1627 VDD.n1626 0.119
R3566 VDD.n1626 VDD.n1625 0.119
R3567 VDD.n1625 VDD.n1624 0.119
R3568 VDD.n1624 VDD.n1623 0.119
R3569 VDD.n1623 VDD.n1622 0.119
R3570 VDD.n1622 VDD.n1621 0.119
R3571 VDD.n1621 VDD.n1618 0.119
R3572 VDD.n1618 VDD.n1615 0.119
R3573 VDD.n1615 VDD.n1611 0.119
R3574 VDD.n1611 VDD.n1608 0.119
R3575 VDD.n1608 VDD.n1603 0.119
R3576 VDD.n1603 VDD.n1600 0.119
R3577 VDD.n1600 VDD.n1597 0.119
R3578 VDD.n1597 VDD.n1594 0.119
R3579 VDD.n1594 VDD.n1591 0.119
R3580 VDD.n1591 VDD.n1587 0.119
R3581 VDD.n1587 VDD.n1584 0.119
R3582 VDD.n1584 VDD.n1581 0.119
R3583 VDD.n1581 VDD.n1576 0.119
R3584 VDD.n1576 VDD.n1573 0.119
R3585 VDD.n1573 VDD.n1570 0.119
R3586 VDD.n1570 VDD.n1565 0.119
R3587 VDD.n1565 VDD.n1562 0.119
R3588 VDD.n1562 VDD.n1559 0.119
R3589 VDD.n1559 VDD.n1556 0.119
R3590 VDD.n1556 VDD.n1549 0.119
R3591 VDD.n1549 VDD.n1546 0.119
R3592 VDD.n1546 VDD.n1541 0.119
R3593 VDD.n1541 VDD.n1538 0.119
R3594 VDD.n1538 VDD.n1535 0.119
R3595 VDD.n1535 VDD.n1532 0.119
R3596 VDD.n1532 VDD.n1528 0.119
R3597 VDD.n1528 VDD.n1525 0.119
R3598 VDD.n1525 VDD.n1520 0.119
R3599 VDD.n1520 VDD.n1517 0.119
R3600 VDD.n1517 VDD.n1514 0.119
R3601 VDD.n1514 VDD.n1511 0.119
R3602 VDD.n1511 VDD.n1508 0.119
R3603 VDD.n1508 VDD.n1504 0.119
R3604 VDD.n1504 VDD.n1501 0.119
R3605 VDD.n1501 VDD.n1498 0.119
R3606 VDD.n1498 VDD.n1493 0.119
R3607 VDD.n1493 VDD.n1490 0.119
R3608 VDD.n1490 VDD.n1487 0.119
R3609 VDD.n1487 VDD.n1482 0.119
R3610 VDD.n1482 VDD.n1479 0.119
R3611 VDD.n1479 VDD.n1476 0.119
R3612 VDD.n1476 VDD.n1473 0.119
R3613 VDD.n1473 VDD.n1466 0.119
R3614 VDD.n1466 VDD.n1463 0.119
R3615 VDD.n1463 VDD.n1458 0.119
R3616 VDD.n1458 VDD.n1455 0.119
R3617 VDD.n1455 VDD.n1452 0.119
R3618 VDD.n1452 VDD.n1449 0.119
R3619 VDD.n1449 VDD.n1445 0.119
R3620 VDD.n1445 VDD.n1442 0.119
R3621 VDD.n1442 VDD.n1437 0.119
R3622 VDD.n1437 VDD.n1434 0.119
R3623 VDD.n1434 VDD.n1431 0.119
R3624 VDD.n1431 VDD.n1428 0.119
R3625 VDD.n1428 VDD.n1425 0.119
R3626 VDD.n1425 VDD.n1421 0.119
R3627 VDD.n1421 VDD.n1418 0.119
R3628 VDD.n1418 VDD.n1415 0.119
R3629 VDD.n1415 VDD.n1410 0.119
R3630 VDD.n1410 VDD.n1407 0.119
R3631 VDD.n1407 VDD.n1404 0.119
R3632 VDD.n1404 VDD.n1399 0.119
R3633 VDD.n1399 VDD.n1396 0.119
R3634 VDD.n1396 VDD.n1393 0.119
R3635 VDD.n1393 VDD.n1390 0.119
R3636 VDD.n1390 VDD.n1383 0.119
R3637 VDD.n1383 VDD.n1380 0.119
R3638 VDD.n1380 VDD.n1375 0.119
R3639 VDD.n1375 VDD.n1372 0.119
R3640 VDD.n1372 VDD.n1369 0.119
R3641 VDD.n1369 VDD.n1366 0.119
R3642 VDD.n1366 VDD.n1362 0.119
R3643 VDD.n1362 VDD.n1359 0.119
R3644 VDD.n1359 VDD.n1354 0.119
R3645 VDD.n1354 VDD.n1351 0.119
R3646 VDD.n1351 VDD.n1348 0.119
R3647 VDD.n1348 VDD.n1345 0.119
R3648 VDD.n1345 VDD.n1342 0.119
R3649 VDD.n1342 VDD.n1338 0.119
R3650 VDD.n1338 VDD.n1335 0.119
R3651 VDD.n1335 VDD.n1332 0.119
R3652 VDD.n1332 VDD.n1327 0.119
R3653 VDD.n1327 VDD.n1324 0.119
R3654 VDD.n1324 VDD.n1321 0.119
R3655 VDD.n1321 VDD.n1316 0.119
R3656 VDD.n1316 VDD.n1313 0.119
R3657 VDD.n1313 VDD.n1310 0.119
R3658 VDD.n1310 VDD.n1307 0.119
R3659 VDD.n1307 VDD.n1300 0.119
R3660 VDD.n1300 VDD.n1297 0.119
R3661 VDD.n1297 VDD.n1292 0.119
R3662 VDD.n1292 VDD.n1289 0.119
R3663 VDD.n1289 VDD.n1286 0.119
R3664 VDD.n1286 VDD.n1283 0.119
R3665 VDD.n1283 VDD.n1279 0.119
R3666 VDD.n1279 VDD.n1276 0.119
R3667 VDD.n1276 VDD.n1271 0.119
R3668 VDD.n1271 VDD.n1268 0.119
R3669 VDD.n1268 VDD.n1265 0.119
R3670 VDD.n1265 VDD.n1262 0.119
R3671 VDD.n1262 VDD.n1259 0.119
R3672 VDD.n1259 VDD.n1255 0.119
R3673 VDD.n1255 VDD.n1252 0.119
R3674 VDD.n1252 VDD.n1249 0.119
R3675 VDD.n1249 VDD.n1244 0.119
R3676 VDD.n1244 VDD.n1241 0.119
R3677 VDD.n1241 VDD.n1238 0.119
R3678 VDD.n1238 VDD.n1233 0.119
R3679 VDD.n1233 VDD.n1230 0.119
R3680 VDD.n1230 VDD.n1227 0.119
R3681 VDD.n1227 VDD.n1224 0.119
R3682 VDD.n1224 VDD.n1217 0.119
R3683 VDD.n1217 VDD.n1214 0.119
R3684 VDD.n1214 VDD.n1209 0.119
R3685 VDD.n1209 VDD.n1206 0.119
R3686 VDD.n1206 VDD.n1203 0.119
R3687 VDD.n1203 VDD.n1200 0.119
R3688 VDD.n1200 VDD.n1196 0.119
R3689 VDD.n1196 VDD.n1193 0.119
R3690 VDD.n1193 VDD.n1188 0.119
R3691 VDD.n1188 VDD.n1185 0.119
R3692 VDD.n1185 VDD.n1182 0.119
R3693 VDD.n1182 VDD.n1179 0.119
R3694 VDD.n1179 VDD.n1176 0.119
R3695 VDD.n1176 VDD.n1172 0.119
R3696 VDD.n1172 VDD.n1169 0.119
R3697 VDD.n1169 VDD.n1166 0.119
R3698 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t2 203.459
R3699 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t5 187.847
R3700 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t3 164.979
R3701 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t4 149.105
R3702 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t1 143.732
R3703 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n1 76
R3704 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n3 73.482
R3705 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n2 50.925
R3706 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_193_47.n0 41.551
R3707 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t4 366.855
R3708 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t5 174.055
R3709 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n0 117.298
R3710 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n1 77.111
R3711 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t2 70
R3712 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n3 68.011
R3713 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t3 63.321
R3714 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.t0 61.666
R3715 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1108_47.n2 57.017
R3716 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1462_47.t1 87.142
R3717 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t2 530.008
R3718 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t4 334.888
R3719 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t6 255.459
R3720 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t3 224.611
R3721 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t7 196.882
R3722 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t5 141.921
R3723 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n9 126.03
R3724 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.t0 99.672
R3725 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n1 92.562
R3726 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n0 44.57
R3727 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n2 38.638
R3728 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n6 15
R3729 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n8 15
R3730 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n4 13.653
R3731 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n7 3.182
R3732 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n3 1.366
R3733 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[0]/a_27_47.n5 1.326
R3734 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t5 332.579
R3735 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t4 168.699
R3736 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n1 104.381
R3737 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n0 101.869
R3738 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t3 96.154
R3739 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n2 92.648
R3740 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n3 65.666
R3741 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t2 65
R3742 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_543_47.t1 45
R3743 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.t1 194.654
R3744 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.t2 168.384
R3745 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_651_413.n0 63.321
R3746 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t3 333.651
R3747 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t2 297.233
R3748 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t4 294.554
R3749 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t5 211.008
R3750 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t1 102.408
R3751 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t0 50.774
R3752 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D.n1 49.535
R3753 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/D 20.838
R3754 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D.n0 9.965
R3755 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D.n4 7.455
R3756 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n3 3.763
R3757 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n2 3.763
R3758 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[0]/D 2.855
R3759 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[0]/D 1.297
R3760 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n0 163.71
R3761 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n1 82.083
R3762 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.t3 63.333
R3763 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.t2 63.321
R3764 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_448_47.t1 29.726
R3765 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/Q.t0 59.048
R3766 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/Q.t1 50.115
R3767 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1270_413.t1 126.642
R3768 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[0]/a_1217_47.t0 94.726
R3769 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t4 350.253
R3770 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t5 189.586
R3771 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n1 97.205
R3772 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t3 89.119
R3773 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n0 79.305
R3774 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n2 66.705
R3775 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t1 63.333
R3776 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n3 41.041
R3777 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_761_289.t0 31.979
R3778 sky130_fd_sc_hd__dfrbp_1_0[1]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_639_47.t0 198.571
R3779 sky130_fd_sc_hd__dfrbp_1_0[1]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_805_47.t1 60
R3780 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t6 389.181
R3781 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t3 256.987
R3782 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t8 212.079
R3783 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t7 174.888
R3784 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t4 163.801
R3785 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n0 161.578
R3786 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t5 139.779
R3787 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n1 129.263
R3788 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n5 102.015
R3789 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t1 63.321
R3790 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t2 63.321
R3791 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n6 46.071
R3792 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n3 37.442
R3793 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n4 23.54
R3794 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1283_21.n2 22.639
R3795 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.t3 239.038
R3796 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.t2 166.738
R3797 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n1 95.895
R3798 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.t0 71.217
R3799 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1847_47.n0 30.051
R3800 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t2 203.459
R3801 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t5 187.847
R3802 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t3 164.979
R3803 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t4 149.105
R3804 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t1 143.732
R3805 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n1 76
R3806 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n3 73.482
R3807 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n2 50.925
R3808 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_193_47.n0 41.551
R3809 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t4 366.855
R3810 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t5 174.055
R3811 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n0 117.298
R3812 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n1 77.111
R3813 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t2 70
R3814 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t3 68.011
R3815 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n3 63.321
R3816 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.t0 61.666
R3817 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1108_47.n2 57.017
R3818 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1462_47.t1 87.142
R3819 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t2 530.008
R3820 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t4 334.888
R3821 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t6 255.459
R3822 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t3 224.611
R3823 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t7 196.882
R3824 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t5 141.921
R3825 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n9 126.03
R3826 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.t0 99.672
R3827 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n1 92.562
R3828 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n0 44.57
R3829 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n2 38.638
R3830 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n6 15
R3831 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n8 15
R3832 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n4 13.653
R3833 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n7 3.182
R3834 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n3 1.366
R3835 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[1]/a_27_47.n5 1.326
R3836 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t5 332.579
R3837 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t4 168.699
R3838 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n1 104.381
R3839 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n0 101.869
R3840 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t3 96.154
R3841 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n2 92.648
R3842 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n3 65.666
R3843 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t2 65
R3844 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_543_47.t1 45
R3845 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.n0 194.654
R3846 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.t2 168.384
R3847 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_651_413.t1 63.321
R3848 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t3 333.651
R3849 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t2 297.233
R3850 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t4 294.554
R3851 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t5 211.008
R3852 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t1 102.408
R3853 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/D.t0 50.774
R3854 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[1]/D.n1 49.535
R3855 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/D 20.838
R3856 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[1]/D.n0 9.965
R3857 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[1]/D.n4 7.455
R3858 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n3 3.763
R3859 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n2 3.763
R3860 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[1]/D 2.855
R3861 sky130_fd_sc_hd__dfrbp_1_0[1]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[1]/D 1.297
R3862 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n0 163.71
R3863 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n1 82.083
R3864 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.t1 63.333
R3865 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.t3 63.321
R3866 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_448_47.t2 29.726
R3867 sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/Q.t0 59.048
R3868 sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/Q.t1 50.115
R3869 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1270_413.t1 126.642
R3870 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[1]/a_1217_47.t1 94.726
R3871 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t4 350.253
R3872 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t5 189.586
R3873 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n1 97.205
R3874 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t0 89.119
R3875 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n0 79.305
R3876 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n2 66.705
R3877 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t2 63.333
R3878 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n3 41.041
R3879 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_761_289.t3 31.979
R3880 sky130_fd_sc_hd__dfrbp_1_0[2]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_639_47.t0 198.571
R3881 sky130_fd_sc_hd__dfrbp_1_0[2]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_805_47.t1 60
R3882 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t6 389.181
R3883 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t3 256.987
R3884 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t8 212.079
R3885 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t7 174.888
R3886 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t4 163.801
R3887 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n0 161.578
R3888 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t5 139.779
R3889 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n1 129.263
R3890 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n5 102.015
R3891 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t1 63.321
R3892 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t2 63.321
R3893 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n6 46.071
R3894 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n3 37.442
R3895 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n4 23.54
R3896 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1283_21.n2 22.639
R3897 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.t3 239.038
R3898 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.t2 166.738
R3899 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n1 95.895
R3900 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.t0 71.217
R3901 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1847_47.n0 30.051
R3902 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t2 203.459
R3903 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t5 187.847
R3904 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t3 164.979
R3905 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t4 149.105
R3906 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t0 143.732
R3907 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n1 76
R3908 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n3 73.482
R3909 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n2 50.925
R3910 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_193_47.n0 41.551
R3911 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t4 366.855
R3912 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t5 174.055
R3913 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n0 117.298
R3914 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n1 77.111
R3915 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t2 70
R3916 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t3 68.011
R3917 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n3 63.321
R3918 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.t0 61.666
R3919 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1108_47.n2 57.017
R3920 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1462_47.t1 87.142
R3921 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t2 530.008
R3922 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t4 334.888
R3923 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t6 255.459
R3924 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t3 224.611
R3925 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t7 196.882
R3926 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t5 141.921
R3927 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n9 126.03
R3928 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.t0 99.672
R3929 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n1 92.562
R3930 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n0 44.57
R3931 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n2 38.638
R3932 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n6 15
R3933 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n8 15
R3934 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n4 13.653
R3935 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n7 3.182
R3936 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n3 1.366
R3937 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[2]/a_27_47.n5 1.326
R3938 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t5 332.579
R3939 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t4 168.699
R3940 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n1 104.381
R3941 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n0 101.869
R3942 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t2 96.154
R3943 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n2 92.648
R3944 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n3 65.666
R3945 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t3 65
R3946 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_543_47.t1 45
R3947 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.n0 194.654
R3948 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.t2 168.384
R3949 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_651_413.t1 63.321
R3950 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t3 333.651
R3951 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t2 297.233
R3952 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t4 294.554
R3953 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t5 211.008
R3954 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t1 102.408
R3955 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/D.t0 50.774
R3956 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D.n1 49.535
R3957 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/D 20.838
R3958 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D.n0 9.965
R3959 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D.n4 7.455
R3960 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n3 3.763
R3961 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n2 3.763
R3962 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[2]/D 2.855
R3963 sky130_fd_sc_hd__dfrbp_1_0[2]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/D 1.297
R3964 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n0 163.71
R3965 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.t2 82.083
R3966 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.t3 63.333
R3967 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.t1 63.321
R3968 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.t0 26.393
R3969 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n2 14.4
R3970 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[2]/a_448_47.n1 3.333
R3971 sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/Q.t0 59.048
R3972 sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/Q.t1 50.115
R3973 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1270_413.t1 126.642
R3974 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[2]/a_1217_47.t1 94.726
R3975 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t4 350.253
R3976 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t5 189.586
R3977 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n1 97.205
R3978 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t0 89.119
R3979 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n0 79.305
R3980 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n2 66.705
R3981 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t2 63.333
R3982 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n3 41.041
R3983 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_761_289.t3 31.979
R3984 sky130_fd_sc_hd__dfrbp_1_0[3]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_639_47.t0 198.571
R3985 sky130_fd_sc_hd__dfrbp_1_0[3]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_805_47.t1 60
R3986 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t6 389.181
R3987 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t3 256.987
R3988 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t8 212.079
R3989 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t7 174.888
R3990 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t4 163.801
R3991 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n0 161.578
R3992 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t5 139.779
R3993 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n1 129.263
R3994 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n5 102.015
R3995 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t1 63.321
R3996 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t2 63.321
R3997 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n6 46.071
R3998 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n3 37.442
R3999 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n4 23.54
R4000 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1283_21.n2 22.639
R4001 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.t3 239.038
R4002 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.t2 166.738
R4003 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n1 95.895
R4004 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.t0 71.217
R4005 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1847_47.n0 30.051
R4006 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t2 203.459
R4007 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t5 187.847
R4008 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t3 164.979
R4009 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t4 149.105
R4010 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t1 143.732
R4011 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n1 76
R4012 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n3 73.482
R4013 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n2 50.925
R4014 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_193_47.n0 41.551
R4015 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t4 366.855
R4016 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t5 174.055
R4017 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n0 117.298
R4018 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n1 77.111
R4019 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t2 70
R4020 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n3 68.011
R4021 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t3 63.321
R4022 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.t1 61.666
R4023 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1108_47.n2 57.017
R4024 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1462_47.t1 87.142
R4025 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t2 530.008
R4026 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t4 334.888
R4027 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t6 255.459
R4028 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t3 224.611
R4029 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t7 196.882
R4030 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t5 141.921
R4031 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n9 126.03
R4032 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.t0 99.672
R4033 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n1 92.562
R4034 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n0 44.57
R4035 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n2 38.638
R4036 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n6 15
R4037 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n8 15
R4038 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n4 13.653
R4039 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n7 3.182
R4040 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n3 1.366
R4041 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[3]/a_27_47.n5 1.326
R4042 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t5 332.579
R4043 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t4 168.699
R4044 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n1 104.381
R4045 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n0 101.869
R4046 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t3 96.154
R4047 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n2 92.648
R4048 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n3 65.666
R4049 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t2 65
R4050 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_543_47.t1 45
R4051 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.n0 194.654
R4052 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.t2 168.384
R4053 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_651_413.t1 63.321
R4054 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t3 333.651
R4055 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t2 297.233
R4056 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t4 294.554
R4057 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t5 211.008
R4058 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t1 102.408
R4059 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/D.t0 50.774
R4060 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D.n1 49.535
R4061 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/D 20.838
R4062 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D.n0 9.965
R4063 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D.n4 7.455
R4064 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n3 3.763
R4065 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n2 3.763
R4066 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[3]/D 2.855
R4067 sky130_fd_sc_hd__dfrbp_1_0[3]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/D 1.297
R4068 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n0 163.71
R4069 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.t2 82.083
R4070 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.t3 63.333
R4071 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.t1 63.321
R4072 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.t0 26.393
R4073 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n2 14.4
R4074 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[3]/a_448_47.n1 3.333
R4075 sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/Q.t0 59.048
R4076 sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/Q.t1 50.115
R4077 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1270_413.t1 126.642
R4078 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[3]/a_1217_47.t1 94.726
R4079 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t4 350.253
R4080 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t5 189.586
R4081 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n1 97.205
R4082 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t1 89.119
R4083 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n0 79.305
R4084 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n2 66.705
R4085 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t2 63.333
R4086 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n3 41.041
R4087 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_761_289.t3 31.979
R4088 sky130_fd_sc_hd__dfrbp_1_0[4]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_639_47.t0 198.571
R4089 sky130_fd_sc_hd__dfrbp_1_0[4]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_805_47.t1 60
R4090 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t6 389.181
R4091 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t3 256.987
R4092 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t8 212.079
R4093 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t7 174.888
R4094 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t4 163.801
R4095 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n5 161.578
R4096 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t5 139.779
R4097 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n0 129.263
R4098 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n3 102.015
R4099 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n6 63.321
R4100 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t2 63.321
R4101 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.t1 46.071
R4102 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n2 37.442
R4103 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n4 23.54
R4104 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1283_21.n1 22.639
R4105 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.t3 239.038
R4106 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.t2 166.738
R4107 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n1 95.895
R4108 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.t0 71.217
R4109 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1847_47.n0 30.051
R4110 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t2 203.459
R4111 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t5 187.847
R4112 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t3 164.979
R4113 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t4 149.105
R4114 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t0 143.732
R4115 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n1 76
R4116 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n3 73.482
R4117 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n2 50.925
R4118 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_193_47.n0 41.551
R4119 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t4 366.855
R4120 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t5 174.055
R4121 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n0 117.298
R4122 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n1 77.111
R4123 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t3 70
R4124 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n3 68.011
R4125 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t2 63.321
R4126 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.t1 61.666
R4127 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1108_47.n2 57.017
R4128 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1462_47.t1 87.142
R4129 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t2 530.008
R4130 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t4 334.888
R4131 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t6 255.459
R4132 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t3 224.611
R4133 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t7 196.882
R4134 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t5 141.921
R4135 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n9 126.03
R4136 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.t0 99.672
R4137 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n1 92.562
R4138 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n0 44.57
R4139 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n2 38.638
R4140 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n6 15
R4141 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n8 15
R4142 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n4 13.653
R4143 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n7 3.182
R4144 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n3 1.366
R4145 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[4]/a_27_47.n5 1.326
R4146 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t5 332.579
R4147 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t4 168.699
R4148 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n1 104.381
R4149 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n0 101.869
R4150 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n3 96.154
R4151 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n2 92.648
R4152 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t2 65.666
R4153 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t1 65
R4154 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_543_47.t3 45
R4155 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.n0 194.654
R4156 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.t2 168.384
R4157 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_651_413.t1 63.321
R4158 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t3 333.651
R4159 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t2 297.233
R4160 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t4 294.554
R4161 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t5 211.008
R4162 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t1 102.408
R4163 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t0 50.774
R4164 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D.n1 49.535
R4165 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/D 20.838
R4166 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D.n0 9.965
R4167 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D.n4 7.455
R4168 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n3 3.763
R4169 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n2 3.763
R4170 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[4]/D 2.855
R4171 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[4]/D 1.297
R4172 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n0 163.71
R4173 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n1 82.083
R4174 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.t0 63.333
R4175 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.t3 63.321
R4176 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_448_47.t2 29.726
R4177 sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[4]/Q.t0 59.048
R4178 sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[4]/Q.t1 50.115
R4179 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1270_413.t1 126.642
R4180 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[4]/a_1217_47.t0 94.726
R4181 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t4 350.253
R4182 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t5 189.586
R4183 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n1 97.205
R4184 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t0 89.119
R4185 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n0 79.305
R4186 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n2 66.705
R4187 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t2 63.333
R4188 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n3 41.041
R4189 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_761_289.t1 31.979
R4190 sky130_fd_sc_hd__dfrbp_1_0[5]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_639_47.t0 198.571
R4191 sky130_fd_sc_hd__dfrbp_1_0[5]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_805_47.t1 60
R4192 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t6 389.181
R4193 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t3 256.987
R4194 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t8 212.079
R4195 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t7 174.888
R4196 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t4 163.801
R4197 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n5 161.578
R4198 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t5 139.779
R4199 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n0 129.263
R4200 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n3 102.015
R4201 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n6 63.321
R4202 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t2 63.321
R4203 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.t1 46.071
R4204 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n2 37.442
R4205 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n4 23.54
R4206 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1283_21.n1 22.639
R4207 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.t3 239.038
R4208 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.t2 166.738
R4209 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n1 95.895
R4210 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.t0 71.217
R4211 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1847_47.n0 30.051
R4212 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t2 203.459
R4213 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t5 187.847
R4214 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t3 164.979
R4215 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t4 149.105
R4216 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t1 143.732
R4217 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n1 76
R4218 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n3 73.482
R4219 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n2 50.925
R4220 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_193_47.n0 41.551
R4221 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t4 366.855
R4222 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t5 174.055
R4223 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n0 117.298
R4224 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n1 77.111
R4225 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t3 70
R4226 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n3 68.011
R4227 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t2 63.321
R4228 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.t1 61.666
R4229 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1108_47.n2 57.017
R4230 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1462_47.t1 87.142
R4231 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t2 530.008
R4232 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t4 334.888
R4233 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t6 255.459
R4234 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t3 224.611
R4235 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t7 196.882
R4236 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t5 141.921
R4237 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n9 126.03
R4238 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.t0 99.672
R4239 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n1 92.562
R4240 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n0 44.57
R4241 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n2 38.638
R4242 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n6 15
R4243 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n8 15
R4244 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n4 13.653
R4245 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n7 3.182
R4246 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n3 1.366
R4247 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[5]/a_27_47.n5 1.326
R4248 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t5 332.579
R4249 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t4 168.699
R4250 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n1 104.381
R4251 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n0 101.869
R4252 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n3 96.154
R4253 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n2 92.648
R4254 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t3 65.666
R4255 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t0 65
R4256 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_543_47.t2 45
R4257 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.n0 194.654
R4258 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.t2 168.384
R4259 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_651_413.t1 63.321
R4260 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t3 333.651
R4261 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t2 297.233
R4262 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t4 294.554
R4263 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t5 211.008
R4264 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t1 102.408
R4265 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/D.t0 50.774
R4266 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D.n1 49.535
R4267 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/D 20.838
R4268 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D.n0 9.965
R4269 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D.n4 7.455
R4270 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n3 3.763
R4271 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n2 3.763
R4272 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[5]/D 2.855
R4273 sky130_fd_sc_hd__dfrbp_1_0[5]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/D 1.297
R4274 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n0 163.71
R4275 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.t3 82.083
R4276 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.t0 63.333
R4277 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.t2 63.321
R4278 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.t1 26.393
R4279 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n2 14.4
R4280 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[5]/a_448_47.n1 3.333
R4281 sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/Q.t0 59.048
R4282 sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/Q.t1 50.115
R4283 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1270_413.t1 126.642
R4284 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[5]/a_1217_47.t0 94.726
R4285 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t4 350.253
R4286 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t5 189.586
R4287 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n1 97.205
R4288 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t0 89.119
R4289 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n0 79.305
R4290 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n2 66.705
R4291 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t3 63.333
R4292 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n3 41.041
R4293 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_761_289.t1 31.979
R4294 sky130_fd_sc_hd__dfrbp_1_0[6]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_639_47.t0 198.571
R4295 sky130_fd_sc_hd__dfrbp_1_0[6]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_805_47.t1 60
R4296 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t6 389.181
R4297 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t3 256.987
R4298 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t8 212.079
R4299 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t7 174.888
R4300 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t4 163.801
R4301 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n0 161.578
R4302 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t5 139.779
R4303 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n1 129.263
R4304 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n5 102.015
R4305 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t1 63.321
R4306 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t2 63.321
R4307 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n6 46.071
R4308 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n3 37.442
R4309 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n4 23.54
R4310 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1283_21.n2 22.639
R4311 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.t3 239.038
R4312 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.t2 166.738
R4313 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n1 95.895
R4314 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.t0 71.217
R4315 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1847_47.n0 30.051
R4316 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t2 203.459
R4317 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t5 187.847
R4318 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t3 164.979
R4319 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t4 149.105
R4320 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t0 143.732
R4321 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n1 76
R4322 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n3 73.482
R4323 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n2 50.925
R4324 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_193_47.n0 41.551
R4325 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t4 366.855
R4326 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t5 174.055
R4327 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n0 117.298
R4328 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n1 77.111
R4329 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t2 70
R4330 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n3 68.011
R4331 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t1 63.321
R4332 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.t3 61.666
R4333 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1108_47.n2 57.017
R4334 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1462_47.t1 87.142
R4335 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t2 530.008
R4336 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t4 334.888
R4337 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t6 255.459
R4338 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t3 224.611
R4339 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t7 196.882
R4340 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t5 141.921
R4341 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n9 126.03
R4342 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.t0 99.672
R4343 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n1 92.562
R4344 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n0 44.57
R4345 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n2 38.638
R4346 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n6 15
R4347 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n8 15
R4348 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n4 13.653
R4349 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n7 3.182
R4350 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n3 1.366
R4351 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[6]/a_27_47.n5 1.326
R4352 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t5 332.579
R4353 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t4 168.699
R4354 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n1 104.381
R4355 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n0 101.869
R4356 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t3 96.154
R4357 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n2 92.648
R4358 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n3 65.666
R4359 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t2 65
R4360 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_543_47.t1 45
R4361 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.n0 194.654
R4362 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.t1 168.384
R4363 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_651_413.t2 63.321
R4364 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t3 333.651
R4365 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t2 297.233
R4366 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t4 294.554
R4367 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t5 211.008
R4368 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t1 102.408
R4369 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/D.t0 50.774
R4370 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D.n1 49.535
R4371 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/D 20.838
R4372 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D.n0 9.965
R4373 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D.n4 7.455
R4374 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n3 3.763
R4375 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n2 3.763
R4376 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[6]/D 2.855
R4377 sky130_fd_sc_hd__dfrbp_1_0[6]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[6]/D 1.297
R4378 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n0 163.71
R4379 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n1 82.083
R4380 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.t1 63.333
R4381 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.t3 63.321
R4382 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_448_47.t2 29.726
R4383 sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/Q.t0 59.048
R4384 sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/Q.t1 50.115
R4385 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1270_413.t1 126.642
R4386 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[6]/a_1217_47.t0 94.726
R4387 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t4 350.253
R4388 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t5 189.586
R4389 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n1 97.205
R4390 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t0 89.119
R4391 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n0 79.305
R4392 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n2 66.705
R4393 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t3 63.333
R4394 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n3 41.041
R4395 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_761_289.t1 31.979
R4396 sky130_fd_sc_hd__dfrbp_1_0[7]/a_639_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_639_47.t1 198.571
R4397 sky130_fd_sc_hd__dfrbp_1_0[7]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_805_47.t1 60
R4398 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t6 389.181
R4399 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t3 256.987
R4400 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t8 212.079
R4401 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t7 174.888
R4402 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t4 163.801
R4403 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n0 161.578
R4404 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t5 139.779
R4405 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n1 129.263
R4406 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n5 102.015
R4407 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t1 63.321
R4408 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t2 63.321
R4409 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n6 46.071
R4410 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n3 37.442
R4411 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n4 23.54
R4412 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1283_21.n2 22.639
R4413 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.t3 239.038
R4414 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.t2 166.738
R4415 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n1 95.895
R4416 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.t0 71.217
R4417 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1847_47.n0 30.051
R4418 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t2 203.459
R4419 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t5 187.847
R4420 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t3 164.979
R4421 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t4 149.105
R4422 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t1 143.732
R4423 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n1 76
R4424 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n3 73.482
R4425 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n2 50.925
R4426 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_193_47.n0 41.551
R4427 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t4 366.855
R4428 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t5 174.055
R4429 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n0 117.298
R4430 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n1 77.111
R4431 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t2 70
R4432 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n3 68.011
R4433 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t1 63.321
R4434 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.t3 61.666
R4435 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1108_47.n2 57.017
R4436 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1462_47.t1 87.142
R4437 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t2 530.008
R4438 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t4 334.888
R4439 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t6 255.459
R4440 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t3 224.611
R4441 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t7 196.882
R4442 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t5 141.921
R4443 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n9 126.03
R4444 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.t0 99.672
R4445 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n1 92.562
R4446 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n0 44.57
R4447 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n2 38.638
R4448 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n6 15
R4449 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n8 15
R4450 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n4 13.653
R4451 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n7 3.182
R4452 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n3 1.366
R4453 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[7]/a_27_47.n5 1.326
R4454 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t5 332.579
R4455 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t4 168.699
R4456 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n1 104.381
R4457 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n0 101.869
R4458 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n3 96.154
R4459 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n2 92.648
R4460 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t2 65.666
R4461 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t1 65
R4462 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_543_47.t3 45
R4463 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.t1 194.654
R4464 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.t2 168.384
R4465 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_651_413.n0 63.321
R4466 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t3 333.651
R4467 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t2 297.233
R4468 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t4 294.554
R4469 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t5 211.008
R4470 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t1 102.408
R4471 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/D.t0 50.774
R4472 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D.n1 49.535
R4473 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/D 20.838
R4474 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D.n0 9.965
R4475 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D.n4 7.455
R4476 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n3 3.763
R4477 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n2 3.763
R4478 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[7]/D 2.855
R4479 sky130_fd_sc_hd__dfrbp_1_0[7]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[7]/D 1.297
R4480 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n0 163.71
R4481 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.t1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n1 82.083
R4482 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.t0 63.333
R4483 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.t3 63.321
R4484 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_448_47.t2 29.726
R4485 sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/Q.t0 59.048
R4486 sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/Q.t1 50.115
R4487 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1270_413.t1 126.642
R4488 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[7]/a_1217_47.t0 94.726
R4489 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t4 350.253
R4490 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t5 189.586
R4491 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n1 97.205
R4492 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t2 89.119
R4493 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n0 79.305
R4494 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n2 66.705
R4495 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t0 63.333
R4496 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n3 41.041
R4497 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_761_289.t1 31.979
R4498 sky130_fd_sc_hd__dfrbp_1_0[8]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_639_47.t0 198.571
R4499 sky130_fd_sc_hd__dfrbp_1_0[8]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_805_47.t1 60
R4500 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t6 389.181
R4501 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t3 256.987
R4502 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t8 212.079
R4503 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t7 174.888
R4504 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t4 163.801
R4505 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n0 161.578
R4506 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t5 139.779
R4507 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n1 129.263
R4508 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n5 102.015
R4509 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t1 63.321
R4510 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t2 63.321
R4511 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n6 46.071
R4512 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n3 37.442
R4513 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n4 23.54
R4514 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1283_21.n2 22.639
R4515 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.t3 239.038
R4516 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.t2 166.738
R4517 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n1 95.895
R4518 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.t0 71.217
R4519 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1847_47.n0 30.051
R4520 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t2 203.459
R4521 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t5 187.847
R4522 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t3 164.979
R4523 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t4 149.105
R4524 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t0 143.732
R4525 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n1 76
R4526 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n3 73.482
R4527 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n2 50.925
R4528 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_193_47.n0 41.551
R4529 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t4 366.855
R4530 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t5 174.055
R4531 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n0 117.298
R4532 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n1 77.111
R4533 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t1 70
R4534 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t3 68.011
R4535 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n3 63.321
R4536 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.t2 61.666
R4537 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1108_47.n2 57.017
R4538 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1462_47.t1 87.142
R4539 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t2 530.008
R4540 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t4 334.888
R4541 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t6 255.459
R4542 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t3 224.611
R4543 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t7 196.882
R4544 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t5 141.921
R4545 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n9 126.03
R4546 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.t0 99.672
R4547 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n1 92.562
R4548 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n0 44.57
R4549 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n2 38.638
R4550 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n6 15
R4551 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n8 15
R4552 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n4 13.653
R4553 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n7 3.182
R4554 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n3 1.366
R4555 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[8]/a_27_47.n5 1.326
R4556 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t5 332.579
R4557 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t4 168.699
R4558 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n1 104.381
R4559 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n0 101.869
R4560 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t2 96.154
R4561 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n2 92.648
R4562 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n3 65.666
R4563 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t3 65
R4564 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_543_47.t1 45
R4565 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.n0 194.654
R4566 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.t2 168.384
R4567 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_651_413.t1 63.321
R4568 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t3 333.651
R4569 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t2 297.233
R4570 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t4 294.554
R4571 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t5 211.008
R4572 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t1 102.408
R4573 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/D.t0 50.774
R4574 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D.n1 49.535
R4575 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/D 20.838
R4576 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D.n0 9.965
R4577 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D.n4 7.455
R4578 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n3 3.763
R4579 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n2 3.763
R4580 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[8]/D 2.855
R4581 sky130_fd_sc_hd__dfrbp_1_0[8]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[8]/D 1.297
R4582 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n0 163.71
R4583 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n1 82.083
R4584 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.t1 63.333
R4585 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.t3 63.321
R4586 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_448_47.t2 29.726
R4587 sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[8]/Q.t0 59.048
R4588 sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[8]/Q.t1 50.115
R4589 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1270_413.t1 126.642
R4590 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[8]/a_1217_47.t1 94.726
R4591 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t4 350.253
R4592 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t5 189.586
R4593 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n1 97.205
R4594 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t1 89.119
R4595 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n0 79.305
R4596 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n2 66.705
R4597 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t2 63.333
R4598 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n3 41.041
R4599 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_761_289.t3 31.979
R4600 sky130_fd_sc_hd__dfrbp_1_0[9]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_639_47.t0 198.571
R4601 sky130_fd_sc_hd__dfrbp_1_0[9]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_805_47.t1 60
R4602 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t6 389.181
R4603 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t3 256.987
R4604 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t8 212.079
R4605 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t7 174.888
R4606 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t4 163.801
R4607 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n5 161.578
R4608 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t5 139.779
R4609 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n0 129.263
R4610 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n3 102.015
R4611 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n6 63.321
R4612 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t2 63.321
R4613 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.t1 46.071
R4614 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n2 37.442
R4615 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n4 23.54
R4616 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1283_21.n1 22.639
R4617 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.t3 239.038
R4618 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.t2 166.738
R4619 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n1 95.895
R4620 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.t0 71.217
R4621 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1847_47.n0 30.051
R4622 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t2 203.459
R4623 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t5 187.847
R4624 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t3 164.979
R4625 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t4 149.105
R4626 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t0 143.732
R4627 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n1 76
R4628 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n3 73.482
R4629 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n2 50.925
R4630 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_193_47.n0 41.551
R4631 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t4 366.855
R4632 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t5 174.055
R4633 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n0 117.298
R4634 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n1 77.111
R4635 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t3 70
R4636 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n3 68.011
R4637 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t2 63.321
R4638 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.t1 61.666
R4639 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1108_47.n2 57.017
R4640 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1462_47.t1 87.142
R4641 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t2 530.008
R4642 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t4 334.888
R4643 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t6 255.459
R4644 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t3 224.611
R4645 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t7 196.882
R4646 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t5 141.921
R4647 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n9 126.03
R4648 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.t0 99.672
R4649 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n1 92.562
R4650 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n0 44.57
R4651 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n2 38.638
R4652 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n6 15
R4653 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n8 15
R4654 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n4 13.653
R4655 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n7 3.182
R4656 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n3 1.366
R4657 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[9]/a_27_47.n5 1.326
R4658 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t5 332.579
R4659 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t4 168.699
R4660 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n1 104.381
R4661 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n0 101.869
R4662 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t2 96.154
R4663 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n2 92.648
R4664 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n3 65.666
R4665 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t3 65
R4666 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_543_47.t1 45
R4667 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.t1 194.654
R4668 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.t2 168.384
R4669 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_651_413.n0 63.321
R4670 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t3 333.651
R4671 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t2 297.233
R4672 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t4 294.554
R4673 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t5 211.008
R4674 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t1 102.408
R4675 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/D.t0 50.774
R4676 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D.n1 49.535
R4677 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/D 20.838
R4678 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D.n0 9.965
R4679 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D.n4 7.455
R4680 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n3 3.763
R4681 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n2 3.763
R4682 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[9]/D 2.855
R4683 sky130_fd_sc_hd__dfrbp_1_0[9]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/D 1.297
R4684 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n0 163.71
R4685 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n1 82.083
R4686 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.t3 63.333
R4687 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.t2 63.321
R4688 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_448_47.t1 29.726
R4689 sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/Q.t0 59.048
R4690 sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/Q.t1 50.115
R4691 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1270_413.t1 126.642
R4692 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/a_1217_47.t1 94.726
R4693 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t4 350.253
R4694 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t5 189.586
R4695 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n1 97.205
R4696 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t1 89.119
R4697 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n0 79.305
R4698 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n2 66.705
R4699 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t0 63.333
R4700 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n3 41.041
R4701 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_761_289.t2 31.979
R4702 sky130_fd_sc_hd__dfrbp_1_0[10]/a_639_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_639_47.t1 198.571
R4703 sky130_fd_sc_hd__dfrbp_1_0[10]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_805_47.t1 60
R4704 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t6 389.181
R4705 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t3 256.987
R4706 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t8 212.079
R4707 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t7 174.888
R4708 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t4 163.801
R4709 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n5 161.578
R4710 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t5 139.779
R4711 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n0 129.263
R4712 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n3 102.015
R4713 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n6 63.321
R4714 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t2 63.321
R4715 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.t1 46.071
R4716 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n2 37.442
R4717 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n4 23.54
R4718 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1283_21.n1 22.639
R4719 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.t3 239.038
R4720 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.t2 166.738
R4721 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n1 95.895
R4722 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.t0 71.217
R4723 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1847_47.n0 30.051
R4724 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t2 203.459
R4725 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t5 187.847
R4726 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t3 164.979
R4727 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t4 149.105
R4728 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t1 143.732
R4729 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n1 76
R4730 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n3 73.482
R4731 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n2 50.925
R4732 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_193_47.n0 41.551
R4733 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t4 366.855
R4734 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t5 174.055
R4735 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n0 117.298
R4736 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n1 77.111
R4737 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t1 70
R4738 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t2 68.011
R4739 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n3 63.321
R4740 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.t3 61.666
R4741 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1108_47.n2 57.017
R4742 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1462_47.t1 87.142
R4743 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t2 530.008
R4744 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t4 334.888
R4745 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t6 255.459
R4746 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t3 224.611
R4747 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t7 196.882
R4748 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t5 141.921
R4749 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n9 126.03
R4750 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.t0 99.672
R4751 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n1 92.562
R4752 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n0 44.57
R4753 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n2 38.638
R4754 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n6 15
R4755 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n8 15
R4756 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n4 13.653
R4757 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n7 3.182
R4758 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n3 1.366
R4759 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[10]/a_27_47.n5 1.326
R4760 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t5 332.579
R4761 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t4 168.699
R4762 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n1 104.381
R4763 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n0 101.869
R4764 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t2 96.154
R4765 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n2 92.648
R4766 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n3 65.666
R4767 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t3 65
R4768 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_543_47.t1 45
R4769 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.t1 194.654
R4770 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.t2 168.384
R4771 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_651_413.n0 63.321
R4772 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t3 333.651
R4773 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t2 297.233
R4774 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t4 294.554
R4775 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t5 211.008
R4776 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t1 102.408
R4777 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/D.t0 50.774
R4778 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D.n1 49.535
R4779 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/D 20.838
R4780 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D.n0 9.965
R4781 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D.n4 7.455
R4782 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n3 3.763
R4783 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n2 3.763
R4784 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[10]/D 2.855
R4785 sky130_fd_sc_hd__dfrbp_1_0[10]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[10]/D 1.297
R4786 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n0 163.71
R4787 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n1 82.083
R4788 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.t1 63.333
R4789 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.t3 63.321
R4790 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_448_47.t2 29.726
R4791 sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/Q.t0 59.048
R4792 sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/Q.t1 50.115
R4793 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1270_413.t1 126.642
R4794 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[10]/a_1217_47.t0 94.726
R4795 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t4 350.253
R4796 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t5 189.586
R4797 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n1 97.205
R4798 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t3 89.119
R4799 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n0 79.305
R4800 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n2 66.705
R4801 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t0 63.333
R4802 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n3 41.041
R4803 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_761_289.t1 31.979
R4804 sky130_fd_sc_hd__dfrbp_1_0[11]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_639_47.t0 198.571
R4805 sky130_fd_sc_hd__dfrbp_1_0[11]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_805_47.t1 60
R4806 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t6 389.181
R4807 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t3 256.987
R4808 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t8 212.079
R4809 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t7 174.888
R4810 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t4 163.801
R4811 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n0 161.578
R4812 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t5 139.779
R4813 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n1 129.263
R4814 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n5 102.015
R4815 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t1 63.321
R4816 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t2 63.321
R4817 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n6 46.071
R4818 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n3 37.442
R4819 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n4 23.54
R4820 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1283_21.n2 22.639
R4821 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.t3 239.038
R4822 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.t2 166.738
R4823 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n1 95.895
R4824 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.t0 71.217
R4825 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1847_47.n0 30.051
R4826 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t2 203.459
R4827 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t5 187.847
R4828 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t3 164.979
R4829 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t4 149.105
R4830 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t1 143.732
R4831 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n1 76
R4832 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n3 73.482
R4833 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n2 50.925
R4834 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_193_47.n0 41.551
R4835 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t4 366.855
R4836 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t5 174.055
R4837 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n0 117.298
R4838 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n1 77.111
R4839 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t1 70
R4840 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t3 68.011
R4841 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n3 63.321
R4842 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.t2 61.666
R4843 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1108_47.n2 57.017
R4844 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1462_47.t1 87.142
R4845 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t2 530.008
R4846 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t4 334.888
R4847 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t6 255.459
R4848 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t3 224.611
R4849 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t7 196.882
R4850 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t5 141.921
R4851 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n9 126.03
R4852 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.t0 99.672
R4853 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n1 92.562
R4854 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n0 44.57
R4855 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n2 38.638
R4856 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n6 15
R4857 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n8 15
R4858 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n4 13.653
R4859 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n7 3.182
R4860 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n3 1.366
R4861 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[11]/a_27_47.n5 1.326
R4862 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t5 332.579
R4863 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t4 168.699
R4864 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n1 104.381
R4865 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n0 101.869
R4866 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t3 96.154
R4867 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n2 92.648
R4868 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n3 65.666
R4869 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t2 65
R4870 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_543_47.t1 45
R4871 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.t1 194.654
R4872 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.t2 168.384
R4873 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_651_413.n0 63.321
R4874 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t3 333.651
R4875 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t2 297.233
R4876 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t4 294.554
R4877 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t5 211.008
R4878 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t1 102.408
R4879 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/D.t0 50.774
R4880 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[11]/D.n1 49.535
R4881 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/D 20.838
R4882 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[11]/D.n0 9.965
R4883 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[11]/D.n4 7.455
R4884 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n3 3.763
R4885 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n2 3.763
R4886 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[11]/D 2.855
R4887 sky130_fd_sc_hd__dfrbp_1_0[11]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[11]/D 1.297
R4888 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n0 163.71
R4889 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n1 82.083
R4890 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.t1 63.333
R4891 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.t3 63.321
R4892 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_448_47.t2 29.726
R4893 sky130_fd_sc_hd__dfrbp_1_0[11]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/Q.t0 59.048
R4894 sky130_fd_sc_hd__dfrbp_1_0[11]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/Q.t1 50.115
R4895 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1270_413.t1 126.642
R4896 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[11]/a_1217_47.t1 94.726
R4897 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t4 350.253
R4898 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t5 189.586
R4899 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n1 97.205
R4900 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t1 89.119
R4901 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n0 79.305
R4902 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n2 66.705
R4903 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t2 63.333
R4904 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n3 41.041
R4905 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_761_289.t0 31.979
R4906 sky130_fd_sc_hd__dfrbp_1_0[12]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_639_47.t0 198.571
R4907 sky130_fd_sc_hd__dfrbp_1_0[12]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_805_47.t1 60
R4908 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t6 389.181
R4909 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t3 256.987
R4910 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t8 212.079
R4911 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t7 174.888
R4912 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t4 163.801
R4913 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n5 161.578
R4914 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t5 139.779
R4915 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n0 129.263
R4916 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n3 102.015
R4917 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n6 63.321
R4918 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t2 63.321
R4919 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.t1 46.071
R4920 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n2 37.442
R4921 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n4 23.54
R4922 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1283_21.n1 22.639
R4923 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.t3 239.038
R4924 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.t2 166.738
R4925 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n1 95.895
R4926 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.t0 71.217
R4927 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1847_47.n0 30.051
R4928 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t2 203.459
R4929 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t5 187.847
R4930 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t3 164.979
R4931 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t4 149.105
R4932 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t0 143.732
R4933 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n1 76
R4934 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n3 73.482
R4935 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n2 50.925
R4936 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_193_47.n0 41.551
R4937 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t4 366.855
R4938 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t5 174.055
R4939 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n0 117.298
R4940 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n1 77.111
R4941 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t1 70
R4942 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n3 68.011
R4943 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t2 63.321
R4944 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.t3 61.666
R4945 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1108_47.n2 57.017
R4946 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1462_47.t1 87.142
R4947 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t2 530.008
R4948 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t4 334.888
R4949 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t6 255.459
R4950 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t3 224.611
R4951 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t7 196.882
R4952 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t5 141.921
R4953 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n9 126.03
R4954 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.t0 99.672
R4955 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n1 92.562
R4956 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n0 44.57
R4957 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n2 38.638
R4958 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n6 15
R4959 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n8 15
R4960 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n4 13.653
R4961 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n7 3.182
R4962 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n3 1.366
R4963 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[12]/a_27_47.n5 1.326
R4964 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t5 332.579
R4965 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t4 168.699
R4966 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n1 104.381
R4967 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n0 101.869
R4968 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t2 96.154
R4969 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n2 92.648
R4970 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n3 65.666
R4971 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t3 65
R4972 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_543_47.t0 45
R4973 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.t1 194.654
R4974 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.t2 168.384
R4975 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_651_413.n0 63.321
R4976 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t3 333.651
R4977 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t2 297.233
R4978 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t4 294.554
R4979 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t5 211.008
R4980 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t1 102.408
R4981 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/D.t0 50.774
R4982 sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D.n1 49.535
R4983 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/D 20.838
R4984 sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D.n0 9.965
R4985 sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D.n4 7.455
R4986 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n3 3.763
R4987 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n2 3.763
R4988 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[12]/D 2.855
R4989 sky130_fd_sc_hd__dfrbp_1_0[12]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/D 1.297
R4990 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n0 163.71
R4991 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.t2 82.083
R4992 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.t3 63.333
R4993 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.t1 63.321
R4994 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.t0 26.393
R4995 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n2 14.4
R4996 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[12]/a_448_47.n1 3.333
R4997 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/Q.t0 59.048
R4998 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/Q.t1 50.115
R4999 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1270_413.t1 126.642
R5000 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[12]/a_1217_47.t0 94.726
R5001 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t4 350.253
R5002 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t5 189.586
R5003 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n1 97.205
R5004 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t1 89.119
R5005 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n0 79.305
R5006 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n2 66.705
R5007 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t2 63.333
R5008 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n3 41.041
R5009 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_761_289.t3 31.979
R5010 sky130_fd_sc_hd__dfrbp_1_0[13]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_639_47.t0 198.571
R5011 sky130_fd_sc_hd__dfrbp_1_0[13]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_805_47.t1 60
R5012 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t6 389.181
R5013 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t3 256.987
R5014 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t8 212.079
R5015 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t7 174.888
R5016 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t4 163.801
R5017 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n5 161.578
R5018 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t5 139.779
R5019 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n0 129.263
R5020 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n3 102.015
R5021 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n6 63.321
R5022 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t2 63.321
R5023 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.t1 46.071
R5024 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n2 37.442
R5025 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n4 23.54
R5026 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1283_21.n1 22.639
R5027 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.t3 239.038
R5028 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.t2 166.738
R5029 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n1 95.895
R5030 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.t0 71.217
R5031 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1847_47.n0 30.051
R5032 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t2 203.459
R5033 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t5 187.847
R5034 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t3 164.979
R5035 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t4 149.105
R5036 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t0 143.732
R5037 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n1 76
R5038 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n3 73.482
R5039 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n2 50.925
R5040 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_193_47.n0 41.551
R5041 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t4 366.855
R5042 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t5 174.055
R5043 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n0 117.298
R5044 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n1 77.111
R5045 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t2 70
R5046 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n3 68.011
R5047 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t1 63.321
R5048 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.t3 61.666
R5049 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1108_47.n2 57.017
R5050 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1462_47.t1 87.142
R5051 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t2 530.008
R5052 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t4 334.888
R5053 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t6 255.459
R5054 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t3 224.611
R5055 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t7 196.882
R5056 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t5 141.921
R5057 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n9 126.03
R5058 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.t0 99.672
R5059 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n1 92.562
R5060 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n0 44.57
R5061 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n2 38.638
R5062 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n6 15
R5063 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n8 15
R5064 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n4 13.653
R5065 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n7 3.182
R5066 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n3 1.366
R5067 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[13]/a_27_47.n5 1.326
R5068 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t5 332.579
R5069 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t4 168.699
R5070 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n1 104.381
R5071 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n0 101.869
R5072 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t3 96.154
R5073 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n2 92.648
R5074 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n3 65.666
R5075 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t2 65
R5076 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_543_47.t0 45
R5077 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.t1 194.654
R5078 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.t2 168.384
R5079 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_651_413.n0 63.321
R5080 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t3 333.651
R5081 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t2 297.233
R5082 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t4 294.554
R5083 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t5 211.008
R5084 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t1 102.408
R5085 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/D.t0 50.774
R5086 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D.n1 49.535
R5087 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/D 20.838
R5088 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D.n0 9.965
R5089 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D.n4 7.455
R5090 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n3 3.763
R5091 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n2 3.763
R5092 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[13]/D 2.855
R5093 sky130_fd_sc_hd__dfrbp_1_0[13]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[13]/D 1.297
R5094 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n0 163.71
R5095 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n1 82.083
R5096 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.t1 63.333
R5097 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.t3 63.321
R5098 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_448_47.t2 29.726
R5099 sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/Q.t0 59.048
R5100 sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/Q.t1 50.115
R5101 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1270_413.t1 126.642
R5102 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[13]/a_1217_47.t1 94.726
R5103 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t4 350.253
R5104 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t5 189.586
R5105 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n1 97.205
R5106 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t3 89.119
R5107 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n0 79.305
R5108 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n2 66.705
R5109 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t2 63.333
R5110 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n3 41.041
R5111 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_761_289.t0 31.979
R5112 sky130_fd_sc_hd__dfrbp_1_0[14]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_639_47.t0 198.571
R5113 sky130_fd_sc_hd__dfrbp_1_0[14]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_805_47.t1 60
R5114 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t6 389.181
R5115 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t3 256.987
R5116 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t8 212.079
R5117 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t7 174.888
R5118 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t4 163.801
R5119 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n5 161.578
R5120 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t5 139.779
R5121 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n0 129.263
R5122 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n3 102.015
R5123 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n6 63.321
R5124 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t2 63.321
R5125 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.t1 46.071
R5126 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n2 37.442
R5127 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n4 23.54
R5128 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1283_21.n1 22.639
R5129 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.t3 239.038
R5130 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.t2 166.738
R5131 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n1 95.895
R5132 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.t0 71.217
R5133 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1847_47.n0 30.051
R5134 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t2 203.459
R5135 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t5 187.847
R5136 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t3 164.979
R5137 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t4 149.105
R5138 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t1 143.732
R5139 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n1 76
R5140 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n3 73.482
R5141 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n2 50.925
R5142 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_193_47.n0 41.551
R5143 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t4 366.855
R5144 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t5 174.055
R5145 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n0 117.298
R5146 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n1 77.111
R5147 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t2 70
R5148 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n3 68.011
R5149 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t3 63.321
R5150 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.t0 61.666
R5151 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1108_47.n2 57.017
R5152 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1462_47.t1 87.142
R5153 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t2 530.008
R5154 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t4 334.888
R5155 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t6 255.459
R5156 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t3 224.611
R5157 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t7 196.882
R5158 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t5 141.921
R5159 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n9 126.03
R5160 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.t0 99.672
R5161 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n1 92.562
R5162 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n0 44.57
R5163 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n2 38.638
R5164 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n6 15
R5165 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n8 15
R5166 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n4 13.653
R5167 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n7 3.182
R5168 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n3 1.366
R5169 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[14]/a_27_47.n5 1.326
R5170 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t5 332.579
R5171 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t4 168.699
R5172 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n1 104.381
R5173 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n0 101.869
R5174 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n3 96.154
R5175 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n2 92.648
R5176 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t2 65.666
R5177 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t1 65
R5178 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_543_47.t3 45
R5179 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.t1 194.654
R5180 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.t2 168.384
R5181 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_651_413.n0 63.321
R5182 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t3 333.651
R5183 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t2 297.233
R5184 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t4 294.554
R5185 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t5 211.008
R5186 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t1 102.408
R5187 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/D.t0 50.774
R5188 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D.n1 49.535
R5189 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/D 20.838
R5190 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D.n0 9.965
R5191 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D.n4 7.455
R5192 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n3 3.763
R5193 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n2 3.763
R5194 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[14]/D 2.855
R5195 sky130_fd_sc_hd__dfrbp_1_0[14]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/D 1.297
R5196 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n0 163.71
R5197 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.t3 82.083
R5198 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.t2 63.333
R5199 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.t1 63.321
R5200 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.t0 26.393
R5201 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n2 14.4
R5202 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[14]/a_448_47.n1 3.333
R5203 sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/Q.t0 59.048
R5204 sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/Q.t1 50.115
R5205 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1270_413.t1 126.642
R5206 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[14]/a_1217_47.t1 94.726
R5207 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t4 350.253
R5208 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t5 189.586
R5209 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n1 97.205
R5210 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t0 89.119
R5211 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n0 79.305
R5212 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n2 66.705
R5213 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t3 63.333
R5214 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n3 41.041
R5215 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_761_289.t1 31.979
R5216 sky130_fd_sc_hd__dfrbp_1_0[15]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_639_47.t0 198.571
R5217 sky130_fd_sc_hd__dfrbp_1_0[15]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_805_47.t1 60
R5218 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t6 389.181
R5219 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t3 256.987
R5220 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t8 212.079
R5221 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t7 174.888
R5222 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t4 163.801
R5223 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n0 161.578
R5224 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t5 139.779
R5225 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n1 129.263
R5226 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n5 102.015
R5227 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t1 63.321
R5228 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t2 63.321
R5229 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n6 46.071
R5230 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n3 37.442
R5231 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n4 23.54
R5232 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1283_21.n2 22.639
R5233 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.t3 239.038
R5234 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.t2 166.738
R5235 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n1 95.895
R5236 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.t0 71.217
R5237 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1847_47.n0 30.051
R5238 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t2 203.459
R5239 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t5 187.847
R5240 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t3 164.979
R5241 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t4 149.105
R5242 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t0 143.732
R5243 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n1 76
R5244 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n3 73.482
R5245 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n2 50.925
R5246 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_193_47.n0 41.551
R5247 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t4 366.855
R5248 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t5 174.055
R5249 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n0 117.298
R5250 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n1 77.111
R5251 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t2 70
R5252 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n3 68.011
R5253 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t3 63.321
R5254 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.t1 61.666
R5255 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1108_47.n2 57.017
R5256 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1462_47.t1 87.142
R5257 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t2 530.008
R5258 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t4 334.888
R5259 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t6 255.459
R5260 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t3 224.611
R5261 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t7 196.882
R5262 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t5 141.921
R5263 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n9 126.03
R5264 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.t0 99.672
R5265 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n1 92.562
R5266 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n0 44.57
R5267 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n2 38.638
R5268 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n6 15
R5269 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n8 15
R5270 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n4 13.653
R5271 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n7 3.182
R5272 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n3 1.366
R5273 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[15]/a_27_47.n5 1.326
R5274 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t5 332.579
R5275 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t4 168.699
R5276 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n1 104.381
R5277 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n0 101.869
R5278 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t3 96.154
R5279 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n2 92.648
R5280 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n3 65.666
R5281 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t2 65
R5282 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_543_47.t1 45
R5283 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.t1 194.654
R5284 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.t2 168.384
R5285 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_651_413.n0 63.321
R5286 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t3 333.651
R5287 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t2 297.233
R5288 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t4 294.554
R5289 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t5 211.008
R5290 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t1 102.408
R5291 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/D.t0 50.774
R5292 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D.n1 49.535
R5293 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/D 20.838
R5294 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D.n0 9.965
R5295 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D.n4 7.455
R5296 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n3 3.763
R5297 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n2 3.763
R5298 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[15]/D 2.855
R5299 sky130_fd_sc_hd__dfrbp_1_0[15]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[15]/D 1.297
R5300 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n0 163.71
R5301 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n1 82.083
R5302 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.t3 63.333
R5303 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.t2 63.321
R5304 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_448_47.t1 29.726
R5305 sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[15]/Q.t0 59.048
R5306 sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[15]/Q.t1 50.115
R5307 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1270_413.t1 126.642
R5308 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1217_47.t1 sky130_fd_sc_hd__dfrbp_1_0[15]/a_1217_47.t0 94.726
R5309 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t4 350.253
R5310 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t5 189.586
R5311 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n1 97.205
R5312 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t1 89.119
R5313 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n0 79.305
R5314 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n2 66.705
R5315 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t2 63.333
R5316 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n3 41.041
R5317 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_761_289.t3 31.979
R5318 sky130_fd_sc_hd__dfrbp_1_0[16]/a_639_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_639_47.t1 198.571
R5319 sky130_fd_sc_hd__dfrbp_1_0[16]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_805_47.t1 60
R5320 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t6 389.181
R5321 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t3 256.987
R5322 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t8 212.079
R5323 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t7 174.888
R5324 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t4 163.801
R5325 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n0 161.578
R5326 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t5 139.779
R5327 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n1 129.263
R5328 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n5 102.015
R5329 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t1 63.321
R5330 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t2 63.321
R5331 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n6 46.071
R5332 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n3 37.442
R5333 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n4 23.54
R5334 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1283_21.n2 22.639
R5335 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.t3 239.038
R5336 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.t2 166.738
R5337 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n1 95.895
R5338 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.t0 71.217
R5339 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1847_47.n0 30.051
R5340 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t2 203.459
R5341 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t5 187.847
R5342 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t3 164.979
R5343 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t4 149.105
R5344 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t0 143.732
R5345 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n1 76
R5346 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n3 73.482
R5347 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n2 50.925
R5348 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_193_47.n0 41.551
R5349 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t4 366.855
R5350 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t5 174.055
R5351 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n0 117.298
R5352 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n1 77.111
R5353 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t3 70
R5354 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n3 68.011
R5355 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t2 63.321
R5356 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.t1 61.666
R5357 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1108_47.n2 57.017
R5358 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1462_47.t1 87.142
R5359 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t2 530.008
R5360 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t4 334.888
R5361 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t6 255.459
R5362 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t3 224.611
R5363 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t7 196.882
R5364 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t5 141.921
R5365 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n9 126.03
R5366 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.t0 99.672
R5367 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n1 92.562
R5368 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n0 44.57
R5369 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n2 38.638
R5370 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n6 15
R5371 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n8 15
R5372 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n4 13.653
R5373 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n7 3.182
R5374 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n3 1.366
R5375 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[16]/a_27_47.n5 1.326
R5376 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t5 332.579
R5377 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t4 168.699
R5378 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n1 104.381
R5379 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n0 101.869
R5380 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n3 96.154
R5381 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n2 92.648
R5382 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t2 65.666
R5383 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t1 65
R5384 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_543_47.t3 45
R5385 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.n0 194.654
R5386 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.t2 168.384
R5387 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_651_413.t1 63.321
R5388 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t3 333.651
R5389 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t2 297.233
R5390 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t4 294.554
R5391 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t5 211.008
R5392 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t1 102.408
R5393 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t0 50.774
R5394 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D.n1 49.535
R5395 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/D 20.838
R5396 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D.n0 9.965
R5397 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D.n4 7.455
R5398 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n3 3.763
R5399 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n2 3.763
R5400 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[16]/D 2.855
R5401 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/D 1.297
R5402 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n0 163.71
R5403 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.t3 82.083
R5404 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.t0 63.333
R5405 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.t2 63.321
R5406 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.t1 26.393
R5407 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n3 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n2 14.4
R5408 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n2 sky130_fd_sc_hd__dfrbp_1_0[16]/a_448_47.n1 3.333
R5409 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/Q.t0 59.048
R5410 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/Q.t1 50.115
R5411 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1270_413.t1 126.642
R5412 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[16]/a_1217_47.t1 94.726
R5413 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t4 350.253
R5414 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t5 189.586
R5415 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n1 97.205
R5416 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t2 89.119
R5417 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n0 79.305
R5418 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n2 66.705
R5419 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t1 63.333
R5420 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n3 41.041
R5421 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_761_289.t0 31.979
R5422 sky130_fd_sc_hd__dfrbp_1_0[17]/a_639_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_639_47.t1 198.571
R5423 sky130_fd_sc_hd__dfrbp_1_0[17]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_805_47.t1 60
R5424 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t6 389.181
R5425 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t3 256.987
R5426 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t8 212.079
R5427 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t7 174.888
R5428 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t4 163.801
R5429 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n0 161.578
R5430 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t5 139.779
R5431 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n1 129.263
R5432 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n5 102.015
R5433 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t1 63.321
R5434 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t2 63.321
R5435 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n6 46.071
R5436 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n3 37.442
R5437 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n4 23.54
R5438 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1283_21.n2 22.639
R5439 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.t3 239.038
R5440 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.t2 166.738
R5441 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n1 95.895
R5442 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.t0 71.217
R5443 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1847_47.n0 30.051
R5444 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t2 203.459
R5445 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t5 187.847
R5446 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t3 164.979
R5447 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t4 149.105
R5448 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t1 143.732
R5449 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n1 76
R5450 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n3 73.482
R5451 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n2 50.925
R5452 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_193_47.n0 41.551
R5453 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t4 366.855
R5454 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t5 174.055
R5455 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n0 117.298
R5456 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n1 77.111
R5457 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t1 70
R5458 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t3 68.011
R5459 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n3 63.321
R5460 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.t0 61.666
R5461 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1108_47.n2 57.017
R5462 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1462_47.t1 87.142
R5463 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t2 530.008
R5464 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t4 334.888
R5465 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t6 255.459
R5466 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t3 224.611
R5467 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t7 196.882
R5468 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t5 141.921
R5469 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n9 126.03
R5470 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.t0 99.672
R5471 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n1 92.562
R5472 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n0 44.57
R5473 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n2 38.638
R5474 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n6 15
R5475 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n8 15
R5476 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n4 13.653
R5477 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n7 3.182
R5478 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n3 1.366
R5479 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[17]/a_27_47.n5 1.326
R5480 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t5 332.579
R5481 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t4 168.699
R5482 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n1 104.381
R5483 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n0 101.869
R5484 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n3 96.154
R5485 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n2 92.648
R5486 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t2 65.666
R5487 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t1 65
R5488 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_543_47.t3 45
R5489 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.t1 194.654
R5490 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.t2 168.384
R5491 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_651_413.n0 63.321
R5492 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t3 333.651
R5493 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t2 297.233
R5494 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t4 294.554
R5495 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t5 211.008
R5496 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t1 102.408
R5497 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/D.t0 50.774
R5498 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[17]/D.n1 49.535
R5499 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/D 20.838
R5500 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[17]/D.n0 9.965
R5501 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[17]/D.n4 7.455
R5502 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n3 3.763
R5503 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n2 3.763
R5504 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[17]/D 2.855
R5505 sky130_fd_sc_hd__dfrbp_1_0[17]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[17]/D 1.297
R5506 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n0 163.71
R5507 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.t1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n1 82.083
R5508 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.t0 63.333
R5509 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.t3 63.321
R5510 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_448_47.t2 29.726
R5511 sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[17]/Q.t0 59.048
R5512 sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[17]/Q.t1 50.115
R5513 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1270_413.t1 126.642
R5514 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[17]/a_1217_47.t1 94.726
R5515 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t4 350.253
R5516 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t5 189.586
R5517 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n1 97.205
R5518 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t2 89.119
R5519 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n0 79.305
R5520 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n2 66.705
R5521 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t0 63.333
R5522 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n3 41.041
R5523 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_761_289.t3 31.979
R5524 sky130_fd_sc_hd__dfrbp_1_0[18]/a_639_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_639_47.t1 198.571
R5525 sky130_fd_sc_hd__dfrbp_1_0[18]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_805_47.t1 60
R5526 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t6 389.181
R5527 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t3 256.987
R5528 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t8 212.079
R5529 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t7 174.888
R5530 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t4 163.801
R5531 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n0 161.578
R5532 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t5 139.779
R5533 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n1 129.263
R5534 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n5 102.015
R5535 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t1 63.321
R5536 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t2 63.321
R5537 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n6 46.071
R5538 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n3 37.442
R5539 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n4 23.54
R5540 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1283_21.n2 22.639
R5541 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.t3 239.038
R5542 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.t2 166.738
R5543 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n1 95.895
R5544 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.t0 71.217
R5545 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1847_47.n0 30.051
R5546 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t2 203.459
R5547 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t5 187.847
R5548 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t3 164.979
R5549 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t4 149.105
R5550 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t1 143.732
R5551 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n1 76
R5552 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n3 73.482
R5553 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n2 50.925
R5554 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_193_47.n0 41.551
R5555 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t4 366.855
R5556 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t5 174.055
R5557 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n0 117.298
R5558 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n1 77.111
R5559 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t0 70
R5560 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t3 68.011
R5561 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n3 63.321
R5562 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.t2 61.666
R5563 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1108_47.n2 57.017
R5564 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1462_47.t1 87.142
R5565 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t2 530.008
R5566 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t4 334.888
R5567 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t6 255.459
R5568 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t3 224.611
R5569 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t7 196.882
R5570 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t5 141.921
R5571 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n9 126.03
R5572 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.t0 99.672
R5573 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n1 92.562
R5574 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n0 44.57
R5575 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n2 38.638
R5576 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n6 15
R5577 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n8 15
R5578 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n4 13.653
R5579 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n7 3.182
R5580 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n3 1.366
R5581 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[18]/a_27_47.n5 1.326
R5582 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t5 332.579
R5583 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t4 168.699
R5584 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n1 104.381
R5585 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n0 101.869
R5586 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t2 96.154
R5587 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n2 92.648
R5588 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n3 65.666
R5589 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t3 65
R5590 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_543_47.t1 45
R5591 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.n0 194.654
R5592 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.t2 168.384
R5593 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_651_413.t1 63.321
R5594 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t3 333.651
R5595 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t2 297.233
R5596 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t4 294.554
R5597 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t5 211.008
R5598 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t1 102.408
R5599 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/D.t0 50.774
R5600 sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D.n1 49.535
R5601 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/D 20.838
R5602 sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D.n0 9.965
R5603 sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D.n4 7.455
R5604 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n3 3.763
R5605 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n3 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n2 3.763
R5606 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n4 sky130_fd_sc_hd__dfrbp_1_0[18]/D 2.855
R5607 sky130_fd_sc_hd__dfrbp_1_0[18]/D.n2 sky130_fd_sc_hd__dfrbp_1_0[18]/D 1.297
R5608 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n0 163.71
R5609 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n1 82.083
R5610 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.t1 63.333
R5611 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.t3 63.321
R5612 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_448_47.t2 29.726
R5613 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/Q.t0 59.048
R5614 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/Q.t1 50.115
R5615 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1270_413.t1 126.642
R5616 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[18]/a_1217_47.t1 94.726
R5617 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t4 350.253
R5618 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t5 189.586
R5619 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n1 97.205
R5620 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t3 89.119
R5621 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n0 79.305
R5622 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n2 66.705
R5623 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t2 63.333
R5624 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n3 41.041
R5625 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_761_289.t1 31.979
R5626 sky130_fd_sc_hd__dfrbp_1_0[19]/a_639_47.t1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_639_47.t0 198.571
R5627 sky130_fd_sc_hd__dfrbp_1_0[19]/a_805_47.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_805_47.t1 60
R5628 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t6 389.181
R5629 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t3 256.987
R5630 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t8 212.079
R5631 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n5 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t7 174.888
R5632 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t4 163.801
R5633 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n0 161.578
R5634 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t5 139.779
R5635 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n1 129.263
R5636 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n5 102.015
R5637 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t1 63.321
R5638 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t2 63.321
R5639 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n6 46.071
R5640 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n4 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n3 37.442
R5641 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n6 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n4 23.54
R5642 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1283_21.n2 22.639
R5643 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.t3 239.038
R5644 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.t2 166.738
R5645 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.t1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n1 95.895
R5646 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.t0 71.217
R5647 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1847_47.n0 30.051
R5648 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t2 203.459
R5649 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t5 187.847
R5650 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t3 164.979
R5651 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t4 149.105
R5652 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t0 143.732
R5653 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n1 76
R5654 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.t1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n3 73.482
R5655 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n2 50.925
R5656 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_193_47.n0 41.551
R5657 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t4 366.855
R5658 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t5 174.055
R5659 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n0 117.298
R5660 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n1 77.111
R5661 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t0 70
R5662 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t3 68.011
R5663 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n3 63.321
R5664 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.t2 61.666
R5665 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1108_47.n2 57.017
R5666 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1462_47.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1462_47.t1 87.142
R5667 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t2 530.008
R5668 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t4 334.888
R5669 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n8 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t6 255.459
R5670 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n4 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t3 224.611
R5671 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t7 196.882
R5672 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t5 141.921
R5673 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n9 126.03
R5674 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.t0 99.672
R5675 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n1 92.562
R5676 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n0 44.57
R5677 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n2 38.638
R5678 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n6 15
R5679 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n8 15
R5680 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n4 13.653
R5681 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n9 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n7 3.182
R5682 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n5 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n3 1.366
R5683 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n7 sky130_fd_sc_hd__dfrbp_1_0[19]/a_27_47.n5 1.326
R5684 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t5 332.579
R5685 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t4 168.699
R5686 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n1 104.381
R5687 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n2 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n0 101.869
R5688 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t3 96.154
R5689 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n3 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n2 92.648
R5690 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n3 65.666
R5691 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t2 65
R5692 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_543_47.t1 45
R5693 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.t1 194.654
R5694 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.t2 168.384
R5695 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_651_413.n0 63.321
R5696 sky130_fd_sc_hd__dfrbp_1_0[19]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/D.t3 333.651
R5697 sky130_fd_sc_hd__dfrbp_1_0[19]/D.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/D.t2 297.233
R5698 sky130_fd_sc_hd__dfrbp_1_0[19]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/D.t1 92.046
R5699 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[19]/D.t0 55.241
R5700 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[19]/D.n0 49.535
R5701 sky130_fd_sc_hd__dfrbp_1_0[19]/D.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/D 20.838
R5702 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[19]/D.n1 6.185
R5703 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n0 163.71
R5704 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n1 82.083
R5705 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.t3 63.333
R5706 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n1 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.t2 63.321
R5707 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.n0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_448_47.t1 29.726
R5708 sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/Q.t0 59.048
R5709 sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/Q.t1 50.115
R5710 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1270_413.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1270_413.t1 126.642
R5711 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1217_47.t0 sky130_fd_sc_hd__dfrbp_1_0[19]/a_1217_47.t1 94.726
Xsky130_fd_sc_hd__dfrbp_1_0[0] Vclk sky130_fd_sc_hd__dfrbp_1_0[0]/D
+ sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[1] sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[1]/D
+ sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[2] sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D
+ sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[3] sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D
+ sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[4] sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D
+ sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[4]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[5] sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D
+ sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[6] sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D
+ sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[7] sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D
+ sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[8] sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D
+ sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[8]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[9] sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D
+ sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[10] sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D
+ sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[11] sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[11]/D
+ sky130_fd_sc_hd__dfrbp_1_0[11]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[12] sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D
+ sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[13] sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D
+ sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[14] sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D
+ sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[15] sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D
+ sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[15]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[16] sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D
+ sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[17] sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[17]/D
+ sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[17]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[18] sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D
+ sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_0[19] sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[19]/D
+ sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/D Vreset
+ GND VDD sky130_fd_sc_hd__dfrbp_1
C77 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t4 0 0.04fF
C78 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t5 0 0.02fF
C79 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t2 0 0.03fF
C80 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t3 0 0.03fF
C81 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n1 0 0.08fF $ **FLOATING
C82 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n2 0 0.08fF $ **FLOATING
C83 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n3 0 1.31fF $ **FLOATING
C84 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n4 0 0.13fF $ **FLOATING
C85 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t4 0 0.04fF
C86 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t5 0 0.02fF
C87 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t2 0 0.03fF
C88 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t3 0 0.03fF
C89 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n1 0 0.08fF $ **FLOATING
C90 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n2 0 0.07fF $ **FLOATING
C91 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n3 0 1.31fF $ **FLOATING
C92 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n4 0 0.13fF $ **FLOATING
C93 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t4 0 0.04fF
C94 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t5 0 0.02fF
C95 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t2 0 0.03fF
C96 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t3 0 0.03fF
C97 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n1 0 0.08fF $ **FLOATING
C98 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n2 0 0.08fF $ **FLOATING
C99 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n3 0 1.31fF $ **FLOATING
C100 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n4 0 0.13fF $ **FLOATING
C101 VDD.t110 0 0.01fF
C102 VDD.t84 0 0.01fF
C103 VDD.t135 0 0.01fF
C104 VDD.t119 0 0.01fF
C105 VDD.t117 0 0.02fF
C106 VDD.t180 0 0.01fF
C107 VDD.t188 0 0.01fF
C108 VDD.t96 0 0.01fF
C109 VDD.t109 0 0.03fF
C110 VDD.t187 0 0.01fF
C111 VDD.t163 0 0.01fF
C112 VDD.t116 0 0.01fF
C113 VDD.n77 0 0.02fF $ **FLOATING
C114 VDD.n78 0 0.02fF $ **FLOATING
C115 VDD.n79 0 0.04fF $ **FLOATING
C116 VDD.n80 0 0.02fF $ **FLOATING
C117 VDD.n81 0 0.03fF $ **FLOATING
C118 VDD.n82 0 0.04fF $ **FLOATING
C119 VDD.n83 0 0.02fF $ **FLOATING
C120 VDD.n84 0 0.03fF $ **FLOATING
C121 VDD.n85 0 0.04fF $ **FLOATING
C122 VDD.t127 0 0.01fF
C123 VDD.t136 0 0.01fF
C124 VDD.n86 0 0.03fF $ **FLOATING
C125 VDD.n87 0 0.04fF $ **FLOATING
C126 VDD.n88 0 0.02fF $ **FLOATING
C127 VDD.n89 0 0.02fF $ **FLOATING
C128 VDD.n90 0 0.04fF $ **FLOATING
C129 VDD.n91 0 0.02fF $ **FLOATING
C130 VDD.n92 0 0.03fF $ **FLOATING
C131 VDD.n93 0 0.04fF $ **FLOATING
C132 VDD.n94 0 0.02fF $ **FLOATING
C133 VDD.n95 0 0.03fF $ **FLOATING
C134 VDD.n96 0 0.04fF $ **FLOATING
C135 VDD.t126 0 0.01fF
C136 VDD.t155 0 0.01fF
C137 VDD.n97 0 0.07fF $ **FLOATING
C138 VDD.n98 0 0.03fF $ **FLOATING
C139 VDD.n99 0 0.02fF $ **FLOATING
C140 VDD.n100 0 0.02fF $ **FLOATING
C141 VDD.n101 0 0.04fF $ **FLOATING
C142 VDD.n102 0 0.02fF $ **FLOATING
C143 VDD.n103 0 0.03fF $ **FLOATING
C144 VDD.n104 0 0.04fF $ **FLOATING
C145 VDD.n105 0 0.02fF $ **FLOATING
C146 VDD.n106 0 0.03fF $ **FLOATING
C147 VDD.n107 0 0.04fF $ **FLOATING
C148 VDD.n108 0 0.02fF $ **FLOATING
C149 VDD.n109 0 0.03fF $ **FLOATING
C150 VDD.n110 0 0.04fF $ **FLOATING
C151 VDD.t90 0 0.02fF
C152 VDD.n111 0 0.04fF $ **FLOATING
C153 VDD.n112 0 0.04fF $ **FLOATING
C154 VDD.t177 0 0.01fF
C155 VDD.n113 0 0.02fF $ **FLOATING
C156 VDD.n114 0 0.03fF $ **FLOATING
C157 VDD.n115 0 0.02fF $ **FLOATING
C158 VDD.n116 0 0.03fF $ **FLOATING
C159 VDD.n117 0 0.04fF $ **FLOATING
C160 VDD.n118 0 0.02fF $ **FLOATING
C161 VDD.n119 0 0.03fF $ **FLOATING
C162 VDD.n120 0 0.04fF $ **FLOATING
C163 VDD.t190 0 0.01fF
C164 VDD.t114 0 0.01fF
C165 VDD.n121 0 0.03fF $ **FLOATING
C166 VDD.n122 0 0.03fF $ **FLOATING
C167 VDD.n123 0 0.02fF $ **FLOATING
C168 VDD.n124 0 0.02fF $ **FLOATING
C169 VDD.n125 0 0.04fF $ **FLOATING
C170 VDD.n126 0 0.02fF $ **FLOATING
C171 VDD.n127 0 0.03fF $ **FLOATING
C172 VDD.n128 0 0.04fF $ **FLOATING
C173 VDD.n129 0 0.02fF $ **FLOATING
C174 VDD.n130 0 0.03fF $ **FLOATING
C175 VDD.n131 0 0.04fF $ **FLOATING
C176 VDD.n132 0 0.02fF $ **FLOATING
C177 VDD.n133 0 0.03fF $ **FLOATING
C178 VDD.n134 0 0.04fF $ **FLOATING
C179 VDD.t128 0 0.03fF
C180 VDD.n135 0 0.06fF $ **FLOATING
C181 VDD.n136 0 0.02fF $ **FLOATING
C182 VDD.n137 0 0.02fF $ **FLOATING
C183 VDD.n138 0 0.04fF $ **FLOATING
C184 VDD.n139 0 0.02fF $ **FLOATING
C185 VDD.n140 0 0.03fF $ **FLOATING
C186 VDD.n141 0 0.04fF $ **FLOATING
C187 VDD.t189 0 0.01fF
C188 VDD.t169 0 0.01fF
C189 VDD.n142 0 0.02fF $ **FLOATING
C190 VDD.n143 0 0.03fF $ **FLOATING
C191 VDD.n144 0 0.02fF $ **FLOATING
C192 VDD.n145 0 0.02fF $ **FLOATING
C193 VDD.n146 0 0.04fF $ **FLOATING
C194 VDD.n147 0 0.02fF $ **FLOATING
C195 VDD.n148 0 0.03fF $ **FLOATING
C196 VDD.n149 0 0.04fF $ **FLOATING
C197 VDD.n150 0 0.02fF $ **FLOATING
C198 VDD.n151 0 0.03fF $ **FLOATING
C199 VDD.n152 0 0.04fF $ **FLOATING
C200 VDD.n153 0 0.02fF $ **FLOATING
C201 VDD.n154 0 0.03fF $ **FLOATING
C202 VDD.n155 0 0.04fF $ **FLOATING
C203 VDD.n156 0 0.02fF $ **FLOATING
C204 VDD.n157 0 0.03fF $ **FLOATING
C205 VDD.n158 0 0.04fF $ **FLOATING
C206 VDD.t151 0 0.01fF
C207 VDD.n159 0 0.05fF $ **FLOATING
C208 VDD.n160 0 0.02fF $ **FLOATING
C209 VDD.n161 0 0.02fF $ **FLOATING
C210 VDD.n162 0 0.04fF $ **FLOATING
C211 VDD.n163 0 0.02fF $ **FLOATING
C212 VDD.n164 0 0.03fF $ **FLOATING
C213 VDD.n165 0 0.04fF $ **FLOATING
C214 VDD.n166 0 0.02fF $ **FLOATING
C215 VDD.n167 0 0.03fF $ **FLOATING
C216 VDD.n168 0 0.04fF $ **FLOATING
C217 VDD.t99 0 0.01fF
C218 VDD.t118 0 0.01fF
C219 VDD.n169 0 0.03fF $ **FLOATING
C220 VDD.n170 0 0.04fF $ **FLOATING
C221 VDD.n171 0 0.02fF $ **FLOATING
C222 VDD.n172 0 0.02fF $ **FLOATING
C223 VDD.n173 0 0.04fF $ **FLOATING
C224 VDD.n174 0 0.02fF $ **FLOATING
C225 VDD.n175 0 0.03fF $ **FLOATING
C226 VDD.n176 0 0.04fF $ **FLOATING
C227 VDD.n177 0 0.02fF $ **FLOATING
C228 VDD.n178 0 0.03fF $ **FLOATING
C229 VDD.n179 0 0.04fF $ **FLOATING
C230 VDD.t181 0 0.01fF
C231 VDD.t138 0 0.01fF
C232 VDD.n180 0 0.07fF $ **FLOATING
C233 VDD.n181 0 0.03fF $ **FLOATING
C234 VDD.n182 0 0.02fF $ **FLOATING
C235 VDD.n183 0 0.02fF $ **FLOATING
C236 VDD.n184 0 0.04fF $ **FLOATING
C237 VDD.n185 0 0.02fF $ **FLOATING
C238 VDD.n186 0 0.03fF $ **FLOATING
C239 VDD.n187 0 0.04fF $ **FLOATING
C240 VDD.n188 0 0.02fF $ **FLOATING
C241 VDD.n189 0 0.03fF $ **FLOATING
C242 VDD.n190 0 0.04fF $ **FLOATING
C243 VDD.n191 0 0.02fF $ **FLOATING
C244 VDD.n192 0 0.03fF $ **FLOATING
C245 VDD.n193 0 0.04fF $ **FLOATING
C246 VDD.t174 0 0.02fF
C247 VDD.n194 0 0.04fF $ **FLOATING
C248 VDD.n195 0 0.04fF $ **FLOATING
C249 VDD.t134 0 0.01fF
C250 VDD.n196 0 0.02fF $ **FLOATING
C251 VDD.n197 0 0.03fF $ **FLOATING
C252 VDD.n198 0 0.02fF $ **FLOATING
C253 VDD.n199 0 0.03fF $ **FLOATING
C254 VDD.n200 0 0.04fF $ **FLOATING
C255 VDD.n201 0 0.02fF $ **FLOATING
C256 VDD.n202 0 0.03fF $ **FLOATING
C257 VDD.n203 0 0.04fF $ **FLOATING
C258 VDD.t192 0 0.01fF
C259 VDD.t185 0 0.01fF
C260 VDD.n204 0 0.03fF $ **FLOATING
C261 VDD.n205 0 0.03fF $ **FLOATING
C262 VDD.n206 0 0.02fF $ **FLOATING
C263 VDD.n207 0 0.02fF $ **FLOATING
C264 VDD.n208 0 0.04fF $ **FLOATING
C265 VDD.n209 0 0.02fF $ **FLOATING
C266 VDD.n210 0 0.03fF $ **FLOATING
C267 VDD.n211 0 0.04fF $ **FLOATING
C268 VDD.n212 0 0.02fF $ **FLOATING
C269 VDD.n213 0 0.03fF $ **FLOATING
C270 VDD.n214 0 0.04fF $ **FLOATING
C271 VDD.n215 0 0.02fF $ **FLOATING
C272 VDD.n216 0 0.03fF $ **FLOATING
C273 VDD.n217 0 0.04fF $ **FLOATING
C274 VDD.t168 0 0.03fF
C275 VDD.n218 0 0.06fF $ **FLOATING
C276 VDD.n219 0 0.02fF $ **FLOATING
C277 VDD.n220 0 0.02fF $ **FLOATING
C278 VDD.n221 0 0.04fF $ **FLOATING
C279 VDD.n222 0 0.02fF $ **FLOATING
C280 VDD.n223 0 0.03fF $ **FLOATING
C281 VDD.n224 0 0.04fF $ **FLOATING
C282 VDD.t191 0 0.01fF
C283 VDD.t45 0 0.01fF
C284 VDD.n225 0 0.02fF $ **FLOATING
C285 VDD.n226 0 0.03fF $ **FLOATING
C286 VDD.n227 0 0.02fF $ **FLOATING
C287 VDD.n228 0 0.02fF $ **FLOATING
C288 VDD.n229 0 0.04fF $ **FLOATING
C289 VDD.n230 0 0.02fF $ **FLOATING
C290 VDD.n231 0 0.03fF $ **FLOATING
C291 VDD.n232 0 0.04fF $ **FLOATING
C292 VDD.n233 0 0.02fF $ **FLOATING
C293 VDD.n234 0 0.03fF $ **FLOATING
C294 VDD.n235 0 0.04fF $ **FLOATING
C295 VDD.n236 0 0.02fF $ **FLOATING
C296 VDD.n237 0 0.03fF $ **FLOATING
C297 VDD.n238 0 0.04fF $ **FLOATING
C298 VDD.n239 0 0.02fF $ **FLOATING
C299 VDD.n240 0 0.03fF $ **FLOATING
C300 VDD.n241 0 0.04fF $ **FLOATING
C301 VDD.t43 0 0.01fF
C302 VDD.n242 0 0.05fF $ **FLOATING
C303 VDD.n243 0 0.02fF $ **FLOATING
C304 VDD.n244 0 0.02fF $ **FLOATING
C305 VDD.n245 0 0.04fF $ **FLOATING
C306 VDD.n246 0 0.02fF $ **FLOATING
C307 VDD.n247 0 0.03fF $ **FLOATING
C308 VDD.n248 0 0.04fF $ **FLOATING
C309 VDD.n249 0 0.02fF $ **FLOATING
C310 VDD.n250 0 0.03fF $ **FLOATING
C311 VDD.n251 0 0.04fF $ **FLOATING
C312 VDD.t130 0 0.01fF
C313 VDD.t50 0 0.01fF
C314 VDD.n252 0 0.03fF $ **FLOATING
C315 VDD.n253 0 0.04fF $ **FLOATING
C316 VDD.n254 0 0.02fF $ **FLOATING
C317 VDD.n255 0 0.02fF $ **FLOATING
C318 VDD.n256 0 0.04fF $ **FLOATING
C319 VDD.n257 0 0.02fF $ **FLOATING
C320 VDD.n258 0 0.03fF $ **FLOATING
C321 VDD.n259 0 0.04fF $ **FLOATING
C322 VDD.n260 0 0.02fF $ **FLOATING
C323 VDD.n261 0 0.03fF $ **FLOATING
C324 VDD.n262 0 0.04fF $ **FLOATING
C325 VDD.t167 0 0.01fF
C326 VDD.t227 0 0.01fF
C327 VDD.n263 0 0.07fF $ **FLOATING
C328 VDD.n264 0 0.03fF $ **FLOATING
C329 VDD.n265 0 0.02fF $ **FLOATING
C330 VDD.n266 0 0.02fF $ **FLOATING
C331 VDD.n267 0 0.04fF $ **FLOATING
C332 VDD.n268 0 0.02fF $ **FLOATING
C333 VDD.n269 0 0.03fF $ **FLOATING
C334 VDD.n270 0 0.04fF $ **FLOATING
C335 VDD.n271 0 0.02fF $ **FLOATING
C336 VDD.n272 0 0.03fF $ **FLOATING
C337 VDD.n273 0 0.04fF $ **FLOATING
C338 VDD.n274 0 0.02fF $ **FLOATING
C339 VDD.n275 0 0.03fF $ **FLOATING
C340 VDD.n276 0 0.04fF $ **FLOATING
C341 VDD.t92 0 0.02fF
C342 VDD.n277 0 0.04fF $ **FLOATING
C343 VDD.n278 0 0.04fF $ **FLOATING
C344 VDD.t129 0 0.01fF
C345 VDD.n279 0 0.02fF $ **FLOATING
C346 VDD.n280 0 0.03fF $ **FLOATING
C347 VDD.n281 0 0.02fF $ **FLOATING
C348 VDD.n282 0 0.03fF $ **FLOATING
C349 VDD.n283 0 0.04fF $ **FLOATING
C350 VDD.n284 0 0.02fF $ **FLOATING
C351 VDD.n285 0 0.03fF $ **FLOATING
C352 VDD.n286 0 0.04fF $ **FLOATING
C353 VDD.t194 0 0.01fF
C354 VDD.t122 0 0.01fF
C355 VDD.n287 0 0.03fF $ **FLOATING
C356 VDD.n288 0 0.03fF $ **FLOATING
C357 VDD.n289 0 0.02fF $ **FLOATING
C358 VDD.n290 0 0.02fF $ **FLOATING
C359 VDD.n291 0 0.04fF $ **FLOATING
C360 VDD.n292 0 0.02fF $ **FLOATING
C361 VDD.n293 0 0.03fF $ **FLOATING
C362 VDD.n294 0 0.04fF $ **FLOATING
C363 VDD.n295 0 0.02fF $ **FLOATING
C364 VDD.n296 0 0.03fF $ **FLOATING
C365 VDD.n297 0 0.04fF $ **FLOATING
C366 VDD.n298 0 0.02fF $ **FLOATING
C367 VDD.n299 0 0.03fF $ **FLOATING
C368 VDD.n300 0 0.04fF $ **FLOATING
C369 VDD.t18 0 0.03fF
C370 VDD.n301 0 0.06fF $ **FLOATING
C371 VDD.n302 0 0.02fF $ **FLOATING
C372 VDD.n303 0 0.02fF $ **FLOATING
C373 VDD.n304 0 0.04fF $ **FLOATING
C374 VDD.n305 0 0.02fF $ **FLOATING
C375 VDD.n306 0 0.03fF $ **FLOATING
C376 VDD.n307 0 0.04fF $ **FLOATING
C377 VDD.t193 0 0.01fF
C378 VDD.t91 0 0.01fF
C379 VDD.n308 0 0.02fF $ **FLOATING
C380 VDD.n309 0 0.03fF $ **FLOATING
C381 VDD.n310 0 0.02fF $ **FLOATING
C382 VDD.n311 0 0.02fF $ **FLOATING
C383 VDD.n312 0 0.04fF $ **FLOATING
C384 VDD.n313 0 0.02fF $ **FLOATING
C385 VDD.n314 0 0.03fF $ **FLOATING
C386 VDD.n315 0 0.04fF $ **FLOATING
C387 VDD.n316 0 0.02fF $ **FLOATING
C388 VDD.n317 0 0.03fF $ **FLOATING
C389 VDD.n318 0 0.04fF $ **FLOATING
C390 VDD.n319 0 0.02fF $ **FLOATING
C391 VDD.n320 0 0.03fF $ **FLOATING
C392 VDD.n321 0 0.04fF $ **FLOATING
C393 VDD.n322 0 0.02fF $ **FLOATING
C394 VDD.n323 0 0.03fF $ **FLOATING
C395 VDD.n324 0 0.04fF $ **FLOATING
C396 VDD.t147 0 0.01fF
C397 VDD.n325 0 0.05fF $ **FLOATING
C398 VDD.n326 0 0.02fF $ **FLOATING
C399 VDD.n327 0 0.02fF $ **FLOATING
C400 VDD.n328 0 0.04fF $ **FLOATING
C401 VDD.n329 0 0.02fF $ **FLOATING
C402 VDD.n330 0 0.03fF $ **FLOATING
C403 VDD.n331 0 0.04fF $ **FLOATING
C404 VDD.n332 0 0.02fF $ **FLOATING
C405 VDD.n333 0 0.03fF $ **FLOATING
C406 VDD.n334 0 0.04fF $ **FLOATING
C407 VDD.t143 0 0.01fF
C408 VDD.t97 0 0.01fF
C409 VDD.n335 0 0.03fF $ **FLOATING
C410 VDD.n336 0 0.04fF $ **FLOATING
C411 VDD.n337 0 0.02fF $ **FLOATING
C412 VDD.n338 0 0.02fF $ **FLOATING
C413 VDD.n339 0 0.04fF $ **FLOATING
C414 VDD.n340 0 0.02fF $ **FLOATING
C415 VDD.n341 0 0.03fF $ **FLOATING
C416 VDD.n342 0 0.04fF $ **FLOATING
C417 VDD.n343 0 0.02fF $ **FLOATING
C418 VDD.n344 0 0.03fF $ **FLOATING
C419 VDD.n345 0 0.04fF $ **FLOATING
C420 VDD.t235 0 0.01fF
C421 VDD.t150 0 0.01fF
C422 VDD.n346 0 0.07fF $ **FLOATING
C423 VDD.n347 0 0.03fF $ **FLOATING
C424 VDD.n348 0 0.02fF $ **FLOATING
C425 VDD.n349 0 0.02fF $ **FLOATING
C426 VDD.n350 0 0.04fF $ **FLOATING
C427 VDD.n351 0 0.02fF $ **FLOATING
C428 VDD.n352 0 0.03fF $ **FLOATING
C429 VDD.n353 0 0.04fF $ **FLOATING
C430 VDD.n354 0 0.02fF $ **FLOATING
C431 VDD.n355 0 0.03fF $ **FLOATING
C432 VDD.n356 0 0.04fF $ **FLOATING
C433 VDD.n357 0 0.02fF $ **FLOATING
C434 VDD.n358 0 0.03fF $ **FLOATING
C435 VDD.n359 0 0.04fF $ **FLOATING
C436 VDD.t106 0 0.02fF
C437 VDD.n360 0 0.04fF $ **FLOATING
C438 VDD.n361 0 0.04fF $ **FLOATING
C439 VDD.t137 0 0.01fF
C440 VDD.n362 0 0.02fF $ **FLOATING
C441 VDD.n363 0 0.03fF $ **FLOATING
C442 VDD.n364 0 0.02fF $ **FLOATING
C443 VDD.n365 0 0.03fF $ **FLOATING
C444 VDD.n366 0 0.04fF $ **FLOATING
C445 VDD.n367 0 0.02fF $ **FLOATING
C446 VDD.n368 0 0.03fF $ **FLOATING
C447 VDD.n369 0 0.04fF $ **FLOATING
C448 VDD.t196 0 0.01fF
C449 VDD.n370 0 0.03fF $ **FLOATING
C450 VDD.n371 0 0.03fF $ **FLOATING
C451 VDD.n372 0 0.02fF $ **FLOATING
C452 VDD.n373 0 0.02fF $ **FLOATING
C453 VDD.n374 0 0.04fF $ **FLOATING
C454 VDD.n375 0 0.02fF $ **FLOATING
C455 VDD.n376 0 0.03fF $ **FLOATING
C456 VDD.n377 0 0.04fF $ **FLOATING
C457 VDD.n378 0 0.02fF $ **FLOATING
C458 VDD.n379 0 0.03fF $ **FLOATING
C459 VDD.n380 0 0.04fF $ **FLOATING
C460 VDD.n381 0 0.02fF $ **FLOATING
C461 VDD.n382 0 0.03fF $ **FLOATING
C462 VDD.n383 0 0.04fF $ **FLOATING
C463 VDD.t140 0 0.03fF
C464 VDD.n384 0 0.06fF $ **FLOATING
C465 VDD.n385 0 0.02fF $ **FLOATING
C466 VDD.n386 0 0.02fF $ **FLOATING
C467 VDD.n387 0 0.04fF $ **FLOATING
C468 VDD.n388 0 0.02fF $ **FLOATING
C469 VDD.n389 0 0.03fF $ **FLOATING
C470 VDD.n390 0 0.04fF $ **FLOATING
C471 VDD.t195 0 0.01fF
C472 VDD.t124 0 0.01fF
C473 VDD.n391 0 0.02fF $ **FLOATING
C474 VDD.n392 0 0.03fF $ **FLOATING
C475 VDD.n393 0 0.02fF $ **FLOATING
C476 VDD.n394 0 0.02fF $ **FLOATING
C477 VDD.n395 0 0.04fF $ **FLOATING
C478 VDD.n396 0 0.02fF $ **FLOATING
C479 VDD.n397 0 0.03fF $ **FLOATING
C480 VDD.n398 0 0.04fF $ **FLOATING
C481 VDD.n399 0 0.02fF $ **FLOATING
C482 VDD.n400 0 0.03fF $ **FLOATING
C483 VDD.n401 0 0.04fF $ **FLOATING
C484 VDD.n402 0 0.02fF $ **FLOATING
C485 VDD.n403 0 0.03fF $ **FLOATING
C486 VDD.n404 0 0.04fF $ **FLOATING
C487 VDD.n405 0 0.02fF $ **FLOATING
C488 VDD.n406 0 0.03fF $ **FLOATING
C489 VDD.n407 0 0.04fF $ **FLOATING
C490 VDD.t228 0 0.01fF
C491 VDD.n408 0 0.05fF $ **FLOATING
C492 VDD.n409 0 0.02fF $ **FLOATING
C493 VDD.n410 0 0.02fF $ **FLOATING
C494 VDD.n411 0 0.04fF $ **FLOATING
C495 VDD.n412 0 0.02fF $ **FLOATING
C496 VDD.n413 0 0.03fF $ **FLOATING
C497 VDD.n414 0 0.04fF $ **FLOATING
C498 VDD.n415 0 0.02fF $ **FLOATING
C499 VDD.n416 0 0.03fF $ **FLOATING
C500 VDD.n417 0 0.04fF $ **FLOATING
C501 VDD.t141 0 0.01fF
C502 VDD.t46 0 0.01fF
C503 VDD.n418 0 0.03fF $ **FLOATING
C504 VDD.n419 0 0.04fF $ **FLOATING
C505 VDD.n420 0 0.02fF $ **FLOATING
C506 VDD.n421 0 0.02fF $ **FLOATING
C507 VDD.n422 0 0.04fF $ **FLOATING
C508 VDD.n423 0 0.02fF $ **FLOATING
C509 VDD.n424 0 0.03fF $ **FLOATING
C510 VDD.n425 0 0.04fF $ **FLOATING
C511 VDD.n426 0 0.02fF $ **FLOATING
C512 VDD.n427 0 0.03fF $ **FLOATING
C513 VDD.n428 0 0.04fF $ **FLOATING
C514 VDD.t183 0 0.01fF
C515 VDD.t39 0 0.01fF
C516 VDD.n429 0 0.07fF $ **FLOATING
C517 VDD.n430 0 0.03fF $ **FLOATING
C518 VDD.n431 0 0.02fF $ **FLOATING
C519 VDD.n432 0 0.02fF $ **FLOATING
C520 VDD.n433 0 0.04fF $ **FLOATING
C521 VDD.n434 0 0.02fF $ **FLOATING
C522 VDD.n435 0 0.03fF $ **FLOATING
C523 VDD.n436 0 0.04fF $ **FLOATING
C524 VDD.n437 0 0.02fF $ **FLOATING
C525 VDD.n438 0 0.03fF $ **FLOATING
C526 VDD.n439 0 0.04fF $ **FLOATING
C527 VDD.n440 0 0.02fF $ **FLOATING
C528 VDD.n441 0 0.03fF $ **FLOATING
C529 VDD.n442 0 0.04fF $ **FLOATING
C530 VDD.t115 0 0.02fF
C531 VDD.n443 0 0.04fF $ **FLOATING
C532 VDD.n444 0 0.04fF $ **FLOATING
C533 VDD.t36 0 0.01fF
C534 VDD.n445 0 0.02fF $ **FLOATING
C535 VDD.n446 0 0.03fF $ **FLOATING
C536 VDD.n447 0 0.02fF $ **FLOATING
C537 VDD.n448 0 0.03fF $ **FLOATING
C538 VDD.n449 0 0.04fF $ **FLOATING
C539 VDD.n450 0 0.02fF $ **FLOATING
C540 VDD.n451 0 0.03fF $ **FLOATING
C541 VDD.n452 0 0.04fF $ **FLOATING
C542 VDD.t198 0 0.01fF
C543 VDD.t154 0 0.01fF
C544 VDD.n453 0 0.03fF $ **FLOATING
C545 VDD.n454 0 0.03fF $ **FLOATING
C546 VDD.n455 0 0.02fF $ **FLOATING
C547 VDD.n456 0 0.02fF $ **FLOATING
C548 VDD.n457 0 0.04fF $ **FLOATING
C549 VDD.n458 0 0.02fF $ **FLOATING
C550 VDD.n459 0 0.03fF $ **FLOATING
C551 VDD.n460 0 0.04fF $ **FLOATING
C552 VDD.n461 0 0.02fF $ **FLOATING
C553 VDD.n462 0 0.03fF $ **FLOATING
C554 VDD.n463 0 0.04fF $ **FLOATING
C555 VDD.n464 0 0.02fF $ **FLOATING
C556 VDD.n465 0 0.03fF $ **FLOATING
C557 VDD.n466 0 0.04fF $ **FLOATING
C558 VDD.t51 0 0.03fF
C559 VDD.n467 0 0.06fF $ **FLOATING
C560 VDD.n468 0 0.02fF $ **FLOATING
C561 VDD.n469 0 0.02fF $ **FLOATING
C562 VDD.n470 0 0.04fF $ **FLOATING
C563 VDD.n471 0 0.02fF $ **FLOATING
C564 VDD.n472 0 0.03fF $ **FLOATING
C565 VDD.n473 0 0.04fF $ **FLOATING
C566 VDD.t197 0 0.01fF
C567 VDD.t107 0 0.01fF
C568 VDD.n474 0 0.02fF $ **FLOATING
C569 VDD.n475 0 0.03fF $ **FLOATING
C570 VDD.n476 0 0.02fF $ **FLOATING
C571 VDD.n477 0 0.02fF $ **FLOATING
C572 VDD.n478 0 0.04fF $ **FLOATING
C573 VDD.n479 0 0.02fF $ **FLOATING
C574 VDD.n480 0 0.03fF $ **FLOATING
C575 VDD.n481 0 0.04fF $ **FLOATING
C576 VDD.n482 0 0.02fF $ **FLOATING
C577 VDD.n483 0 0.03fF $ **FLOATING
C578 VDD.n484 0 0.04fF $ **FLOATING
C579 VDD.n485 0 0.02fF $ **FLOATING
C580 VDD.n486 0 0.03fF $ **FLOATING
C581 VDD.n487 0 0.04fF $ **FLOATING
C582 VDD.n488 0 0.02fF $ **FLOATING
C583 VDD.n489 0 0.03fF $ **FLOATING
C584 VDD.n490 0 0.04fF $ **FLOATING
C585 VDD.t31 0 0.01fF
C586 VDD.n491 0 0.05fF $ **FLOATING
C587 VDD.n492 0 0.02fF $ **FLOATING
C588 VDD.n493 0 0.02fF $ **FLOATING
C589 VDD.n494 0 0.04fF $ **FLOATING
C590 VDD.n495 0 0.02fF $ **FLOATING
C591 VDD.n496 0 0.03fF $ **FLOATING
C592 VDD.n497 0 0.04fF $ **FLOATING
C593 VDD.n498 0 0.02fF $ **FLOATING
C594 VDD.n499 0 0.03fF $ **FLOATING
C595 VDD.n500 0 0.04fF $ **FLOATING
C596 VDD.t166 0 0.01fF
C597 VDD.t172 0 0.01fF
C598 VDD.n501 0 0.03fF $ **FLOATING
C599 VDD.n502 0 0.04fF $ **FLOATING
C600 VDD.n503 0 0.02fF $ **FLOATING
C601 VDD.n504 0 0.02fF $ **FLOATING
C602 VDD.n505 0 0.04fF $ **FLOATING
C603 VDD.n506 0 0.02fF $ **FLOATING
C604 VDD.n507 0 0.03fF $ **FLOATING
C605 VDD.n508 0 0.04fF $ **FLOATING
C606 VDD.n509 0 0.02fF $ **FLOATING
C607 VDD.n510 0 0.03fF $ **FLOATING
C608 VDD.n511 0 0.04fF $ **FLOATING
C609 VDD.t179 0 0.01fF
C610 VDD.t125 0 0.01fF
C611 VDD.n512 0 0.07fF $ **FLOATING
C612 VDD.n513 0 0.03fF $ **FLOATING
C613 VDD.n514 0 0.02fF $ **FLOATING
C614 VDD.n515 0 0.02fF $ **FLOATING
C615 VDD.n516 0 0.04fF $ **FLOATING
C616 VDD.n517 0 0.02fF $ **FLOATING
C617 VDD.n518 0 0.03fF $ **FLOATING
C618 VDD.n519 0 0.04fF $ **FLOATING
C619 VDD.n520 0 0.02fF $ **FLOATING
C620 VDD.n521 0 0.03fF $ **FLOATING
C621 VDD.n522 0 0.04fF $ **FLOATING
C622 VDD.n523 0 0.02fF $ **FLOATING
C623 VDD.n524 0 0.03fF $ **FLOATING
C624 VDD.n525 0 0.04fF $ **FLOATING
C625 VDD.t121 0 0.02fF
C626 VDD.n526 0 0.04fF $ **FLOATING
C627 VDD.n527 0 0.04fF $ **FLOATING
C628 VDD.t76 0 0.01fF
C629 VDD.n528 0 0.02fF $ **FLOATING
C630 VDD.n529 0 0.03fF $ **FLOATING
C631 VDD.n530 0 0.02fF $ **FLOATING
C632 VDD.n531 0 0.03fF $ **FLOATING
C633 VDD.n532 0 0.04fF $ **FLOATING
C634 VDD.n533 0 0.02fF $ **FLOATING
C635 VDD.n534 0 0.03fF $ **FLOATING
C636 VDD.n535 0 0.04fF $ **FLOATING
C637 VDD.t200 0 0.01fF
C638 VDD.t88 0 0.01fF
C639 VDD.n536 0 0.03fF $ **FLOATING
C640 VDD.n537 0 0.03fF $ **FLOATING
C641 VDD.n538 0 0.02fF $ **FLOATING
C642 VDD.n539 0 0.02fF $ **FLOATING
C643 VDD.n540 0 0.04fF $ **FLOATING
C644 VDD.n541 0 0.02fF $ **FLOATING
C645 VDD.n542 0 0.03fF $ **FLOATING
C646 VDD.n543 0 0.04fF $ **FLOATING
C647 VDD.n544 0 0.02fF $ **FLOATING
C648 VDD.n545 0 0.03fF $ **FLOATING
C649 VDD.n546 0 0.04fF $ **FLOATING
C650 VDD.n547 0 0.02fF $ **FLOATING
C651 VDD.n548 0 0.03fF $ **FLOATING
C652 VDD.n549 0 0.04fF $ **FLOATING
C653 VDD.t66 0 0.03fF
C654 VDD.n550 0 0.06fF $ **FLOATING
C655 VDD.n551 0 0.02fF $ **FLOATING
C656 VDD.n552 0 0.02fF $ **FLOATING
C657 VDD.n553 0 0.04fF $ **FLOATING
C658 VDD.n554 0 0.02fF $ **FLOATING
C659 VDD.n555 0 0.03fF $ **FLOATING
C660 VDD.n556 0 0.04fF $ **FLOATING
C661 VDD.t199 0 0.01fF
C662 VDD.t105 0 0.01fF
C663 VDD.n557 0 0.02fF $ **FLOATING
C664 VDD.n558 0 0.03fF $ **FLOATING
C665 VDD.n559 0 0.02fF $ **FLOATING
C666 VDD.n560 0 0.02fF $ **FLOATING
C667 VDD.n561 0 0.04fF $ **FLOATING
C668 VDD.n562 0 0.02fF $ **FLOATING
C669 VDD.n563 0 0.03fF $ **FLOATING
C670 VDD.n564 0 0.04fF $ **FLOATING
C671 VDD.n565 0 0.02fF $ **FLOATING
C672 VDD.n566 0 0.03fF $ **FLOATING
C673 VDD.n567 0 0.04fF $ **FLOATING
C674 VDD.n568 0 0.02fF $ **FLOATING
C675 VDD.n569 0 0.03fF $ **FLOATING
C676 VDD.n570 0 0.04fF $ **FLOATING
C677 VDD.n571 0 0.02fF $ **FLOATING
C678 VDD.n572 0 0.03fF $ **FLOATING
C679 VDD.n573 0 0.04fF $ **FLOATING
C680 VDD.n574 0 0.05fF $ **FLOATING
C681 VDD.n575 0 0.02fF $ **FLOATING
C682 VDD.n576 0 0.02fF $ **FLOATING
C683 VDD.n577 0 0.04fF $ **FLOATING
C684 VDD.n578 0 0.02fF $ **FLOATING
C685 VDD.n579 0 0.03fF $ **FLOATING
C686 VDD.n580 0 0.04fF $ **FLOATING
C687 VDD.n581 0 0.02fF $ **FLOATING
C688 VDD.n582 0 0.03fF $ **FLOATING
C689 VDD.n583 0 0.04fF $ **FLOATING
C690 VDD.t148 0 0.01fF
C691 VDD.t35 0 0.01fF
C692 VDD.n584 0 0.03fF $ **FLOATING
C693 VDD.n585 0 0.04fF $ **FLOATING
C694 VDD.n586 0 0.02fF $ **FLOATING
C695 VDD.n587 0 0.02fF $ **FLOATING
C696 VDD.n588 0 0.04fF $ **FLOATING
C697 VDD.n589 0 0.02fF $ **FLOATING
C698 VDD.n590 0 0.03fF $ **FLOATING
C699 VDD.n591 0 0.04fF $ **FLOATING
C700 VDD.n592 0 0.02fF $ **FLOATING
C701 VDD.n593 0 0.03fF $ **FLOATING
C702 VDD.n594 0 0.04fF $ **FLOATING
C703 VDD.t89 0 0.01fF
C704 VDD.t145 0 0.01fF
C705 VDD.n595 0 0.07fF $ **FLOATING
C706 VDD.n596 0 0.03fF $ **FLOATING
C707 VDD.n597 0 0.02fF $ **FLOATING
C708 VDD.n598 0 0.02fF $ **FLOATING
C709 VDD.n599 0 0.04fF $ **FLOATING
C710 VDD.n600 0 0.02fF $ **FLOATING
C711 VDD.n601 0 0.03fF $ **FLOATING
C712 VDD.n602 0 0.04fF $ **FLOATING
C713 VDD.n603 0 0.02fF $ **FLOATING
C714 VDD.n604 0 0.03fF $ **FLOATING
C715 VDD.n605 0 0.04fF $ **FLOATING
C716 VDD.n606 0 0.02fF $ **FLOATING
C717 VDD.n607 0 0.03fF $ **FLOATING
C718 VDD.n608 0 0.04fF $ **FLOATING
C719 VDD.t79 0 0.02fF
C720 VDD.n609 0 0.04fF $ **FLOATING
C721 VDD.n610 0 0.04fF $ **FLOATING
C722 VDD.t55 0 0.01fF
C723 VDD.n611 0 0.02fF $ **FLOATING
C724 VDD.n612 0 0.03fF $ **FLOATING
C725 VDD.n613 0 0.02fF $ **FLOATING
C726 VDD.n614 0 0.03fF $ **FLOATING
C727 VDD.n615 0 0.04fF $ **FLOATING
C728 VDD.n616 0 0.02fF $ **FLOATING
C729 VDD.n617 0 0.03fF $ **FLOATING
C730 VDD.n618 0 0.04fF $ **FLOATING
C731 VDD.t202 0 0.01fF
C732 VDD.t58 0 0.01fF
C733 VDD.n619 0 0.03fF $ **FLOATING
C734 VDD.n620 0 0.03fF $ **FLOATING
C735 VDD.n621 0 0.02fF $ **FLOATING
C736 VDD.n622 0 0.02fF $ **FLOATING
C737 VDD.n623 0 0.04fF $ **FLOATING
C738 VDD.n624 0 0.02fF $ **FLOATING
C739 VDD.n625 0 0.03fF $ **FLOATING
C740 VDD.n626 0 0.04fF $ **FLOATING
C741 VDD.n627 0 0.02fF $ **FLOATING
C742 VDD.n628 0 0.03fF $ **FLOATING
C743 VDD.n629 0 0.04fF $ **FLOATING
C744 VDD.n630 0 0.02fF $ **FLOATING
C745 VDD.n631 0 0.03fF $ **FLOATING
C746 VDD.n632 0 0.04fF $ **FLOATING
C747 VDD.t112 0 0.03fF
C748 VDD.n633 0 0.06fF $ **FLOATING
C749 VDD.n634 0 0.02fF $ **FLOATING
C750 VDD.n635 0 0.02fF $ **FLOATING
C751 VDD.n636 0 0.04fF $ **FLOATING
C752 VDD.n637 0 0.02fF $ **FLOATING
C753 VDD.n638 0 0.03fF $ **FLOATING
C754 VDD.n639 0 0.04fF $ **FLOATING
C755 VDD.t201 0 0.01fF
C756 VDD.t186 0 0.01fF
C757 VDD.n640 0 0.02fF $ **FLOATING
C758 VDD.n641 0 0.03fF $ **FLOATING
C759 VDD.n642 0 0.02fF $ **FLOATING
C760 VDD.n643 0 0.02fF $ **FLOATING
C761 VDD.n644 0 0.04fF $ **FLOATING
C762 VDD.n645 0 0.02fF $ **FLOATING
C763 VDD.n646 0 0.03fF $ **FLOATING
C764 VDD.n647 0 0.04fF $ **FLOATING
C765 VDD.n648 0 0.02fF $ **FLOATING
C766 VDD.n649 0 0.03fF $ **FLOATING
C767 VDD.n650 0 0.04fF $ **FLOATING
C768 VDD.n651 0 0.02fF $ **FLOATING
C769 VDD.n652 0 0.03fF $ **FLOATING
C770 VDD.n653 0 0.04fF $ **FLOATING
C771 VDD.n654 0 0.02fF $ **FLOATING
C772 VDD.n655 0 0.03fF $ **FLOATING
C773 VDD.n656 0 0.04fF $ **FLOATING
C774 VDD.t94 0 0.01fF
C775 VDD.n657 0 0.05fF $ **FLOATING
C776 VDD.n658 0 0.02fF $ **FLOATING
C777 VDD.n659 0 0.02fF $ **FLOATING
C778 VDD.n660 0 0.04fF $ **FLOATING
C779 VDD.n661 0 0.02fF $ **FLOATING
C780 VDD.n662 0 0.03fF $ **FLOATING
C781 VDD.n663 0 0.04fF $ **FLOATING
C782 VDD.n664 0 0.02fF $ **FLOATING
C783 VDD.n665 0 0.03fF $ **FLOATING
C784 VDD.n666 0 0.04fF $ **FLOATING
C785 VDD.t233 0 0.01fF
C786 VDD.t72 0 0.01fF
C787 VDD.n667 0 0.03fF $ **FLOATING
C788 VDD.n668 0 0.04fF $ **FLOATING
C789 VDD.n669 0 0.02fF $ **FLOATING
C790 VDD.n670 0 0.02fF $ **FLOATING
C791 VDD.n671 0 0.04fF $ **FLOATING
C792 VDD.n672 0 0.02fF $ **FLOATING
C793 VDD.n673 0 0.03fF $ **FLOATING
C794 VDD.n674 0 0.04fF $ **FLOATING
C795 VDD.n675 0 0.02fF $ **FLOATING
C796 VDD.n676 0 0.03fF $ **FLOATING
C797 VDD.n677 0 0.04fF $ **FLOATING
C798 VDD.t170 0 0.01fF
C799 VDD.t152 0 0.01fF
C800 VDD.n678 0 0.07fF $ **FLOATING
C801 VDD.n679 0 0.03fF $ **FLOATING
C802 VDD.n680 0 0.02fF $ **FLOATING
C803 VDD.n681 0 0.02fF $ **FLOATING
C804 VDD.n682 0 0.04fF $ **FLOATING
C805 VDD.n683 0 0.02fF $ **FLOATING
C806 VDD.n684 0 0.03fF $ **FLOATING
C807 VDD.n685 0 0.04fF $ **FLOATING
C808 VDD.n686 0 0.02fF $ **FLOATING
C809 VDD.n687 0 0.03fF $ **FLOATING
C810 VDD.n688 0 0.04fF $ **FLOATING
C811 VDD.n689 0 0.02fF $ **FLOATING
C812 VDD.n690 0 0.03fF $ **FLOATING
C813 VDD.n691 0 0.04fF $ **FLOATING
C814 VDD.t16 0 0.02fF
C815 VDD.n692 0 0.04fF $ **FLOATING
C816 VDD.n693 0 0.04fF $ **FLOATING
C817 VDD.t173 0 0.01fF
C818 VDD.n694 0 0.02fF $ **FLOATING
C819 VDD.n695 0 0.03fF $ **FLOATING
C820 VDD.n696 0 0.02fF $ **FLOATING
C821 VDD.n697 0 0.03fF $ **FLOATING
C822 VDD.n698 0 0.04fF $ **FLOATING
C823 VDD.n699 0 0.02fF $ **FLOATING
C824 VDD.n700 0 0.03fF $ **FLOATING
C825 VDD.n701 0 0.04fF $ **FLOATING
C826 VDD.t204 0 0.01fF
C827 VDD.t87 0 0.01fF
C828 VDD.n702 0 0.03fF $ **FLOATING
C829 VDD.n703 0 0.03fF $ **FLOATING
C830 VDD.n704 0 0.02fF $ **FLOATING
C831 VDD.n705 0 0.02fF $ **FLOATING
C832 VDD.n706 0 0.04fF $ **FLOATING
C833 VDD.n707 0 0.02fF $ **FLOATING
C834 VDD.n708 0 0.03fF $ **FLOATING
C835 VDD.n709 0 0.04fF $ **FLOATING
C836 VDD.n710 0 0.02fF $ **FLOATING
C837 VDD.n711 0 0.03fF $ **FLOATING
C838 VDD.n712 0 0.04fF $ **FLOATING
C839 VDD.n713 0 0.02fF $ **FLOATING
C840 VDD.n714 0 0.03fF $ **FLOATING
C841 VDD.n715 0 0.04fF $ **FLOATING
C842 VDD.t101 0 0.03fF
C843 VDD.n716 0 0.06fF $ **FLOATING
C844 VDD.n717 0 0.02fF $ **FLOATING
C845 VDD.n718 0 0.02fF $ **FLOATING
C846 VDD.n719 0 0.04fF $ **FLOATING
C847 VDD.n720 0 0.02fF $ **FLOATING
C848 VDD.n721 0 0.03fF $ **FLOATING
C849 VDD.n722 0 0.04fF $ **FLOATING
C850 VDD.t203 0 0.01fF
C851 VDD.t40 0 0.01fF
C852 VDD.n723 0 0.02fF $ **FLOATING
C853 VDD.n724 0 0.03fF $ **FLOATING
C854 VDD.n725 0 0.02fF $ **FLOATING
C855 VDD.n726 0 0.02fF $ **FLOATING
C856 VDD.n727 0 0.04fF $ **FLOATING
C857 VDD.n728 0 0.02fF $ **FLOATING
C858 VDD.n729 0 0.03fF $ **FLOATING
C859 VDD.n730 0 0.04fF $ **FLOATING
C860 VDD.n731 0 0.02fF $ **FLOATING
C861 VDD.n732 0 0.03fF $ **FLOATING
C862 VDD.n733 0 0.04fF $ **FLOATING
C863 VDD.n734 0 0.02fF $ **FLOATING
C864 VDD.n735 0 0.03fF $ **FLOATING
C865 VDD.n736 0 0.04fF $ **FLOATING
C866 VDD.n737 0 0.02fF $ **FLOATING
C867 VDD.n738 0 0.03fF $ **FLOATING
C868 VDD.n739 0 0.04fF $ **FLOATING
C869 VDD.t81 0 0.01fF
C870 VDD.n740 0 0.05fF $ **FLOATING
C871 VDD.n741 0 0.02fF $ **FLOATING
C872 VDD.n742 0 0.02fF $ **FLOATING
C873 VDD.n743 0 0.04fF $ **FLOATING
C874 VDD.n744 0 0.02fF $ **FLOATING
C875 VDD.n745 0 0.03fF $ **FLOATING
C876 VDD.n746 0 0.04fF $ **FLOATING
C877 VDD.n747 0 0.02fF $ **FLOATING
C878 VDD.n748 0 0.03fF $ **FLOATING
C879 VDD.n749 0 0.04fF $ **FLOATING
C880 VDD.t120 0 0.01fF
C881 VDD.t61 0 0.01fF
C882 VDD.n750 0 0.03fF $ **FLOATING
C883 VDD.n751 0 0.04fF $ **FLOATING
C884 VDD.n752 0 0.02fF $ **FLOATING
C885 VDD.n753 0 0.02fF $ **FLOATING
C886 VDD.n754 0 0.04fF $ **FLOATING
C887 VDD.n755 0 0.02fF $ **FLOATING
C888 VDD.n756 0 0.03fF $ **FLOATING
C889 VDD.n757 0 0.04fF $ **FLOATING
C890 VDD.n758 0 0.02fF $ **FLOATING
C891 VDD.n759 0 0.03fF $ **FLOATING
C892 VDD.n760 0 0.04fF $ **FLOATING
C893 VDD.t73 0 0.01fF
C894 VDD.t95 0 0.01fF
C895 VDD.n761 0 0.07fF $ **FLOATING
C896 VDD.n762 0 0.03fF $ **FLOATING
C897 VDD.n763 0 0.02fF $ **FLOATING
C898 VDD.n764 0 0.02fF $ **FLOATING
C899 VDD.n765 0 0.04fF $ **FLOATING
C900 VDD.n766 0 0.02fF $ **FLOATING
C901 VDD.n767 0 0.03fF $ **FLOATING
C902 VDD.n768 0 0.04fF $ **FLOATING
C903 VDD.n769 0 0.02fF $ **FLOATING
C904 VDD.n770 0 0.03fF $ **FLOATING
C905 VDD.n771 0 0.04fF $ **FLOATING
C906 VDD.n772 0 0.02fF $ **FLOATING
C907 VDD.n773 0 0.03fF $ **FLOATING
C908 VDD.n774 0 0.04fF $ **FLOATING
C909 VDD.t108 0 0.02fF
C910 VDD.n775 0 0.04fF $ **FLOATING
C911 VDD.n776 0 0.04fF $ **FLOATING
C912 VDD.t15 0 0.01fF
C913 VDD.n777 0 0.02fF $ **FLOATING
C914 VDD.n778 0 0.03fF $ **FLOATING
C915 VDD.n779 0 0.02fF $ **FLOATING
C916 VDD.n780 0 0.03fF $ **FLOATING
C917 VDD.n781 0 0.04fF $ **FLOATING
C918 VDD.n782 0 0.02fF $ **FLOATING
C919 VDD.n783 0 0.03fF $ **FLOATING
C920 VDD.n784 0 0.04fF $ **FLOATING
C921 VDD.t206 0 0.01fF
C922 VDD.t69 0 0.01fF
C923 VDD.n785 0 0.03fF $ **FLOATING
C924 VDD.n786 0 0.03fF $ **FLOATING
C925 VDD.n787 0 0.02fF $ **FLOATING
C926 VDD.n788 0 0.02fF $ **FLOATING
C927 VDD.n789 0 0.04fF $ **FLOATING
C928 VDD.n790 0 0.02fF $ **FLOATING
C929 VDD.n791 0 0.03fF $ **FLOATING
C930 VDD.n792 0 0.04fF $ **FLOATING
C931 VDD.n793 0 0.02fF $ **FLOATING
C932 VDD.n794 0 0.03fF $ **FLOATING
C933 VDD.n795 0 0.04fF $ **FLOATING
C934 VDD.n796 0 0.02fF $ **FLOATING
C935 VDD.n797 0 0.03fF $ **FLOATING
C936 VDD.n798 0 0.04fF $ **FLOATING
C937 VDD.t164 0 0.03fF
C938 VDD.n799 0 0.06fF $ **FLOATING
C939 VDD.n800 0 0.02fF $ **FLOATING
C940 VDD.n801 0 0.02fF $ **FLOATING
C941 VDD.n802 0 0.04fF $ **FLOATING
C942 VDD.n803 0 0.02fF $ **FLOATING
C943 VDD.n804 0 0.03fF $ **FLOATING
C944 VDD.n805 0 0.04fF $ **FLOATING
C945 VDD.t205 0 0.01fF
C946 VDD.t32 0 0.01fF
C947 VDD.n806 0 0.02fF $ **FLOATING
C948 VDD.n807 0 0.03fF $ **FLOATING
C949 VDD.n808 0 0.02fF $ **FLOATING
C950 VDD.n809 0 0.02fF $ **FLOATING
C951 VDD.n810 0 0.04fF $ **FLOATING
C952 VDD.n811 0 0.02fF $ **FLOATING
C953 VDD.n812 0 0.03fF $ **FLOATING
C954 VDD.n813 0 0.04fF $ **FLOATING
C955 VDD.n814 0 0.02fF $ **FLOATING
C956 VDD.n815 0 0.03fF $ **FLOATING
C957 VDD.n816 0 0.04fF $ **FLOATING
C958 VDD.n817 0 0.02fF $ **FLOATING
C959 VDD.n818 0 0.03fF $ **FLOATING
C960 VDD.n819 0 0.04fF $ **FLOATING
C961 VDD.n820 0 0.02fF $ **FLOATING
C962 VDD.n821 0 0.03fF $ **FLOATING
C963 VDD.n822 0 0.04fF $ **FLOATING
C964 VDD.t111 0 0.01fF
C965 VDD.n823 0 0.05fF $ **FLOATING
C966 VDD.n824 0 0.02fF $ **FLOATING
C967 VDD.n825 0 0.02fF $ **FLOATING
C968 VDD.n826 0 0.04fF $ **FLOATING
C969 VDD.n827 0 0.02fF $ **FLOATING
C970 VDD.n828 0 0.03fF $ **FLOATING
C971 VDD.n829 0 0.04fF $ **FLOATING
C972 VDD.n830 0 0.02fF $ **FLOATING
C973 VDD.n831 0 0.03fF $ **FLOATING
C974 VDD.n832 0 0.04fF $ **FLOATING
C975 VDD.t229 0 0.01fF
C976 VDD.n833 0 0.03fF $ **FLOATING
C977 VDD.n834 0 0.04fF $ **FLOATING
C978 VDD.n835 0 0.02fF $ **FLOATING
C979 VDD.n836 0 0.02fF $ **FLOATING
C980 VDD.n837 0 0.04fF $ **FLOATING
C981 VDD.n838 0 0.02fF $ **FLOATING
C982 VDD.n839 0 0.03fF $ **FLOATING
C983 VDD.n840 0 0.04fF $ **FLOATING
C984 VDD.n841 0 0.02fF $ **FLOATING
C985 VDD.n842 0 0.03fF $ **FLOATING
C986 VDD.n843 0 0.04fF $ **FLOATING
C987 VDD.t171 0 0.01fF
C988 VDD.t48 0 0.01fF
C989 VDD.n844 0 0.07fF $ **FLOATING
C990 VDD.n845 0 0.03fF $ **FLOATING
C991 VDD.n846 0 0.02fF $ **FLOATING
C992 VDD.n847 0 0.02fF $ **FLOATING
C993 VDD.n848 0 0.04fF $ **FLOATING
C994 VDD.n849 0 0.02fF $ **FLOATING
C995 VDD.n850 0 0.03fF $ **FLOATING
C996 VDD.n851 0 0.04fF $ **FLOATING
C997 VDD.n852 0 0.02fF $ **FLOATING
C998 VDD.n853 0 0.03fF $ **FLOATING
C999 VDD.n854 0 0.04fF $ **FLOATING
C1000 VDD.n855 0 0.02fF $ **FLOATING
C1001 VDD.n856 0 0.03fF $ **FLOATING
C1002 VDD.n857 0 0.04fF $ **FLOATING
C1003 VDD.t149 0 0.02fF
C1004 VDD.n858 0 0.04fF $ **FLOATING
C1005 VDD.n859 0 0.04fF $ **FLOATING
C1006 VDD.t142 0 0.01fF
C1007 VDD.n860 0 0.02fF $ **FLOATING
C1008 VDD.n861 0 0.03fF $ **FLOATING
C1009 VDD.n862 0 0.02fF $ **FLOATING
C1010 VDD.n863 0 0.03fF $ **FLOATING
C1011 VDD.n864 0 0.04fF $ **FLOATING
C1012 VDD.n865 0 0.02fF $ **FLOATING
C1013 VDD.n866 0 0.03fF $ **FLOATING
C1014 VDD.n867 0 0.04fF $ **FLOATING
C1015 VDD.t208 0 0.01fF
C1016 VDD.t146 0 0.01fF
C1017 VDD.n868 0 0.03fF $ **FLOATING
C1018 VDD.n869 0 0.03fF $ **FLOATING
C1019 VDD.n870 0 0.02fF $ **FLOATING
C1020 VDD.n871 0 0.02fF $ **FLOATING
C1021 VDD.n872 0 0.04fF $ **FLOATING
C1022 VDD.n873 0 0.02fF $ **FLOATING
C1023 VDD.n874 0 0.03fF $ **FLOATING
C1024 VDD.n875 0 0.04fF $ **FLOATING
C1025 VDD.n876 0 0.02fF $ **FLOATING
C1026 VDD.n877 0 0.03fF $ **FLOATING
C1027 VDD.n878 0 0.04fF $ **FLOATING
C1028 VDD.n879 0 0.02fF $ **FLOATING
C1029 VDD.n880 0 0.03fF $ **FLOATING
C1030 VDD.n881 0 0.04fF $ **FLOATING
C1031 VDD.t49 0 0.03fF
C1032 VDD.n882 0 0.06fF $ **FLOATING
C1033 VDD.n883 0 0.02fF $ **FLOATING
C1034 VDD.n884 0 0.02fF $ **FLOATING
C1035 VDD.n885 0 0.04fF $ **FLOATING
C1036 VDD.n886 0 0.02fF $ **FLOATING
C1037 VDD.n887 0 0.03fF $ **FLOATING
C1038 VDD.n888 0 0.04fF $ **FLOATING
C1039 VDD.t207 0 0.01fF
C1040 VDD.t93 0 0.01fF
C1041 VDD.n889 0 0.02fF $ **FLOATING
C1042 VDD.n890 0 0.03fF $ **FLOATING
C1043 VDD.n891 0 0.02fF $ **FLOATING
C1044 VDD.n892 0 0.02fF $ **FLOATING
C1045 VDD.n893 0 0.04fF $ **FLOATING
C1046 VDD.n894 0 0.02fF $ **FLOATING
C1047 VDD.n895 0 0.03fF $ **FLOATING
C1048 VDD.n896 0 0.04fF $ **FLOATING
C1049 VDD.n897 0 0.02fF $ **FLOATING
C1050 VDD.n898 0 0.03fF $ **FLOATING
C1051 VDD.n899 0 0.04fF $ **FLOATING
C1052 VDD.n900 0 0.02fF $ **FLOATING
C1053 VDD.n901 0 0.03fF $ **FLOATING
C1054 VDD.n902 0 0.04fF $ **FLOATING
C1055 VDD.n903 0 0.02fF $ **FLOATING
C1056 VDD.n904 0 0.03fF $ **FLOATING
C1057 VDD.n905 0 0.04fF $ **FLOATING
C1058 VDD.t176 0 0.01fF
C1059 VDD.n906 0 0.05fF $ **FLOATING
C1060 VDD.n907 0 0.02fF $ **FLOATING
C1061 VDD.n908 0 0.02fF $ **FLOATING
C1062 VDD.n909 0 0.04fF $ **FLOATING
C1063 VDD.n910 0 0.02fF $ **FLOATING
C1064 VDD.n911 0 0.03fF $ **FLOATING
C1065 VDD.n912 0 0.04fF $ **FLOATING
C1066 VDD.n913 0 0.02fF $ **FLOATING
C1067 VDD.n914 0 0.03fF $ **FLOATING
C1068 VDD.n915 0 0.04fF $ **FLOATING
C1069 VDD.t153 0 0.01fF
C1070 VDD.t161 0 0.01fF
C1071 VDD.n916 0 0.03fF $ **FLOATING
C1072 VDD.n917 0 0.04fF $ **FLOATING
C1073 VDD.n918 0 0.02fF $ **FLOATING
C1074 VDD.n919 0 0.02fF $ **FLOATING
C1075 VDD.n920 0 0.04fF $ **FLOATING
C1076 VDD.n921 0 0.02fF $ **FLOATING
C1077 VDD.n922 0 0.03fF $ **FLOATING
C1078 VDD.n923 0 0.04fF $ **FLOATING
C1079 VDD.n924 0 0.02fF $ **FLOATING
C1080 VDD.n925 0 0.03fF $ **FLOATING
C1081 VDD.n926 0 0.04fF $ **FLOATING
C1082 VDD.t230 0 0.01fF
C1083 VDD.t162 0 0.01fF
C1084 VDD.n927 0 0.07fF $ **FLOATING
C1085 VDD.n928 0 0.03fF $ **FLOATING
C1086 VDD.n929 0 0.02fF $ **FLOATING
C1087 VDD.n930 0 0.02fF $ **FLOATING
C1088 VDD.n931 0 0.04fF $ **FLOATING
C1089 VDD.n932 0 0.02fF $ **FLOATING
C1090 VDD.n933 0 0.03fF $ **FLOATING
C1091 VDD.n934 0 0.04fF $ **FLOATING
C1092 VDD.n935 0 0.02fF $ **FLOATING
C1093 VDD.n936 0 0.03fF $ **FLOATING
C1094 VDD.n937 0 0.04fF $ **FLOATING
C1095 VDD.n938 0 0.02fF $ **FLOATING
C1096 VDD.n939 0 0.03fF $ **FLOATING
C1097 VDD.n940 0 0.04fF $ **FLOATING
C1098 VDD.n941 0 0.04fF $ **FLOATING
C1099 VDD.n942 0 0.04fF $ **FLOATING
C1100 VDD.t184 0 0.01fF
C1101 VDD.n943 0 0.02fF $ **FLOATING
C1102 VDD.n944 0 0.03fF $ **FLOATING
C1103 VDD.n945 0 0.02fF $ **FLOATING
C1104 VDD.n946 0 0.03fF $ **FLOATING
C1105 VDD.n947 0 0.04fF $ **FLOATING
C1106 VDD.n948 0 0.02fF $ **FLOATING
C1107 VDD.n949 0 0.03fF $ **FLOATING
C1108 VDD.n950 0 0.04fF $ **FLOATING
C1109 VDD.t210 0 0.01fF
C1110 VDD.t78 0 0.01fF
C1111 VDD.n951 0 0.03fF $ **FLOATING
C1112 VDD.n952 0 0.03fF $ **FLOATING
C1113 VDD.n953 0 0.02fF $ **FLOATING
C1114 VDD.n954 0 0.02fF $ **FLOATING
C1115 VDD.n955 0 0.04fF $ **FLOATING
C1116 VDD.n956 0 0.02fF $ **FLOATING
C1117 VDD.n957 0 0.03fF $ **FLOATING
C1118 VDD.n958 0 0.04fF $ **FLOATING
C1119 VDD.n959 0 0.02fF $ **FLOATING
C1120 VDD.n960 0 0.03fF $ **FLOATING
C1121 VDD.n961 0 0.04fF $ **FLOATING
C1122 VDD.n962 0 0.02fF $ **FLOATING
C1123 VDD.n963 0 0.03fF $ **FLOATING
C1124 VDD.n964 0 0.04fF $ **FLOATING
C1125 VDD.t178 0 0.03fF
C1126 VDD.n965 0 0.06fF $ **FLOATING
C1127 VDD.n966 0 0.02fF $ **FLOATING
C1128 VDD.n967 0 0.02fF $ **FLOATING
C1129 VDD.n968 0 0.04fF $ **FLOATING
C1130 VDD.n969 0 0.02fF $ **FLOATING
C1131 VDD.n970 0 0.03fF $ **FLOATING
C1132 VDD.n971 0 0.04fF $ **FLOATING
C1133 VDD.t209 0 0.01fF
C1134 VDD.t44 0 0.01fF
C1135 VDD.n972 0 0.02fF $ **FLOATING
C1136 VDD.n973 0 0.03fF $ **FLOATING
C1137 VDD.n974 0 0.02fF $ **FLOATING
C1138 VDD.n975 0 0.02fF $ **FLOATING
C1139 VDD.n976 0 0.04fF $ **FLOATING
C1140 VDD.n977 0 0.02fF $ **FLOATING
C1141 VDD.n978 0 0.03fF $ **FLOATING
C1142 VDD.n979 0 0.04fF $ **FLOATING
C1143 VDD.n980 0 0.02fF $ **FLOATING
C1144 VDD.n981 0 0.03fF $ **FLOATING
C1145 VDD.n982 0 0.04fF $ **FLOATING
C1146 VDD.n983 0 0.02fF $ **FLOATING
C1147 VDD.n984 0 0.03fF $ **FLOATING
C1148 VDD.n985 0 0.04fF $ **FLOATING
C1149 VDD.n986 0 0.02fF $ **FLOATING
C1150 VDD.n987 0 0.03fF $ **FLOATING
C1151 VDD.n988 0 0.04fF $ **FLOATING
C1152 VDD.t102 0 0.01fF
C1153 VDD.n989 0 0.05fF $ **FLOATING
C1154 VDD.n990 0 0.02fF $ **FLOATING
C1155 VDD.n991 0 0.02fF $ **FLOATING
C1156 VDD.n992 0 0.04fF $ **FLOATING
C1157 VDD.n993 0 0.02fF $ **FLOATING
C1158 VDD.n994 0 0.03fF $ **FLOATING
C1159 VDD.n995 0 0.04fF $ **FLOATING
C1160 VDD.n996 0 0.02fF $ **FLOATING
C1161 VDD.n997 0 0.03fF $ **FLOATING
C1162 VDD.n998 0 0.04fF $ **FLOATING
C1163 VDD.t182 0 0.01fF
C1164 VDD.t231 0 0.01fF
C1165 VDD.n999 0 0.03fF $ **FLOATING
C1166 VDD.n1000 0 0.04fF $ **FLOATING
C1167 VDD.n1001 0 0.02fF $ **FLOATING
C1168 VDD.n1002 0 0.02fF $ **FLOATING
C1169 VDD.n1003 0 0.04fF $ **FLOATING
C1170 VDD.n1004 0 0.02fF $ **FLOATING
C1171 VDD.n1005 0 0.03fF $ **FLOATING
C1172 VDD.n1006 0 0.04fF $ **FLOATING
C1173 VDD.n1007 0 0.02fF $ **FLOATING
C1174 VDD.n1008 0 0.03fF $ **FLOATING
C1175 VDD.n1009 0 0.04fF $ **FLOATING
C1176 VDD.t13 0 0.01fF
C1177 VDD.t68 0 0.01fF
C1178 VDD.n1010 0 0.07fF $ **FLOATING
C1179 VDD.n1011 0 0.03fF $ **FLOATING
C1180 VDD.n1012 0 0.02fF $ **FLOATING
C1181 VDD.n1013 0 0.02fF $ **FLOATING
C1182 VDD.n1014 0 0.04fF $ **FLOATING
C1183 VDD.n1015 0 0.02fF $ **FLOATING
C1184 VDD.n1016 0 0.03fF $ **FLOATING
C1185 VDD.n1017 0 0.04fF $ **FLOATING
C1186 VDD.n1018 0 0.02fF $ **FLOATING
C1187 VDD.n1019 0 0.03fF $ **FLOATING
C1188 VDD.n1020 0 0.04fF $ **FLOATING
C1189 VDD.n1021 0 0.02fF $ **FLOATING
C1190 VDD.n1022 0 0.03fF $ **FLOATING
C1191 VDD.n1023 0 0.04fF $ **FLOATING
C1192 VDD.t22 0 0.02fF
C1193 VDD.n1024 0 0.04fF $ **FLOATING
C1194 VDD.n1025 0 0.04fF $ **FLOATING
C1195 VDD.t113 0 0.01fF
C1196 VDD.n1026 0 0.02fF $ **FLOATING
C1197 VDD.n1027 0 0.03fF $ **FLOATING
C1198 VDD.n1028 0 0.02fF $ **FLOATING
C1199 VDD.n1029 0 0.03fF $ **FLOATING
C1200 VDD.n1030 0 0.04fF $ **FLOATING
C1201 VDD.n1031 0 0.02fF $ **FLOATING
C1202 VDD.n1032 0 0.03fF $ **FLOATING
C1203 VDD.n1033 0 0.04fF $ **FLOATING
C1204 VDD.t212 0 0.01fF
C1205 VDD.t236 0 0.01fF
C1206 VDD.n1034 0 0.03fF $ **FLOATING
C1207 VDD.n1035 0 0.03fF $ **FLOATING
C1208 VDD.n1036 0 0.02fF $ **FLOATING
C1209 VDD.n1037 0 0.02fF $ **FLOATING
C1210 VDD.n1038 0 0.04fF $ **FLOATING
C1211 VDD.n1039 0 0.02fF $ **FLOATING
C1212 VDD.n1040 0 0.03fF $ **FLOATING
C1213 VDD.n1041 0 0.04fF $ **FLOATING
C1214 VDD.n1042 0 0.02fF $ **FLOATING
C1215 VDD.n1043 0 0.03fF $ **FLOATING
C1216 VDD.n1044 0 0.04fF $ **FLOATING
C1217 VDD.n1045 0 0.02fF $ **FLOATING
C1218 VDD.n1046 0 0.03fF $ **FLOATING
C1219 VDD.n1047 0 0.04fF $ **FLOATING
C1220 VDD.t100 0 0.03fF
C1221 VDD.n1048 0 0.06fF $ **FLOATING
C1222 VDD.n1049 0 0.02fF $ **FLOATING
C1223 VDD.n1050 0 0.02fF $ **FLOATING
C1224 VDD.n1051 0 0.04fF $ **FLOATING
C1225 VDD.n1052 0 0.02fF $ **FLOATING
C1226 VDD.n1053 0 0.03fF $ **FLOATING
C1227 VDD.n1054 0 0.04fF $ **FLOATING
C1228 VDD.t211 0 0.01fF
C1229 VDD.t85 0 0.01fF
C1230 VDD.n1055 0 0.02fF $ **FLOATING
C1231 VDD.n1056 0 0.03fF $ **FLOATING
C1232 VDD.n1057 0 0.02fF $ **FLOATING
C1233 VDD.n1058 0 0.02fF $ **FLOATING
C1234 VDD.n1059 0 0.04fF $ **FLOATING
C1235 VDD.n1060 0 0.02fF $ **FLOATING
C1236 VDD.n1061 0 0.03fF $ **FLOATING
C1237 VDD.n1062 0 0.04fF $ **FLOATING
C1238 VDD.n1063 0 0.02fF $ **FLOATING
C1239 VDD.n1064 0 0.03fF $ **FLOATING
C1240 VDD.n1065 0 0.04fF $ **FLOATING
C1241 VDD.n1066 0 0.02fF $ **FLOATING
C1242 VDD.n1067 0 0.03fF $ **FLOATING
C1243 VDD.n1068 0 0.04fF $ **FLOATING
C1244 VDD.n1069 0 0.02fF $ **FLOATING
C1245 VDD.n1070 0 0.03fF $ **FLOATING
C1246 VDD.n1071 0 0.04fF $ **FLOATING
C1247 VDD.t159 0 0.01fF
C1248 VDD.n1072 0 0.05fF $ **FLOATING
C1249 VDD.n1073 0 0.02fF $ **FLOATING
C1250 VDD.n1074 0 0.02fF $ **FLOATING
C1251 VDD.n1075 0 0.04fF $ **FLOATING
C1252 VDD.n1076 0 0.02fF $ **FLOATING
C1253 VDD.n1077 0 0.03fF $ **FLOATING
C1254 VDD.n1078 0 0.04fF $ **FLOATING
C1255 VDD.n1079 0 0.02fF $ **FLOATING
C1256 VDD.n1080 0 0.03fF $ **FLOATING
C1257 VDD.n1081 0 0.04fF $ **FLOATING
C1258 VDD.t104 0 0.01fF
C1259 VDD.t54 0 0.01fF
C1260 VDD.n1082 0 0.03fF $ **FLOATING
C1261 VDD.n1083 0 0.04fF $ **FLOATING
C1262 VDD.n1084 0 0.02fF $ **FLOATING
C1263 VDD.n1085 0 0.02fF $ **FLOATING
C1264 VDD.n1086 0 0.04fF $ **FLOATING
C1265 VDD.n1087 0 0.02fF $ **FLOATING
C1266 VDD.n1088 0 0.03fF $ **FLOATING
C1267 VDD.n1089 0 0.04fF $ **FLOATING
C1268 VDD.n1090 0 0.02fF $ **FLOATING
C1269 VDD.n1091 0 0.03fF $ **FLOATING
C1270 VDD.n1092 0 0.04fF $ **FLOATING
C1271 VDD.t14 0 0.01fF
C1272 VDD.t160 0 0.01fF
C1273 VDD.n1093 0 0.07fF $ **FLOATING
C1274 VDD.n1094 0 0.03fF $ **FLOATING
C1275 VDD.n1095 0 0.02fF $ **FLOATING
C1276 VDD.n1096 0 0.02fF $ **FLOATING
C1277 VDD.n1097 0 0.04fF $ **FLOATING
C1278 VDD.n1098 0 0.02fF $ **FLOATING
C1279 VDD.n1099 0 0.03fF $ **FLOATING
C1280 VDD.n1100 0 0.04fF $ **FLOATING
C1281 VDD.n1101 0 0.02fF $ **FLOATING
C1282 VDD.n1102 0 0.03fF $ **FLOATING
C1283 VDD.n1103 0 0.04fF $ **FLOATING
C1284 VDD.n1104 0 0.02fF $ **FLOATING
C1285 VDD.n1105 0 0.03fF $ **FLOATING
C1286 VDD.n1106 0 0.04fF $ **FLOATING
C1287 VDD.t157 0 0.02fF
C1288 VDD.n1107 0 0.04fF $ **FLOATING
C1289 VDD.n1108 0 0.04fF $ **FLOATING
C1290 VDD.t103 0 0.01fF
C1291 VDD.n1109 0 0.02fF $ **FLOATING
C1292 VDD.n1110 0 0.03fF $ **FLOATING
C1293 VDD.n1111 0 0.02fF $ **FLOATING
C1294 VDD.n1112 0 0.03fF $ **FLOATING
C1295 VDD.n1113 0 0.04fF $ **FLOATING
C1296 VDD.n1114 0 0.02fF $ **FLOATING
C1297 VDD.n1115 0 0.03fF $ **FLOATING
C1298 VDD.n1116 0 0.04fF $ **FLOATING
C1299 VDD.t214 0 0.01fF
C1300 VDD.t139 0 0.01fF
C1301 VDD.n1117 0 0.03fF $ **FLOATING
C1302 VDD.n1118 0 0.03fF $ **FLOATING
C1303 VDD.n1119 0 0.02fF $ **FLOATING
C1304 VDD.n1120 0 0.02fF $ **FLOATING
C1305 VDD.n1121 0 0.04fF $ **FLOATING
C1306 VDD.n1122 0 0.02fF $ **FLOATING
C1307 VDD.n1123 0 0.03fF $ **FLOATING
C1308 VDD.n1124 0 0.04fF $ **FLOATING
C1309 VDD.n1125 0 0.02fF $ **FLOATING
C1310 VDD.n1126 0 0.03fF $ **FLOATING
C1311 VDD.n1127 0 0.04fF $ **FLOATING
C1312 VDD.n1128 0 0.02fF $ **FLOATING
C1313 VDD.n1129 0 0.03fF $ **FLOATING
C1314 VDD.n1130 0 0.04fF $ **FLOATING
C1315 VDD.t65 0 0.03fF
C1316 VDD.n1131 0 0.06fF $ **FLOATING
C1317 VDD.n1132 0 0.02fF $ **FLOATING
C1318 VDD.n1133 0 0.02fF $ **FLOATING
C1319 VDD.n1134 0 0.04fF $ **FLOATING
C1320 VDD.n1135 0 0.02fF $ **FLOATING
C1321 VDD.n1136 0 0.03fF $ **FLOATING
C1322 VDD.n1137 0 0.04fF $ **FLOATING
C1323 VDD.t213 0 0.01fF
C1324 VDD.t156 0 0.01fF
C1325 VDD.n1138 0 0.02fF $ **FLOATING
C1326 VDD.n1139 0 0.03fF $ **FLOATING
C1327 VDD.n1140 0 0.02fF $ **FLOATING
C1328 VDD.n1141 0 0.02fF $ **FLOATING
C1329 VDD.n1142 0 0.04fF $ **FLOATING
C1330 VDD.n1143 0 0.02fF $ **FLOATING
C1331 VDD.n1144 0 0.03fF $ **FLOATING
C1332 VDD.n1145 0 0.04fF $ **FLOATING
C1333 VDD.n1146 0 0.02fF $ **FLOATING
C1334 VDD.n1147 0 0.03fF $ **FLOATING
C1335 VDD.n1148 0 0.04fF $ **FLOATING
C1336 VDD.n1149 0 0.02fF $ **FLOATING
C1337 VDD.n1150 0 0.03fF $ **FLOATING
C1338 VDD.n1151 0 0.04fF $ **FLOATING
C1339 VDD.n1152 0 0.02fF $ **FLOATING
C1340 VDD.n1153 0 0.03fF $ **FLOATING
C1341 VDD.n1154 0 0.04fF $ **FLOATING
C1342 VDD.n1155 0 0.04fF $ **FLOATING
C1343 VDD.n1156 0 0.04fF $ **FLOATING
C1344 VDD.n1157 0 0.04fF $ **FLOATING
C1345 VDD.n1158 0 0.04fF $ **FLOATING
C1346 VDD.n1159 0 0.04fF $ **FLOATING
C1347 VDD.n1160 0 0.04fF $ **FLOATING
C1348 VDD.n1161 0 0.05fF $ **FLOATING
C1349 VDD.t37 0 0.01fF
C1350 VDD.t123 0 0.01fF
C1351 VDD.n1162 0 0.03fF $ **FLOATING
C1352 VDD.n1163 0 0.04fF $ **FLOATING
C1353 VDD.n1164 0 0.02fF $ **FLOATING
C1354 VDD.n1165 0 0.02fF $ **FLOATING
C1355 VDD.n1166 0 0.09fF $ **FLOATING
C1356 VDD.n1167 0 0.02fF $ **FLOATING
C1357 VDD.n1168 0 0.03fF $ **FLOATING
C1358 VDD.n1169 0 0.04fF $ **FLOATING
C1359 VDD.n1170 0 0.02fF $ **FLOATING
C1360 VDD.n1171 0 0.03fF $ **FLOATING
C1361 VDD.n1172 0 0.04fF $ **FLOATING
C1362 VDD.t25 0 0.01fF
C1363 VDD.n1173 0 0.05fF $ **FLOATING
C1364 VDD.n1174 0 0.02fF $ **FLOATING
C1365 VDD.n1175 0 0.02fF $ **FLOATING
C1366 VDD.n1176 0 0.04fF $ **FLOATING
C1367 VDD.n1177 0 0.02fF $ **FLOATING
C1368 VDD.n1178 0 0.03fF $ **FLOATING
C1369 VDD.n1179 0 0.04fF $ **FLOATING
C1370 VDD.n1180 0 0.02fF $ **FLOATING
C1371 VDD.n1181 0 0.03fF $ **FLOATING
C1372 VDD.n1182 0 0.04fF $ **FLOATING
C1373 VDD.n1183 0 0.02fF $ **FLOATING
C1374 VDD.n1184 0 0.03fF $ **FLOATING
C1375 VDD.n1185 0 0.04fF $ **FLOATING
C1376 VDD.n1186 0 0.02fF $ **FLOATING
C1377 VDD.n1187 0 0.03fF $ **FLOATING
C1378 VDD.n1188 0 0.04fF $ **FLOATING
C1379 VDD.t225 0 0.01fF
C1380 VDD.t70 0 0.01fF
C1381 VDD.n1189 0 0.02fF $ **FLOATING
C1382 VDD.n1190 0 0.03fF $ **FLOATING
C1383 VDD.n1191 0 0.02fF $ **FLOATING
C1384 VDD.n1192 0 0.02fF $ **FLOATING
C1385 VDD.n1193 0 0.04fF $ **FLOATING
C1386 VDD.n1194 0 0.02fF $ **FLOATING
C1387 VDD.n1195 0 0.03fF $ **FLOATING
C1388 VDD.n1196 0 0.04fF $ **FLOATING
C1389 VDD.t33 0 0.03fF
C1390 VDD.n1197 0 0.06fF $ **FLOATING
C1391 VDD.n1198 0 0.02fF $ **FLOATING
C1392 VDD.n1199 0 0.02fF $ **FLOATING
C1393 VDD.n1200 0 0.04fF $ **FLOATING
C1394 VDD.n1201 0 0.02fF $ **FLOATING
C1395 VDD.n1202 0 0.03fF $ **FLOATING
C1396 VDD.n1203 0 0.04fF $ **FLOATING
C1397 VDD.n1204 0 0.02fF $ **FLOATING
C1398 VDD.n1205 0 0.03fF $ **FLOATING
C1399 VDD.n1206 0 0.04fF $ **FLOATING
C1400 VDD.n1207 0 0.02fF $ **FLOATING
C1401 VDD.n1208 0 0.03fF $ **FLOATING
C1402 VDD.n1209 0 0.04fF $ **FLOATING
C1403 VDD.t226 0 0.01fF
C1404 VDD.t132 0 0.01fF
C1405 VDD.n1210 0 0.03fF $ **FLOATING
C1406 VDD.n1211 0 0.03fF $ **FLOATING
C1407 VDD.n1212 0 0.02fF $ **FLOATING
C1408 VDD.n1213 0 0.02fF $ **FLOATING
C1409 VDD.n1214 0 0.04fF $ **FLOATING
C1410 VDD.n1215 0 0.02fF $ **FLOATING
C1411 VDD.n1216 0 0.03fF $ **FLOATING
C1412 VDD.n1217 0 0.04fF $ **FLOATING
C1413 VDD.t131 0 0.02fF
C1414 VDD.n1218 0 0.04fF $ **FLOATING
C1415 VDD.n1219 0 0.04fF $ **FLOATING
C1416 VDD.t83 0 0.01fF
C1417 VDD.n1220 0 0.02fF $ **FLOATING
C1418 VDD.n1221 0 0.03fF $ **FLOATING
C1419 VDD.n1222 0 0.02fF $ **FLOATING
C1420 VDD.n1223 0 0.03fF $ **FLOATING
C1421 VDD.n1224 0 0.04fF $ **FLOATING
C1422 VDD.n1225 0 0.02fF $ **FLOATING
C1423 VDD.n1226 0 0.03fF $ **FLOATING
C1424 VDD.n1227 0 0.04fF $ **FLOATING
C1425 VDD.n1228 0 0.02fF $ **FLOATING
C1426 VDD.n1229 0 0.03fF $ **FLOATING
C1427 VDD.n1230 0 0.04fF $ **FLOATING
C1428 VDD.n1231 0 0.02fF $ **FLOATING
C1429 VDD.n1232 0 0.03fF $ **FLOATING
C1430 VDD.n1233 0 0.04fF $ **FLOATING
C1431 VDD.t133 0 0.01fF
C1432 VDD.t165 0 0.01fF
C1433 VDD.n1234 0 0.07fF $ **FLOATING
C1434 VDD.n1235 0 0.03fF $ **FLOATING
C1435 VDD.n1236 0 0.02fF $ **FLOATING
C1436 VDD.n1237 0 0.02fF $ **FLOATING
C1437 VDD.n1238 0 0.04fF $ **FLOATING
C1438 VDD.n1239 0 0.02fF $ **FLOATING
C1439 VDD.n1240 0 0.03fF $ **FLOATING
C1440 VDD.n1241 0 0.04fF $ **FLOATING
C1441 VDD.n1242 0 0.02fF $ **FLOATING
C1442 VDD.n1243 0 0.03fF $ **FLOATING
C1443 VDD.n1244 0 0.04fF $ **FLOATING
C1444 VDD.t42 0 0.01fF
C1445 VDD.t57 0 0.01fF
C1446 VDD.n1245 0 0.03fF $ **FLOATING
C1447 VDD.n1246 0 0.04fF $ **FLOATING
C1448 VDD.n1247 0 0.02fF $ **FLOATING
C1449 VDD.n1248 0 0.02fF $ **FLOATING
C1450 VDD.n1249 0 0.04fF $ **FLOATING
C1451 VDD.n1250 0 0.02fF $ **FLOATING
C1452 VDD.n1251 0 0.03fF $ **FLOATING
C1453 VDD.n1252 0 0.04fF $ **FLOATING
C1454 VDD.n1253 0 0.02fF $ **FLOATING
C1455 VDD.n1254 0 0.03fF $ **FLOATING
C1456 VDD.n1255 0 0.04fF $ **FLOATING
C1457 VDD.t59 0 0.01fF
C1458 VDD.n1256 0 0.05fF $ **FLOATING
C1459 VDD.n1257 0 0.02fF $ **FLOATING
C1460 VDD.n1258 0 0.02fF $ **FLOATING
C1461 VDD.n1259 0 0.04fF $ **FLOATING
C1462 VDD.n1260 0 0.02fF $ **FLOATING
C1463 VDD.n1261 0 0.03fF $ **FLOATING
C1464 VDD.n1262 0 0.04fF $ **FLOATING
C1465 VDD.n1263 0 0.02fF $ **FLOATING
C1466 VDD.n1264 0 0.03fF $ **FLOATING
C1467 VDD.n1265 0 0.04fF $ **FLOATING
C1468 VDD.n1266 0 0.02fF $ **FLOATING
C1469 VDD.n1267 0 0.03fF $ **FLOATING
C1470 VDD.n1268 0 0.04fF $ **FLOATING
C1471 VDD.n1269 0 0.02fF $ **FLOATING
C1472 VDD.n1270 0 0.03fF $ **FLOATING
C1473 VDD.n1271 0 0.04fF $ **FLOATING
C1474 VDD.t223 0 0.01fF
C1475 VDD.t30 0 0.01fF
C1476 VDD.n1272 0 0.02fF $ **FLOATING
C1477 VDD.n1273 0 0.03fF $ **FLOATING
C1478 VDD.n1274 0 0.02fF $ **FLOATING
C1479 VDD.n1275 0 0.02fF $ **FLOATING
C1480 VDD.n1276 0 0.04fF $ **FLOATING
C1481 VDD.n1277 0 0.02fF $ **FLOATING
C1482 VDD.n1278 0 0.03fF $ **FLOATING
C1483 VDD.n1279 0 0.04fF $ **FLOATING
C1484 VDD.t63 0 0.03fF
C1485 VDD.n1280 0 0.06fF $ **FLOATING
C1486 VDD.n1281 0 0.02fF $ **FLOATING
C1487 VDD.n1282 0 0.02fF $ **FLOATING
C1488 VDD.n1283 0 0.04fF $ **FLOATING
C1489 VDD.n1284 0 0.02fF $ **FLOATING
C1490 VDD.n1285 0 0.03fF $ **FLOATING
C1491 VDD.n1286 0 0.04fF $ **FLOATING
C1492 VDD.n1287 0 0.02fF $ **FLOATING
C1493 VDD.n1288 0 0.03fF $ **FLOATING
C1494 VDD.n1289 0 0.04fF $ **FLOATING
C1495 VDD.n1290 0 0.02fF $ **FLOATING
C1496 VDD.n1291 0 0.03fF $ **FLOATING
C1497 VDD.n1292 0 0.04fF $ **FLOATING
C1498 VDD.t224 0 0.01fF
C1499 VDD.t34 0 0.01fF
C1500 VDD.n1293 0 0.03fF $ **FLOATING
C1501 VDD.n1294 0 0.03fF $ **FLOATING
C1502 VDD.n1295 0 0.02fF $ **FLOATING
C1503 VDD.n1296 0 0.02fF $ **FLOATING
C1504 VDD.n1297 0 0.04fF $ **FLOATING
C1505 VDD.n1298 0 0.02fF $ **FLOATING
C1506 VDD.n1299 0 0.03fF $ **FLOATING
C1507 VDD.n1300 0 0.04fF $ **FLOATING
C1508 VDD.t158 0 0.02fF
C1509 VDD.n1301 0 0.04fF $ **FLOATING
C1510 VDD.n1302 0 0.04fF $ **FLOATING
C1511 VDD.t74 0 0.01fF
C1512 VDD.n1303 0 0.02fF $ **FLOATING
C1513 VDD.n1304 0 0.03fF $ **FLOATING
C1514 VDD.n1305 0 0.02fF $ **FLOATING
C1515 VDD.n1306 0 0.03fF $ **FLOATING
C1516 VDD.n1307 0 0.04fF $ **FLOATING
C1517 VDD.n1308 0 0.02fF $ **FLOATING
C1518 VDD.n1309 0 0.03fF $ **FLOATING
C1519 VDD.n1310 0 0.04fF $ **FLOATING
C1520 VDD.n1311 0 0.02fF $ **FLOATING
C1521 VDD.n1312 0 0.03fF $ **FLOATING
C1522 VDD.n1313 0 0.04fF $ **FLOATING
C1523 VDD.n1314 0 0.02fF $ **FLOATING
C1524 VDD.n1315 0 0.03fF $ **FLOATING
C1525 VDD.n1316 0 0.04fF $ **FLOATING
C1526 VDD.t60 0 0.01fF
C1527 VDD.t28 0 0.01fF
C1528 VDD.n1317 0 0.07fF $ **FLOATING
C1529 VDD.n1318 0 0.03fF $ **FLOATING
C1530 VDD.n1319 0 0.02fF $ **FLOATING
C1531 VDD.n1320 0 0.02fF $ **FLOATING
C1532 VDD.n1321 0 0.04fF $ **FLOATING
C1533 VDD.n1322 0 0.02fF $ **FLOATING
C1534 VDD.n1323 0 0.03fF $ **FLOATING
C1535 VDD.n1324 0 0.04fF $ **FLOATING
C1536 VDD.n1325 0 0.02fF $ **FLOATING
C1537 VDD.n1326 0 0.03fF $ **FLOATING
C1538 VDD.n1327 0 0.04fF $ **FLOATING
C1539 VDD.t75 0 0.01fF
C1540 VDD.t17 0 0.01fF
C1541 VDD.n1328 0 0.03fF $ **FLOATING
C1542 VDD.n1329 0 0.04fF $ **FLOATING
C1543 VDD.n1330 0 0.02fF $ **FLOATING
C1544 VDD.n1331 0 0.02fF $ **FLOATING
C1545 VDD.n1332 0 0.04fF $ **FLOATING
C1546 VDD.n1333 0 0.02fF $ **FLOATING
C1547 VDD.n1334 0 0.03fF $ **FLOATING
C1548 VDD.n1335 0 0.04fF $ **FLOATING
C1549 VDD.n1336 0 0.02fF $ **FLOATING
C1550 VDD.n1337 0 0.03fF $ **FLOATING
C1551 VDD.n1338 0 0.04fF $ **FLOATING
C1552 VDD.t67 0 0.01fF
C1553 VDD.n1339 0 0.05fF $ **FLOATING
C1554 VDD.n1340 0 0.02fF $ **FLOATING
C1555 VDD.n1341 0 0.02fF $ **FLOATING
C1556 VDD.n1342 0 0.04fF $ **FLOATING
C1557 VDD.n1343 0 0.02fF $ **FLOATING
C1558 VDD.n1344 0 0.03fF $ **FLOATING
C1559 VDD.n1345 0 0.04fF $ **FLOATING
C1560 VDD.n1346 0 0.02fF $ **FLOATING
C1561 VDD.n1347 0 0.03fF $ **FLOATING
C1562 VDD.n1348 0 0.04fF $ **FLOATING
C1563 VDD.n1349 0 0.02fF $ **FLOATING
C1564 VDD.n1350 0 0.03fF $ **FLOATING
C1565 VDD.n1351 0 0.04fF $ **FLOATING
C1566 VDD.n1352 0 0.02fF $ **FLOATING
C1567 VDD.n1353 0 0.03fF $ **FLOATING
C1568 VDD.n1354 0 0.04fF $ **FLOATING
C1569 VDD.t221 0 0.01fF
C1570 VDD.t23 0 0.01fF
C1571 VDD.n1355 0 0.02fF $ **FLOATING
C1572 VDD.n1356 0 0.03fF $ **FLOATING
C1573 VDD.n1357 0 0.02fF $ **FLOATING
C1574 VDD.n1358 0 0.02fF $ **FLOATING
C1575 VDD.n1359 0 0.04fF $ **FLOATING
C1576 VDD.n1360 0 0.02fF $ **FLOATING
C1577 VDD.n1361 0 0.03fF $ **FLOATING
C1578 VDD.n1362 0 0.04fF $ **FLOATING
C1579 VDD.t86 0 0.03fF
C1580 VDD.n1363 0 0.06fF $ **FLOATING
C1581 VDD.n1364 0 0.02fF $ **FLOATING
C1582 VDD.n1365 0 0.02fF $ **FLOATING
C1583 VDD.n1366 0 0.04fF $ **FLOATING
C1584 VDD.n1367 0 0.02fF $ **FLOATING
C1585 VDD.n1368 0 0.03fF $ **FLOATING
C1586 VDD.n1369 0 0.04fF $ **FLOATING
C1587 VDD.n1370 0 0.02fF $ **FLOATING
C1588 VDD.n1371 0 0.03fF $ **FLOATING
C1589 VDD.n1372 0 0.04fF $ **FLOATING
C1590 VDD.n1373 0 0.02fF $ **FLOATING
C1591 VDD.n1374 0 0.03fF $ **FLOATING
C1592 VDD.n1375 0 0.04fF $ **FLOATING
C1593 VDD.t222 0 0.01fF
C1594 VDD.t234 0 0.01fF
C1595 VDD.n1376 0 0.03fF $ **FLOATING
C1596 VDD.n1377 0 0.03fF $ **FLOATING
C1597 VDD.n1378 0 0.02fF $ **FLOATING
C1598 VDD.n1379 0 0.02fF $ **FLOATING
C1599 VDD.n1380 0 0.04fF $ **FLOATING
C1600 VDD.n1381 0 0.02fF $ **FLOATING
C1601 VDD.n1382 0 0.03fF $ **FLOATING
C1602 VDD.n1383 0 0.04fF $ **FLOATING
C1603 VDD.t27 0 0.02fF
C1604 VDD.n1384 0 0.04fF $ **FLOATING
C1605 VDD.n1385 0 0.04fF $ **FLOATING
C1606 VDD.t82 0 0.01fF
C1607 VDD.n1386 0 0.02fF $ **FLOATING
C1608 VDD.n1387 0 0.03fF $ **FLOATING
C1609 VDD.n1388 0 0.02fF $ **FLOATING
C1610 VDD.n1389 0 0.03fF $ **FLOATING
C1611 VDD.n1390 0 0.04fF $ **FLOATING
C1612 VDD.n1391 0 0.02fF $ **FLOATING
C1613 VDD.n1392 0 0.03fF $ **FLOATING
C1614 VDD.n1393 0 0.04fF $ **FLOATING
C1615 VDD.n1394 0 0.02fF $ **FLOATING
C1616 VDD.n1395 0 0.03fF $ **FLOATING
C1617 VDD.n1396 0 0.04fF $ **FLOATING
C1618 VDD.n1397 0 0.02fF $ **FLOATING
C1619 VDD.n1398 0 0.03fF $ **FLOATING
C1620 VDD.n1399 0 0.04fF $ **FLOATING
C1621 VDD.t62 0 0.01fF
C1622 VDD.t24 0 0.01fF
C1623 VDD.n1400 0 0.07fF $ **FLOATING
C1624 VDD.n1401 0 0.03fF $ **FLOATING
C1625 VDD.n1402 0 0.02fF $ **FLOATING
C1626 VDD.n1403 0 0.02fF $ **FLOATING
C1627 VDD.n1404 0 0.04fF $ **FLOATING
C1628 VDD.n1405 0 0.02fF $ **FLOATING
C1629 VDD.n1406 0 0.03fF $ **FLOATING
C1630 VDD.n1407 0 0.04fF $ **FLOATING
C1631 VDD.n1408 0 0.02fF $ **FLOATING
C1632 VDD.n1409 0 0.03fF $ **FLOATING
C1633 VDD.n1410 0 0.04fF $ **FLOATING
C1634 VDD.t29 0 0.01fF
C1635 VDD.t21 0 0.01fF
C1636 VDD.n1411 0 0.03fF $ **FLOATING
C1637 VDD.n1412 0 0.04fF $ **FLOATING
C1638 VDD.n1413 0 0.02fF $ **FLOATING
C1639 VDD.n1414 0 0.02fF $ **FLOATING
C1640 VDD.n1415 0 0.04fF $ **FLOATING
C1641 VDD.n1416 0 0.02fF $ **FLOATING
C1642 VDD.n1417 0 0.03fF $ **FLOATING
C1643 VDD.n1418 0 0.04fF $ **FLOATING
C1644 VDD.n1419 0 0.02fF $ **FLOATING
C1645 VDD.n1420 0 0.03fF $ **FLOATING
C1646 VDD.n1421 0 0.04fF $ **FLOATING
C1647 VDD.t98 0 0.01fF
C1648 VDD.n1422 0 0.05fF $ **FLOATING
C1649 VDD.n1423 0 0.02fF $ **FLOATING
C1650 VDD.n1424 0 0.02fF $ **FLOATING
C1651 VDD.n1425 0 0.04fF $ **FLOATING
C1652 VDD.n1426 0 0.02fF $ **FLOATING
C1653 VDD.n1427 0 0.03fF $ **FLOATING
C1654 VDD.n1428 0 0.04fF $ **FLOATING
C1655 VDD.n1429 0 0.02fF $ **FLOATING
C1656 VDD.n1430 0 0.03fF $ **FLOATING
C1657 VDD.n1431 0 0.04fF $ **FLOATING
C1658 VDD.n1432 0 0.02fF $ **FLOATING
C1659 VDD.n1433 0 0.03fF $ **FLOATING
C1660 VDD.n1434 0 0.04fF $ **FLOATING
C1661 VDD.n1435 0 0.02fF $ **FLOATING
C1662 VDD.n1436 0 0.03fF $ **FLOATING
C1663 VDD.n1437 0 0.04fF $ **FLOATING
C1664 VDD.t219 0 0.01fF
C1665 VDD.t20 0 0.01fF
C1666 VDD.n1438 0 0.02fF $ **FLOATING
C1667 VDD.n1439 0 0.03fF $ **FLOATING
C1668 VDD.n1440 0 0.02fF $ **FLOATING
C1669 VDD.n1441 0 0.02fF $ **FLOATING
C1670 VDD.n1442 0 0.04fF $ **FLOATING
C1671 VDD.n1443 0 0.02fF $ **FLOATING
C1672 VDD.n1444 0 0.03fF $ **FLOATING
C1673 VDD.n1445 0 0.04fF $ **FLOATING
C1674 VDD.t52 0 0.03fF
C1675 VDD.n1446 0 0.06fF $ **FLOATING
C1676 VDD.n1447 0 0.02fF $ **FLOATING
C1677 VDD.n1448 0 0.02fF $ **FLOATING
C1678 VDD.n1449 0 0.04fF $ **FLOATING
C1679 VDD.n1450 0 0.02fF $ **FLOATING
C1680 VDD.n1451 0 0.03fF $ **FLOATING
C1681 VDD.n1452 0 0.04fF $ **FLOATING
C1682 VDD.n1453 0 0.02fF $ **FLOATING
C1683 VDD.n1454 0 0.03fF $ **FLOATING
C1684 VDD.n1455 0 0.04fF $ **FLOATING
C1685 VDD.n1456 0 0.02fF $ **FLOATING
C1686 VDD.n1457 0 0.03fF $ **FLOATING
C1687 VDD.n1458 0 0.04fF $ **FLOATING
C1688 VDD.t220 0 0.01fF
C1689 VDD.t80 0 0.01fF
C1690 VDD.n1459 0 0.03fF $ **FLOATING
C1691 VDD.n1460 0 0.03fF $ **FLOATING
C1692 VDD.n1461 0 0.02fF $ **FLOATING
C1693 VDD.n1462 0 0.02fF $ **FLOATING
C1694 VDD.n1463 0 0.04fF $ **FLOATING
C1695 VDD.n1464 0 0.02fF $ **FLOATING
C1696 VDD.n1465 0 0.03fF $ **FLOATING
C1697 VDD.n1466 0 0.04fF $ **FLOATING
C1698 VDD.t19 0 0.02fF
C1699 VDD.n1467 0 0.04fF $ **FLOATING
C1700 VDD.n1468 0 0.04fF $ **FLOATING
C1701 VDD.t41 0 0.01fF
C1702 VDD.n1469 0 0.02fF $ **FLOATING
C1703 VDD.n1470 0 0.03fF $ **FLOATING
C1704 VDD.n1471 0 0.02fF $ **FLOATING
C1705 VDD.n1472 0 0.03fF $ **FLOATING
C1706 VDD.n1473 0 0.04fF $ **FLOATING
C1707 VDD.n1474 0 0.02fF $ **FLOATING
C1708 VDD.n1475 0 0.03fF $ **FLOATING
C1709 VDD.n1476 0 0.04fF $ **FLOATING
C1710 VDD.n1477 0 0.02fF $ **FLOATING
C1711 VDD.n1478 0 0.03fF $ **FLOATING
C1712 VDD.n1479 0 0.04fF $ **FLOATING
C1713 VDD.n1480 0 0.02fF $ **FLOATING
C1714 VDD.n1481 0 0.03fF $ **FLOATING
C1715 VDD.n1482 0 0.04fF $ **FLOATING
C1716 VDD.t64 0 0.01fF
C1717 VDD.n1483 0 0.07fF $ **FLOATING
C1718 VDD.n1484 0 0.03fF $ **FLOATING
C1719 VDD.n1485 0 0.02fF $ **FLOATING
C1720 VDD.n1486 0 0.02fF $ **FLOATING
C1721 VDD.n1487 0 0.04fF $ **FLOATING
C1722 VDD.n1488 0 0.02fF $ **FLOATING
C1723 VDD.n1489 0 0.03fF $ **FLOATING
C1724 VDD.n1490 0 0.04fF $ **FLOATING
C1725 VDD.n1491 0 0.02fF $ **FLOATING
C1726 VDD.n1492 0 0.03fF $ **FLOATING
C1727 VDD.n1493 0 0.04fF $ **FLOATING
C1728 VDD.t144 0 0.01fF
C1729 VDD.t238 0 0.01fF
C1730 VDD.n1494 0 0.03fF $ **FLOATING
C1731 VDD.n1495 0 0.04fF $ **FLOATING
C1732 VDD.n1496 0 0.02fF $ **FLOATING
C1733 VDD.n1497 0 0.02fF $ **FLOATING
C1734 VDD.n1498 0 0.04fF $ **FLOATING
C1735 VDD.n1499 0 0.02fF $ **FLOATING
C1736 VDD.n1500 0 0.03fF $ **FLOATING
C1737 VDD.n1501 0 0.04fF $ **FLOATING
C1738 VDD.n1502 0 0.02fF $ **FLOATING
C1739 VDD.n1503 0 0.03fF $ **FLOATING
C1740 VDD.n1504 0 0.04fF $ **FLOATING
C1741 VDD.t56 0 0.01fF
C1742 VDD.n1505 0 0.05fF $ **FLOATING
C1743 VDD.n1506 0 0.02fF $ **FLOATING
C1744 VDD.n1507 0 0.02fF $ **FLOATING
C1745 VDD.n1508 0 0.04fF $ **FLOATING
C1746 VDD.n1509 0 0.02fF $ **FLOATING
C1747 VDD.n1510 0 0.03fF $ **FLOATING
C1748 VDD.n1511 0 0.04fF $ **FLOATING
C1749 VDD.n1512 0 0.02fF $ **FLOATING
C1750 VDD.n1513 0 0.03fF $ **FLOATING
C1751 VDD.n1514 0 0.04fF $ **FLOATING
C1752 VDD.n1515 0 0.02fF $ **FLOATING
C1753 VDD.n1516 0 0.03fF $ **FLOATING
C1754 VDD.n1517 0 0.04fF $ **FLOATING
C1755 VDD.n1518 0 0.02fF $ **FLOATING
C1756 VDD.n1519 0 0.03fF $ **FLOATING
C1757 VDD.n1520 0 0.04fF $ **FLOATING
C1758 VDD.t217 0 0.01fF
C1759 VDD.t77 0 0.01fF
C1760 VDD.n1521 0 0.02fF $ **FLOATING
C1761 VDD.n1522 0 0.03fF $ **FLOATING
C1762 VDD.n1523 0 0.02fF $ **FLOATING
C1763 VDD.n1524 0 0.02fF $ **FLOATING
C1764 VDD.n1525 0 0.04fF $ **FLOATING
C1765 VDD.n1526 0 0.02fF $ **FLOATING
C1766 VDD.n1527 0 0.03fF $ **FLOATING
C1767 VDD.n1528 0 0.04fF $ **FLOATING
C1768 VDD.n1529 0 0.06fF $ **FLOATING
C1769 VDD.n1530 0 0.02fF $ **FLOATING
C1770 VDD.n1531 0 0.02fF $ **FLOATING
C1771 VDD.n1532 0 0.04fF $ **FLOATING
C1772 VDD.n1533 0 0.02fF $ **FLOATING
C1773 VDD.n1534 0 0.03fF $ **FLOATING
C1774 VDD.n1535 0 0.04fF $ **FLOATING
C1775 VDD.n1536 0 0.02fF $ **FLOATING
C1776 VDD.n1537 0 0.03fF $ **FLOATING
C1777 VDD.n1538 0 0.04fF $ **FLOATING
C1778 VDD.n1539 0 0.02fF $ **FLOATING
C1779 VDD.n1540 0 0.03fF $ **FLOATING
C1780 VDD.n1541 0 0.04fF $ **FLOATING
C1781 VDD.t218 0 0.01fF
C1782 VDD.t38 0 0.01fF
C1783 VDD.n1542 0 0.03fF $ **FLOATING
C1784 VDD.n1543 0 0.03fF $ **FLOATING
C1785 VDD.n1544 0 0.02fF $ **FLOATING
C1786 VDD.n1545 0 0.02fF $ **FLOATING
C1787 VDD.n1546 0 0.04fF $ **FLOATING
C1788 VDD.n1547 0 0.02fF $ **FLOATING
C1789 VDD.n1548 0 0.03fF $ **FLOATING
C1790 VDD.n1549 0 0.04fF $ **FLOATING
C1791 VDD.t232 0 0.02fF
C1792 VDD.n1550 0 0.04fF $ **FLOATING
C1793 VDD.n1551 0 0.04fF $ **FLOATING
C1794 VDD.n1552 0 0.02fF $ **FLOATING
C1795 VDD.n1553 0 0.03fF $ **FLOATING
C1796 VDD.n1554 0 0.02fF $ **FLOATING
C1797 VDD.n1555 0 0.03fF $ **FLOATING
C1798 VDD.n1556 0 0.04fF $ **FLOATING
C1799 VDD.n1557 0 0.02fF $ **FLOATING
C1800 VDD.n1558 0 0.03fF $ **FLOATING
C1801 VDD.n1559 0 0.04fF $ **FLOATING
C1802 VDD.n1560 0 0.02fF $ **FLOATING
C1803 VDD.n1561 0 0.03fF $ **FLOATING
C1804 VDD.n1562 0 0.04fF $ **FLOATING
C1805 VDD.n1563 0 0.02fF $ **FLOATING
C1806 VDD.n1564 0 0.03fF $ **FLOATING
C1807 VDD.n1565 0 0.04fF $ **FLOATING
C1808 VDD.t71 0 0.01fF
C1809 VDD.n1566 0 0.07fF $ **FLOATING
C1810 VDD.n1567 0 0.03fF $ **FLOATING
C1811 VDD.n1568 0 0.02fF $ **FLOATING
C1812 VDD.n1569 0 0.02fF $ **FLOATING
C1813 VDD.n1570 0 0.04fF $ **FLOATING
C1814 VDD.n1571 0 0.02fF $ **FLOATING
C1815 VDD.n1572 0 0.03fF $ **FLOATING
C1816 VDD.n1573 0 0.04fF $ **FLOATING
C1817 VDD.n1574 0 0.02fF $ **FLOATING
C1818 VDD.n1575 0 0.03fF $ **FLOATING
C1819 VDD.n1576 0 0.04fF $ **FLOATING
C1820 VDD.t12 0 0.01fF
C1821 VDD.n1577 0 0.03fF $ **FLOATING
C1822 VDD.n1578 0 0.04fF $ **FLOATING
C1823 VDD.n1579 0 0.02fF $ **FLOATING
C1824 VDD.n1580 0 0.02fF $ **FLOATING
C1825 VDD.n1581 0 0.04fF $ **FLOATING
C1826 VDD.n1582 0 0.02fF $ **FLOATING
C1827 VDD.n1583 0 0.03fF $ **FLOATING
C1828 VDD.n1584 0 0.04fF $ **FLOATING
C1829 VDD.n1585 0 0.02fF $ **FLOATING
C1830 VDD.n1586 0 0.03fF $ **FLOATING
C1831 VDD.n1587 0 0.04fF $ **FLOATING
C1832 VDD.n1588 0 0.05fF $ **FLOATING
C1833 VDD.n1589 0 0.02fF $ **FLOATING
C1834 VDD.n1590 0 0.02fF $ **FLOATING
C1835 VDD.n1591 0 0.04fF $ **FLOATING
C1836 VDD.n1592 0 0.02fF $ **FLOATING
C1837 VDD.n1593 0 0.03fF $ **FLOATING
C1838 VDD.n1594 0 0.04fF $ **FLOATING
C1839 VDD.n1595 0 0.02fF $ **FLOATING
C1840 VDD.n1596 0 0.03fF $ **FLOATING
C1841 VDD.n1597 0 0.04fF $ **FLOATING
C1842 VDD.n1598 0 0.02fF $ **FLOATING
C1843 VDD.n1599 0 0.03fF $ **FLOATING
C1844 VDD.n1600 0 0.04fF $ **FLOATING
C1845 VDD.n1601 0 0.02fF $ **FLOATING
C1846 VDD.n1602 0 0.03fF $ **FLOATING
C1847 VDD.n1603 0 0.04fF $ **FLOATING
C1848 VDD.t215 0 0.01fF
C1849 VDD.t53 0 0.01fF
C1850 VDD.n1604 0 0.02fF $ **FLOATING
C1851 VDD.n1605 0 0.03fF $ **FLOATING
C1852 VDD.n1606 0 0.02fF $ **FLOATING
C1853 VDD.n1607 0 0.02fF $ **FLOATING
C1854 VDD.n1608 0 0.04fF $ **FLOATING
C1855 VDD.n1609 0 0.02fF $ **FLOATING
C1856 VDD.n1610 0 0.03fF $ **FLOATING
C1857 VDD.n1611 0 0.04fF $ **FLOATING
C1858 VDD.t239 0 0.03fF
C1859 VDD.n1612 0 0.06fF $ **FLOATING
C1860 VDD.n1613 0 0.02fF $ **FLOATING
C1861 VDD.n1614 0 0.02fF $ **FLOATING
C1862 VDD.n1615 0 0.04fF $ **FLOATING
C1863 VDD.n1616 0 0.02fF $ **FLOATING
C1864 VDD.n1617 0 0.03fF $ **FLOATING
C1865 VDD.n1618 0 0.04fF $ **FLOATING
C1866 VDD.n1619 0 0.02fF $ **FLOATING
C1867 VDD.n1620 0 0.03fF $ **FLOATING
C1868 VDD.n1621 0 0.04fF $ **FLOATING
C1869 VDD.n1622 0 0.04fF $ **FLOATING
C1870 VDD.n1623 0 0.04fF $ **FLOATING
C1871 VDD.n1624 0 0.04fF $ **FLOATING
C1872 VDD.n1625 0 0.04fF $ **FLOATING
C1873 VDD.n1626 0 0.04fF $ **FLOATING
C1874 VDD.n1627 0 0.04fF $ **FLOATING
C1875 VDD.n1628 0 0.04fF $ **FLOATING
C1876 VDD.n1629 0 0.04fF $ **FLOATING
C1877 VDD.n1630 0 0.02fF $ **FLOATING
C1878 VDD.t175 0 0.01fF
C1879 VDD.n1631 0 0.02fF $ **FLOATING
C1880 VDD.t216 0 0.01fF
C1881 VDD.t26 0 0.01fF
C1882 VDD.n1632 0 0.03fF $ **FLOATING
C1883 VDD.n1633 0 0.02fF $ **FLOATING
C1884 VDD.n1634 0 0.03fF $ **FLOATING
C1885 VDD.n1635 0 0.03fF $ **FLOATING
C1886 VDD.n1636 0 0.02fF $ **FLOATING
C1887 VDD.n1637 0 0.02fF $ **FLOATING
C1888 VDD.n1638 0 0.02fF $ **FLOATING
C1889 VDD.n1639 0 0.03fF $ **FLOATING
C1890 VDD.n1640 0 0.03fF $ **FLOATING
C1891 VDD.n1641 0 0.02fF $ **FLOATING
C1892 VDD.n1642 0 0.03fF $ **FLOATING
C1893 VDD.t47 0 0.02fF
C1894 VDD.n1643 0 0.04fF $ **FLOATING
C1895 VDD.n1644 0 0.04fF $ **FLOATING
C1896 VDD.n1645 0 0.02fF $ **FLOATING
C1897 VDD.n1646 0 0.03fF $ **FLOATING
C1898 VDD.n1647 0 0.02fF $ **FLOATING
C1899 VDD.n1648 0 0.03fF $ **FLOATING
C1900 VDD.n1649 0 0.02fF $ **FLOATING
C1901 VDD.n1650 0 0.03fF $ **FLOATING
C1902 VDD.n1651 0 0.02fF $ **FLOATING
C1903 VDD.n1652 0 0.02fF $ **FLOATING
C1904 VDD.t237 0 0.01fF
C1905 VDD.n1653 0 0.01fF $ **FLOATING
C1906 VDD.n1654 0 0.02fF $ **FLOATING
C1907 VDD.n1655 0 0.02fF $ **FLOATING
C1908 sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0 0.07fF
C1909 sky130_fd_sc_hd__dfrbp_1_0[19]/D 0 0.62fF
C1910 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t8 0 0.01fF $ **FLOATING
C1911 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t5 0 0.01fF $ **FLOATING
C1912 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n0 0 0.03fF $ **FLOATING
C1913 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t0 0 0.01fF $ **FLOATING
C1914 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n1 0 0.01fF $ **FLOATING
C1915 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n2 0 0.03fF $ **FLOATING
C1916 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n3 0 0.01fF $ **FLOATING
C1917 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n4 0 0.03fF $ **FLOATING
C1918 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n5 0 0.01fF $ **FLOATING
C1919 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n6 0 0.03fF $ **FLOATING
C1920 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n7 0 0.01fF $ **FLOATING
C1921 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n8 0 0.02fF $ **FLOATING
C1922 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n9 0 0.04fF $ **FLOATING
C1923 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n10 0 0.01fF $ **FLOATING
C1924 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n11 0 0.03fF $ **FLOATING
C1925 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n12 0 0.01fF $ **FLOATING
C1926 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n13 0 0.03fF $ **FLOATING
C1927 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n14 0 0.01fF $ **FLOATING
C1928 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t4 0 0.01fF $ **FLOATING
C1929 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t1 0 0.00fF $ **FLOATING
C1930 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n15 0 0.06fF $ **FLOATING
C1931 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n16 0 0.01fF $ **FLOATING
C1932 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n17 0 0.03fF $ **FLOATING
C1933 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n18 0 0.02fF $ **FLOATING
C1934 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n19 0 0.06fF $ **FLOATING
C1935 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n20 0 0.12fF $ **FLOATING
C1936 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n21 0 0.01fF $ **FLOATING
C1937 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n22 0 0.03fF $ **FLOATING
C1938 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n23 0 0.04fF $ **FLOATING
C1939 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n24 0 0.01fF $ **FLOATING
C1940 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n25 0 0.02fF $ **FLOATING
C1941 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n26 0 0.04fF $ **FLOATING
C1942 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t2 0 0.01fF $ **FLOATING
C1943 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n27 0 0.03fF $ **FLOATING
C1944 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n28 0 0.03fF $ **FLOATING
C1945 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t6 0 0.01fF $ **FLOATING
C1946 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n29 0 0.02fF $ **FLOATING
C1947 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n30 0 0.03fF $ **FLOATING
C1948 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n31 0 0.01fF $ **FLOATING
C1949 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n32 0 0.02fF $ **FLOATING
C1950 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n33 0 0.04fF $ **FLOATING
C1951 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n34 0 0.01fF $ **FLOATING
C1952 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n35 0 0.02fF $ **FLOATING
C1953 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n36 0 0.04fF $ **FLOATING
C1954 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t7 0 0.00fF $ **FLOATING
C1955 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t3 0 0.01fF $ **FLOATING
C1956 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n37 0 0.02fF $ **FLOATING
C1957 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n38 0 0.02fF $ **FLOATING
C1958 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n39 0 0.01fF $ **FLOATING
C1959 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n40 0 0.02fF $ **FLOATING
C1960 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n41 0 0.04fF $ **FLOATING
C1961 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n42 0 0.01fF $ **FLOATING
C1962 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n43 0 0.03fF $ **FLOATING
C1963 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n44 0 0.04fF $ **FLOATING
C1964 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n45 0 0.01fF $ **FLOATING
C1965 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n46 0 0.03fF $ **FLOATING
C1966 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n47 0 0.04fF $ **FLOATING
C1967 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n48 0 0.01fF $ **FLOATING
C1968 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n49 0 0.03fF $ **FLOATING
C1969 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n50 0 0.04fF $ **FLOATING
C1970 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t9 0 0.03fF $ **FLOATING
C1971 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n51 0 0.05fF $ **FLOATING
C1972 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n52 0 0.01fF $ **FLOATING
C1973 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n53 0 0.02fF $ **FLOATING
C1974 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n54 0 0.04fF $ **FLOATING
C1975 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n55 0 0.01fF $ **FLOATING
C1976 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n56 0 0.02fF $ **FLOATING
C1977 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n57 0 0.04fF $ **FLOATING
C1978 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t11 0 0.00fF $ **FLOATING
C1979 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.t10 0 0.01fF $ **FLOATING
C1980 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n58 0 0.02fF $ **FLOATING
C1981 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n59 0 0.03fF $ **FLOATING
C1982 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n60 0 0.01fF $ **FLOATING
C1983 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n61 0 0.02fF $ **FLOATING
C1984 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n62 0 0.04fF $ **FLOATING
C1985 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n63 0 0.01fF $ **FLOATING
C1986 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n64 0 0.02fF $ **FLOATING
C1987 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n65 0 0.04fF $ **FLOATING
C1988 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n66 0 0.04fF $ **FLOATING
C1989 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n67 0 0.04fF $ **FLOATING
C1990 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n68 0 0.04fF $ **FLOATING
C1991 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n69 0 0.04fF $ **FLOATING
C1992 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n70 0 0.04fF $ **FLOATING
C1993 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n71 0 0.04fF $ **FLOATING
C1994 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n72 0 0.07fF $ **FLOATING
C1995 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n73 0 0.01fF $ **FLOATING
C1996 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n74 0 0.02fF $ **FLOATING
C1997 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n75 0 0.04fF $ **FLOATING
C1998 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB.n76 0 0.01fF $ **FLOATING
C1999 sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0 0.07fF
C2000 sky130_fd_sc_hd__dfrbp_1_0[17]/D 0 0.88fF
C2001 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t8 0 0.01fF $ **FLOATING
C2002 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t5 0 0.01fF $ **FLOATING
C2003 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n0 0 0.03fF $ **FLOATING
C2004 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t0 0 0.01fF $ **FLOATING
C2005 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n1 0 0.01fF $ **FLOATING
C2006 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n2 0 0.03fF $ **FLOATING
C2007 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n3 0 0.01fF $ **FLOATING
C2008 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n4 0 0.03fF $ **FLOATING
C2009 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n5 0 0.01fF $ **FLOATING
C2010 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n6 0 0.03fF $ **FLOATING
C2011 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n7 0 0.01fF $ **FLOATING
C2012 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n8 0 0.02fF $ **FLOATING
C2013 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n9 0 0.04fF $ **FLOATING
C2014 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n10 0 0.01fF $ **FLOATING
C2015 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n11 0 0.03fF $ **FLOATING
C2016 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n12 0 0.01fF $ **FLOATING
C2017 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n13 0 0.03fF $ **FLOATING
C2018 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n14 0 0.01fF $ **FLOATING
C2019 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t4 0 0.01fF $ **FLOATING
C2020 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t1 0 0.00fF $ **FLOATING
C2021 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n15 0 0.06fF $ **FLOATING
C2022 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n16 0 0.01fF $ **FLOATING
C2023 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n17 0 0.03fF $ **FLOATING
C2024 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n18 0 0.02fF $ **FLOATING
C2025 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n19 0 0.06fF $ **FLOATING
C2026 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n20 0 0.12fF $ **FLOATING
C2027 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n21 0 0.01fF $ **FLOATING
C2028 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n22 0 0.03fF $ **FLOATING
C2029 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n23 0 0.04fF $ **FLOATING
C2030 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n24 0 0.01fF $ **FLOATING
C2031 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n25 0 0.02fF $ **FLOATING
C2032 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n26 0 0.04fF $ **FLOATING
C2033 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t2 0 0.01fF $ **FLOATING
C2034 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n27 0 0.03fF $ **FLOATING
C2035 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n28 0 0.03fF $ **FLOATING
C2036 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t6 0 0.01fF $ **FLOATING
C2037 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n29 0 0.02fF $ **FLOATING
C2038 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n30 0 0.03fF $ **FLOATING
C2039 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n31 0 0.01fF $ **FLOATING
C2040 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n32 0 0.02fF $ **FLOATING
C2041 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n33 0 0.04fF $ **FLOATING
C2042 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n34 0 0.01fF $ **FLOATING
C2043 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n35 0 0.02fF $ **FLOATING
C2044 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n36 0 0.04fF $ **FLOATING
C2045 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t7 0 0.00fF $ **FLOATING
C2046 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t3 0 0.01fF $ **FLOATING
C2047 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n37 0 0.02fF $ **FLOATING
C2048 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n38 0 0.02fF $ **FLOATING
C2049 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n39 0 0.01fF $ **FLOATING
C2050 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n40 0 0.02fF $ **FLOATING
C2051 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n41 0 0.04fF $ **FLOATING
C2052 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n42 0 0.01fF $ **FLOATING
C2053 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n43 0 0.03fF $ **FLOATING
C2054 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n44 0 0.04fF $ **FLOATING
C2055 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n45 0 0.01fF $ **FLOATING
C2056 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n46 0 0.03fF $ **FLOATING
C2057 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n47 0 0.04fF $ **FLOATING
C2058 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n48 0 0.01fF $ **FLOATING
C2059 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n49 0 0.03fF $ **FLOATING
C2060 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n50 0 0.04fF $ **FLOATING
C2061 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t9 0 0.03fF $ **FLOATING
C2062 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n51 0 0.05fF $ **FLOATING
C2063 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n52 0 0.01fF $ **FLOATING
C2064 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n53 0 0.02fF $ **FLOATING
C2065 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n54 0 0.04fF $ **FLOATING
C2066 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n55 0 0.01fF $ **FLOATING
C2067 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n56 0 0.02fF $ **FLOATING
C2068 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n57 0 0.04fF $ **FLOATING
C2069 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t11 0 0.00fF $ **FLOATING
C2070 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.t10 0 0.01fF $ **FLOATING
C2071 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n58 0 0.02fF $ **FLOATING
C2072 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n59 0 0.03fF $ **FLOATING
C2073 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n60 0 0.01fF $ **FLOATING
C2074 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n61 0 0.02fF $ **FLOATING
C2075 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n62 0 0.04fF $ **FLOATING
C2076 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n63 0 0.01fF $ **FLOATING
C2077 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n64 0 0.02fF $ **FLOATING
C2078 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n65 0 0.04fF $ **FLOATING
C2079 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n66 0 0.04fF $ **FLOATING
C2080 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n67 0 0.04fF $ **FLOATING
C2081 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n68 0 0.04fF $ **FLOATING
C2082 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n69 0 0.04fF $ **FLOATING
C2083 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n70 0 0.04fF $ **FLOATING
C2084 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n71 0 0.04fF $ **FLOATING
C2085 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n72 0 0.07fF $ **FLOATING
C2086 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n73 0 0.01fF $ **FLOATING
C2087 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n74 0 0.02fF $ **FLOATING
C2088 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n75 0 0.04fF $ **FLOATING
C2089 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB.n76 0 0.01fF $ **FLOATING
C2090 sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0 0.07fF
C2091 sky130_fd_sc_hd__dfrbp_1_0[16]/D 0 2.14fF
C2092 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t8 0 0.01fF $ **FLOATING
C2093 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t5 0 0.01fF $ **FLOATING
C2094 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n0 0 0.03fF $ **FLOATING
C2095 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t0 0 0.01fF $ **FLOATING
C2096 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n1 0 0.01fF $ **FLOATING
C2097 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n2 0 0.03fF $ **FLOATING
C2098 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n3 0 0.01fF $ **FLOATING
C2099 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n4 0 0.03fF $ **FLOATING
C2100 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n5 0 0.01fF $ **FLOATING
C2101 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n6 0 0.03fF $ **FLOATING
C2102 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n7 0 0.01fF $ **FLOATING
C2103 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n8 0 0.02fF $ **FLOATING
C2104 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n9 0 0.04fF $ **FLOATING
C2105 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n10 0 0.01fF $ **FLOATING
C2106 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n11 0 0.03fF $ **FLOATING
C2107 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n12 0 0.01fF $ **FLOATING
C2108 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n13 0 0.03fF $ **FLOATING
C2109 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n14 0 0.01fF $ **FLOATING
C2110 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t4 0 0.01fF $ **FLOATING
C2111 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t1 0 0.00fF $ **FLOATING
C2112 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n15 0 0.06fF $ **FLOATING
C2113 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n16 0 0.01fF $ **FLOATING
C2114 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n17 0 0.03fF $ **FLOATING
C2115 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n18 0 0.02fF $ **FLOATING
C2116 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n19 0 0.06fF $ **FLOATING
C2117 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n20 0 0.12fF $ **FLOATING
C2118 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n21 0 0.01fF $ **FLOATING
C2119 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n22 0 0.03fF $ **FLOATING
C2120 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n23 0 0.04fF $ **FLOATING
C2121 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n24 0 0.01fF $ **FLOATING
C2122 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n25 0 0.02fF $ **FLOATING
C2123 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n26 0 0.04fF $ **FLOATING
C2124 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t2 0 0.01fF $ **FLOATING
C2125 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n27 0 0.03fF $ **FLOATING
C2126 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n28 0 0.03fF $ **FLOATING
C2127 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t6 0 0.01fF $ **FLOATING
C2128 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n29 0 0.02fF $ **FLOATING
C2129 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n30 0 0.03fF $ **FLOATING
C2130 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n31 0 0.01fF $ **FLOATING
C2131 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n32 0 0.02fF $ **FLOATING
C2132 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n33 0 0.04fF $ **FLOATING
C2133 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n34 0 0.01fF $ **FLOATING
C2134 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n35 0 0.02fF $ **FLOATING
C2135 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n36 0 0.04fF $ **FLOATING
C2136 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t7 0 0.00fF $ **FLOATING
C2137 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t3 0 0.01fF $ **FLOATING
C2138 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n37 0 0.02fF $ **FLOATING
C2139 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n38 0 0.02fF $ **FLOATING
C2140 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n39 0 0.01fF $ **FLOATING
C2141 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n40 0 0.02fF $ **FLOATING
C2142 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n41 0 0.04fF $ **FLOATING
C2143 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n42 0 0.01fF $ **FLOATING
C2144 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n43 0 0.03fF $ **FLOATING
C2145 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n44 0 0.04fF $ **FLOATING
C2146 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n45 0 0.01fF $ **FLOATING
C2147 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n46 0 0.03fF $ **FLOATING
C2148 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n47 0 0.04fF $ **FLOATING
C2149 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n48 0 0.01fF $ **FLOATING
C2150 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n49 0 0.03fF $ **FLOATING
C2151 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n50 0 0.04fF $ **FLOATING
C2152 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t9 0 0.03fF $ **FLOATING
C2153 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n51 0 0.05fF $ **FLOATING
C2154 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n52 0 0.01fF $ **FLOATING
C2155 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n53 0 0.02fF $ **FLOATING
C2156 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n54 0 0.04fF $ **FLOATING
C2157 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n55 0 0.01fF $ **FLOATING
C2158 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n56 0 0.02fF $ **FLOATING
C2159 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n57 0 0.04fF $ **FLOATING
C2160 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t11 0 0.00fF $ **FLOATING
C2161 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.t10 0 0.01fF $ **FLOATING
C2162 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n58 0 0.02fF $ **FLOATING
C2163 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n59 0 0.03fF $ **FLOATING
C2164 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n60 0 0.01fF $ **FLOATING
C2165 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n61 0 0.02fF $ **FLOATING
C2166 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n62 0 0.04fF $ **FLOATING
C2167 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n63 0 0.01fF $ **FLOATING
C2168 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n64 0 0.02fF $ **FLOATING
C2169 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n65 0 0.04fF $ **FLOATING
C2170 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n66 0 0.04fF $ **FLOATING
C2171 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n67 0 0.04fF $ **FLOATING
C2172 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n68 0 0.04fF $ **FLOATING
C2173 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n69 0 0.04fF $ **FLOATING
C2174 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n70 0 0.04fF $ **FLOATING
C2175 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n71 0 0.04fF $ **FLOATING
C2176 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n72 0 0.07fF $ **FLOATING
C2177 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n73 0 0.01fF $ **FLOATING
C2178 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n74 0 0.02fF $ **FLOATING
C2179 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n75 0 0.04fF $ **FLOATING
C2180 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB.n76 0 0.01fF $ **FLOATING
C2181 sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0 0.07fF
C2182 sky130_fd_sc_hd__dfrbp_1_0[15]/D 0 0.28fF
C2183 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t0 0 0.05fF
C2184 sky130_fd_sc_hd__dfrbp_1_0[16]/D.t1 0 0.06fF
C2185 sky130_fd_sc_hd__dfrbp_1_0[16]/D.n0 0 0.07fF $ **FLOATING
C2186 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t8 0 0.01fF $ **FLOATING
C2187 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t5 0 0.01fF $ **FLOATING
C2188 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n0 0 0.03fF $ **FLOATING
C2189 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t0 0 0.01fF $ **FLOATING
C2190 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n1 0 0.01fF $ **FLOATING
C2191 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n2 0 0.03fF $ **FLOATING
C2192 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n3 0 0.01fF $ **FLOATING
C2193 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n4 0 0.03fF $ **FLOATING
C2194 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n5 0 0.01fF $ **FLOATING
C2195 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n6 0 0.03fF $ **FLOATING
C2196 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n7 0 0.01fF $ **FLOATING
C2197 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n8 0 0.02fF $ **FLOATING
C2198 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n9 0 0.04fF $ **FLOATING
C2199 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n10 0 0.01fF $ **FLOATING
C2200 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n11 0 0.03fF $ **FLOATING
C2201 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n12 0 0.01fF $ **FLOATING
C2202 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n13 0 0.03fF $ **FLOATING
C2203 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n14 0 0.01fF $ **FLOATING
C2204 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t4 0 0.01fF $ **FLOATING
C2205 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t1 0 0.00fF $ **FLOATING
C2206 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n15 0 0.06fF $ **FLOATING
C2207 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n16 0 0.01fF $ **FLOATING
C2208 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n17 0 0.03fF $ **FLOATING
C2209 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n18 0 0.02fF $ **FLOATING
C2210 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n19 0 0.06fF $ **FLOATING
C2211 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n20 0 0.12fF $ **FLOATING
C2212 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n21 0 0.01fF $ **FLOATING
C2213 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n22 0 0.03fF $ **FLOATING
C2214 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n23 0 0.04fF $ **FLOATING
C2215 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n24 0 0.01fF $ **FLOATING
C2216 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n25 0 0.02fF $ **FLOATING
C2217 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n26 0 0.04fF $ **FLOATING
C2218 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t2 0 0.01fF $ **FLOATING
C2219 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n27 0 0.03fF $ **FLOATING
C2220 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n28 0 0.03fF $ **FLOATING
C2221 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t6 0 0.01fF $ **FLOATING
C2222 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n29 0 0.02fF $ **FLOATING
C2223 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n30 0 0.03fF $ **FLOATING
C2224 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n31 0 0.01fF $ **FLOATING
C2225 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n32 0 0.02fF $ **FLOATING
C2226 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n33 0 0.04fF $ **FLOATING
C2227 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n34 0 0.01fF $ **FLOATING
C2228 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n35 0 0.02fF $ **FLOATING
C2229 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n36 0 0.04fF $ **FLOATING
C2230 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t7 0 0.00fF $ **FLOATING
C2231 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t3 0 0.01fF $ **FLOATING
C2232 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n37 0 0.02fF $ **FLOATING
C2233 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n38 0 0.02fF $ **FLOATING
C2234 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n39 0 0.01fF $ **FLOATING
C2235 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n40 0 0.02fF $ **FLOATING
C2236 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n41 0 0.04fF $ **FLOATING
C2237 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n42 0 0.01fF $ **FLOATING
C2238 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n43 0 0.03fF $ **FLOATING
C2239 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n44 0 0.04fF $ **FLOATING
C2240 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n45 0 0.01fF $ **FLOATING
C2241 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n46 0 0.03fF $ **FLOATING
C2242 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n47 0 0.04fF $ **FLOATING
C2243 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n48 0 0.01fF $ **FLOATING
C2244 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n49 0 0.03fF $ **FLOATING
C2245 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n50 0 0.04fF $ **FLOATING
C2246 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t9 0 0.03fF $ **FLOATING
C2247 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n51 0 0.05fF $ **FLOATING
C2248 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n52 0 0.01fF $ **FLOATING
C2249 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n53 0 0.02fF $ **FLOATING
C2250 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n54 0 0.04fF $ **FLOATING
C2251 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n55 0 0.01fF $ **FLOATING
C2252 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n56 0 0.02fF $ **FLOATING
C2253 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n57 0 0.04fF $ **FLOATING
C2254 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t11 0 0.00fF $ **FLOATING
C2255 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.t10 0 0.01fF $ **FLOATING
C2256 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n58 0 0.02fF $ **FLOATING
C2257 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n59 0 0.03fF $ **FLOATING
C2258 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n60 0 0.01fF $ **FLOATING
C2259 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n61 0 0.02fF $ **FLOATING
C2260 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n62 0 0.04fF $ **FLOATING
C2261 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n63 0 0.01fF $ **FLOATING
C2262 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n64 0 0.02fF $ **FLOATING
C2263 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n65 0 0.04fF $ **FLOATING
C2264 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n66 0 0.04fF $ **FLOATING
C2265 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n67 0 0.04fF $ **FLOATING
C2266 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n68 0 0.04fF $ **FLOATING
C2267 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n69 0 0.04fF $ **FLOATING
C2268 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n70 0 0.04fF $ **FLOATING
C2269 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n71 0 0.04fF $ **FLOATING
C2270 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n72 0 0.07fF $ **FLOATING
C2271 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n73 0 0.01fF $ **FLOATING
C2272 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n74 0 0.02fF $ **FLOATING
C2273 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n75 0 0.04fF $ **FLOATING
C2274 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB.n76 0 0.01fF $ **FLOATING
C2275 sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0 0.07fF
C2276 sky130_fd_sc_hd__dfrbp_1_0[14]/D 0 1.69fF
C2277 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t8 0 0.01fF $ **FLOATING
C2278 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t5 0 0.01fF $ **FLOATING
C2279 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n0 0 0.03fF $ **FLOATING
C2280 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t0 0 0.01fF $ **FLOATING
C2281 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n1 0 0.01fF $ **FLOATING
C2282 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n2 0 0.03fF $ **FLOATING
C2283 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n3 0 0.01fF $ **FLOATING
C2284 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n4 0 0.03fF $ **FLOATING
C2285 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n5 0 0.01fF $ **FLOATING
C2286 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n6 0 0.03fF $ **FLOATING
C2287 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n7 0 0.01fF $ **FLOATING
C2288 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n8 0 0.02fF $ **FLOATING
C2289 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n9 0 0.04fF $ **FLOATING
C2290 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n10 0 0.01fF $ **FLOATING
C2291 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n11 0 0.03fF $ **FLOATING
C2292 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n12 0 0.01fF $ **FLOATING
C2293 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n13 0 0.03fF $ **FLOATING
C2294 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n14 0 0.01fF $ **FLOATING
C2295 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t4 0 0.01fF $ **FLOATING
C2296 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t1 0 0.00fF $ **FLOATING
C2297 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n15 0 0.06fF $ **FLOATING
C2298 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n16 0 0.01fF $ **FLOATING
C2299 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n17 0 0.03fF $ **FLOATING
C2300 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n18 0 0.02fF $ **FLOATING
C2301 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n19 0 0.06fF $ **FLOATING
C2302 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n20 0 0.12fF $ **FLOATING
C2303 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n21 0 0.01fF $ **FLOATING
C2304 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n22 0 0.03fF $ **FLOATING
C2305 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n23 0 0.04fF $ **FLOATING
C2306 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n24 0 0.01fF $ **FLOATING
C2307 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n25 0 0.02fF $ **FLOATING
C2308 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n26 0 0.04fF $ **FLOATING
C2309 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t2 0 0.01fF $ **FLOATING
C2310 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n27 0 0.03fF $ **FLOATING
C2311 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n28 0 0.03fF $ **FLOATING
C2312 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t6 0 0.01fF $ **FLOATING
C2313 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n29 0 0.02fF $ **FLOATING
C2314 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n30 0 0.03fF $ **FLOATING
C2315 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n31 0 0.01fF $ **FLOATING
C2316 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n32 0 0.02fF $ **FLOATING
C2317 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n33 0 0.04fF $ **FLOATING
C2318 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n34 0 0.01fF $ **FLOATING
C2319 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n35 0 0.02fF $ **FLOATING
C2320 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n36 0 0.04fF $ **FLOATING
C2321 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t7 0 0.00fF $ **FLOATING
C2322 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t3 0 0.01fF $ **FLOATING
C2323 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n37 0 0.02fF $ **FLOATING
C2324 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n38 0 0.02fF $ **FLOATING
C2325 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n39 0 0.01fF $ **FLOATING
C2326 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n40 0 0.02fF $ **FLOATING
C2327 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n41 0 0.04fF $ **FLOATING
C2328 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n42 0 0.01fF $ **FLOATING
C2329 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n43 0 0.03fF $ **FLOATING
C2330 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n44 0 0.04fF $ **FLOATING
C2331 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n45 0 0.01fF $ **FLOATING
C2332 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n46 0 0.03fF $ **FLOATING
C2333 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n47 0 0.04fF $ **FLOATING
C2334 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n48 0 0.01fF $ **FLOATING
C2335 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n49 0 0.03fF $ **FLOATING
C2336 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n50 0 0.04fF $ **FLOATING
C2337 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t9 0 0.03fF $ **FLOATING
C2338 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n51 0 0.05fF $ **FLOATING
C2339 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n52 0 0.01fF $ **FLOATING
C2340 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n53 0 0.02fF $ **FLOATING
C2341 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n54 0 0.04fF $ **FLOATING
C2342 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n55 0 0.01fF $ **FLOATING
C2343 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n56 0 0.02fF $ **FLOATING
C2344 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n57 0 0.04fF $ **FLOATING
C2345 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t11 0 0.00fF $ **FLOATING
C2346 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.t10 0 0.01fF $ **FLOATING
C2347 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n58 0 0.02fF $ **FLOATING
C2348 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n59 0 0.03fF $ **FLOATING
C2349 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n60 0 0.01fF $ **FLOATING
C2350 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n61 0 0.02fF $ **FLOATING
C2351 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n62 0 0.04fF $ **FLOATING
C2352 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n63 0 0.01fF $ **FLOATING
C2353 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n64 0 0.02fF $ **FLOATING
C2354 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n65 0 0.04fF $ **FLOATING
C2355 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n66 0 0.04fF $ **FLOATING
C2356 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n67 0 0.04fF $ **FLOATING
C2357 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n68 0 0.04fF $ **FLOATING
C2358 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n69 0 0.04fF $ **FLOATING
C2359 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n70 0 0.04fF $ **FLOATING
C2360 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n71 0 0.04fF $ **FLOATING
C2361 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n72 0 0.07fF $ **FLOATING
C2362 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n73 0 0.01fF $ **FLOATING
C2363 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n74 0 0.02fF $ **FLOATING
C2364 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n75 0 0.04fF $ **FLOATING
C2365 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB.n76 0 0.01fF $ **FLOATING
C2366 sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0 0.07fF
C2367 sky130_fd_sc_hd__dfrbp_1_0[13]/D 0 0.24fF
C2368 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t8 0 0.01fF $ **FLOATING
C2369 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t5 0 0.01fF $ **FLOATING
C2370 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n0 0 0.03fF $ **FLOATING
C2371 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t0 0 0.01fF $ **FLOATING
C2372 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n1 0 0.01fF $ **FLOATING
C2373 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n2 0 0.03fF $ **FLOATING
C2374 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n3 0 0.01fF $ **FLOATING
C2375 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n4 0 0.03fF $ **FLOATING
C2376 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n5 0 0.01fF $ **FLOATING
C2377 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n6 0 0.03fF $ **FLOATING
C2378 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n7 0 0.01fF $ **FLOATING
C2379 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n8 0 0.02fF $ **FLOATING
C2380 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n9 0 0.04fF $ **FLOATING
C2381 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n10 0 0.01fF $ **FLOATING
C2382 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n11 0 0.03fF $ **FLOATING
C2383 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n12 0 0.01fF $ **FLOATING
C2384 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n13 0 0.03fF $ **FLOATING
C2385 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n14 0 0.01fF $ **FLOATING
C2386 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t4 0 0.01fF $ **FLOATING
C2387 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t1 0 0.00fF $ **FLOATING
C2388 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n15 0 0.06fF $ **FLOATING
C2389 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n16 0 0.01fF $ **FLOATING
C2390 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n17 0 0.03fF $ **FLOATING
C2391 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n18 0 0.02fF $ **FLOATING
C2392 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n19 0 0.06fF $ **FLOATING
C2393 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n20 0 0.12fF $ **FLOATING
C2394 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n21 0 0.01fF $ **FLOATING
C2395 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n22 0 0.03fF $ **FLOATING
C2396 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n23 0 0.04fF $ **FLOATING
C2397 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n24 0 0.01fF $ **FLOATING
C2398 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n25 0 0.02fF $ **FLOATING
C2399 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n26 0 0.04fF $ **FLOATING
C2400 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t2 0 0.01fF $ **FLOATING
C2401 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n27 0 0.03fF $ **FLOATING
C2402 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n28 0 0.03fF $ **FLOATING
C2403 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t6 0 0.01fF $ **FLOATING
C2404 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n29 0 0.02fF $ **FLOATING
C2405 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n30 0 0.03fF $ **FLOATING
C2406 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n31 0 0.01fF $ **FLOATING
C2407 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n32 0 0.02fF $ **FLOATING
C2408 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n33 0 0.04fF $ **FLOATING
C2409 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n34 0 0.01fF $ **FLOATING
C2410 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n35 0 0.02fF $ **FLOATING
C2411 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n36 0 0.04fF $ **FLOATING
C2412 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t7 0 0.00fF $ **FLOATING
C2413 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t3 0 0.01fF $ **FLOATING
C2414 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n37 0 0.02fF $ **FLOATING
C2415 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n38 0 0.02fF $ **FLOATING
C2416 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n39 0 0.01fF $ **FLOATING
C2417 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n40 0 0.02fF $ **FLOATING
C2418 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n41 0 0.04fF $ **FLOATING
C2419 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n42 0 0.01fF $ **FLOATING
C2420 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n43 0 0.03fF $ **FLOATING
C2421 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n44 0 0.04fF $ **FLOATING
C2422 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n45 0 0.01fF $ **FLOATING
C2423 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n46 0 0.03fF $ **FLOATING
C2424 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n47 0 0.04fF $ **FLOATING
C2425 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n48 0 0.01fF $ **FLOATING
C2426 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n49 0 0.03fF $ **FLOATING
C2427 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n50 0 0.04fF $ **FLOATING
C2428 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t9 0 0.03fF $ **FLOATING
C2429 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n51 0 0.05fF $ **FLOATING
C2430 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n52 0 0.01fF $ **FLOATING
C2431 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n53 0 0.02fF $ **FLOATING
C2432 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n54 0 0.04fF $ **FLOATING
C2433 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n55 0 0.01fF $ **FLOATING
C2434 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n56 0 0.02fF $ **FLOATING
C2435 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n57 0 0.04fF $ **FLOATING
C2436 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t11 0 0.00fF $ **FLOATING
C2437 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.t10 0 0.01fF $ **FLOATING
C2438 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n58 0 0.02fF $ **FLOATING
C2439 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n59 0 0.03fF $ **FLOATING
C2440 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n60 0 0.01fF $ **FLOATING
C2441 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n61 0 0.02fF $ **FLOATING
C2442 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n62 0 0.04fF $ **FLOATING
C2443 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n63 0 0.01fF $ **FLOATING
C2444 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n64 0 0.02fF $ **FLOATING
C2445 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n65 0 0.04fF $ **FLOATING
C2446 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n66 0 0.04fF $ **FLOATING
C2447 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n67 0 0.04fF $ **FLOATING
C2448 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n68 0 0.04fF $ **FLOATING
C2449 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n69 0 0.04fF $ **FLOATING
C2450 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n70 0 0.04fF $ **FLOATING
C2451 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n71 0 0.04fF $ **FLOATING
C2452 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n72 0 0.07fF $ **FLOATING
C2453 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n73 0 0.01fF $ **FLOATING
C2454 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n74 0 0.02fF $ **FLOATING
C2455 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n75 0 0.04fF $ **FLOATING
C2456 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB.n76 0 0.01fF $ **FLOATING
C2457 sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0 0.07fF
C2458 sky130_fd_sc_hd__dfrbp_1_0[12]/D 0 1.60fF
C2459 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t8 0 0.01fF $ **FLOATING
C2460 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t5 0 0.01fF $ **FLOATING
C2461 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n0 0 0.03fF $ **FLOATING
C2462 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t0 0 0.01fF $ **FLOATING
C2463 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n1 0 0.01fF $ **FLOATING
C2464 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n2 0 0.03fF $ **FLOATING
C2465 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n3 0 0.01fF $ **FLOATING
C2466 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n4 0 0.03fF $ **FLOATING
C2467 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n5 0 0.01fF $ **FLOATING
C2468 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n6 0 0.03fF $ **FLOATING
C2469 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n7 0 0.01fF $ **FLOATING
C2470 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n8 0 0.02fF $ **FLOATING
C2471 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n9 0 0.04fF $ **FLOATING
C2472 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n10 0 0.01fF $ **FLOATING
C2473 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n11 0 0.03fF $ **FLOATING
C2474 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n12 0 0.01fF $ **FLOATING
C2475 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n13 0 0.03fF $ **FLOATING
C2476 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n14 0 0.01fF $ **FLOATING
C2477 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t4 0 0.01fF $ **FLOATING
C2478 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t1 0 0.00fF $ **FLOATING
C2479 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n15 0 0.06fF $ **FLOATING
C2480 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n16 0 0.01fF $ **FLOATING
C2481 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n17 0 0.03fF $ **FLOATING
C2482 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n18 0 0.02fF $ **FLOATING
C2483 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n19 0 0.06fF $ **FLOATING
C2484 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n20 0 0.12fF $ **FLOATING
C2485 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n21 0 0.01fF $ **FLOATING
C2486 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n22 0 0.03fF $ **FLOATING
C2487 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n23 0 0.04fF $ **FLOATING
C2488 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n24 0 0.01fF $ **FLOATING
C2489 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n25 0 0.02fF $ **FLOATING
C2490 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n26 0 0.04fF $ **FLOATING
C2491 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t2 0 0.01fF $ **FLOATING
C2492 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n27 0 0.03fF $ **FLOATING
C2493 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n28 0 0.03fF $ **FLOATING
C2494 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t6 0 0.01fF $ **FLOATING
C2495 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n29 0 0.02fF $ **FLOATING
C2496 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n30 0 0.03fF $ **FLOATING
C2497 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n31 0 0.01fF $ **FLOATING
C2498 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n32 0 0.02fF $ **FLOATING
C2499 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n33 0 0.04fF $ **FLOATING
C2500 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n34 0 0.01fF $ **FLOATING
C2501 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n35 0 0.02fF $ **FLOATING
C2502 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n36 0 0.04fF $ **FLOATING
C2503 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t7 0 0.00fF $ **FLOATING
C2504 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t3 0 0.01fF $ **FLOATING
C2505 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n37 0 0.02fF $ **FLOATING
C2506 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n38 0 0.02fF $ **FLOATING
C2507 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n39 0 0.01fF $ **FLOATING
C2508 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n40 0 0.02fF $ **FLOATING
C2509 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n41 0 0.04fF $ **FLOATING
C2510 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n42 0 0.01fF $ **FLOATING
C2511 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n43 0 0.03fF $ **FLOATING
C2512 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n44 0 0.04fF $ **FLOATING
C2513 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n45 0 0.01fF $ **FLOATING
C2514 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n46 0 0.03fF $ **FLOATING
C2515 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n47 0 0.04fF $ **FLOATING
C2516 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n48 0 0.01fF $ **FLOATING
C2517 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n49 0 0.03fF $ **FLOATING
C2518 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n50 0 0.04fF $ **FLOATING
C2519 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t9 0 0.03fF $ **FLOATING
C2520 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n51 0 0.05fF $ **FLOATING
C2521 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n52 0 0.01fF $ **FLOATING
C2522 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n53 0 0.02fF $ **FLOATING
C2523 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n54 0 0.04fF $ **FLOATING
C2524 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n55 0 0.01fF $ **FLOATING
C2525 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n56 0 0.02fF $ **FLOATING
C2526 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n57 0 0.04fF $ **FLOATING
C2527 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t11 0 0.00fF $ **FLOATING
C2528 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.t10 0 0.01fF $ **FLOATING
C2529 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n58 0 0.02fF $ **FLOATING
C2530 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n59 0 0.03fF $ **FLOATING
C2531 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n60 0 0.01fF $ **FLOATING
C2532 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n61 0 0.02fF $ **FLOATING
C2533 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n62 0 0.04fF $ **FLOATING
C2534 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n63 0 0.01fF $ **FLOATING
C2535 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n64 0 0.02fF $ **FLOATING
C2536 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n65 0 0.04fF $ **FLOATING
C2537 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n66 0 0.04fF $ **FLOATING
C2538 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n67 0 0.04fF $ **FLOATING
C2539 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n68 0 0.04fF $ **FLOATING
C2540 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n69 0 0.04fF $ **FLOATING
C2541 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n70 0 0.04fF $ **FLOATING
C2542 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n71 0 0.04fF $ **FLOATING
C2543 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n72 0 0.07fF $ **FLOATING
C2544 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n73 0 0.01fF $ **FLOATING
C2545 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n74 0 0.02fF $ **FLOATING
C2546 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n75 0 0.04fF $ **FLOATING
C2547 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB.n76 0 0.01fF $ **FLOATING
C2548 sky130_fd_sc_hd__dfrbp_1_0[12]/Q 0 0.07fF
C2549 sky130_fd_sc_hd__dfrbp_1_0[11]/D 0 0.23fF
C2550 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t8 0 0.01fF $ **FLOATING
C2551 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t5 0 0.01fF $ **FLOATING
C2552 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n0 0 0.03fF $ **FLOATING
C2553 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t0 0 0.01fF $ **FLOATING
C2554 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n1 0 0.01fF $ **FLOATING
C2555 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n2 0 0.03fF $ **FLOATING
C2556 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n3 0 0.01fF $ **FLOATING
C2557 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n4 0 0.03fF $ **FLOATING
C2558 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n5 0 0.01fF $ **FLOATING
C2559 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n6 0 0.03fF $ **FLOATING
C2560 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n7 0 0.01fF $ **FLOATING
C2561 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n8 0 0.02fF $ **FLOATING
C2562 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n9 0 0.04fF $ **FLOATING
C2563 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n10 0 0.01fF $ **FLOATING
C2564 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n11 0 0.03fF $ **FLOATING
C2565 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n12 0 0.01fF $ **FLOATING
C2566 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n13 0 0.03fF $ **FLOATING
C2567 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n14 0 0.01fF $ **FLOATING
C2568 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t4 0 0.01fF $ **FLOATING
C2569 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t1 0 0.00fF $ **FLOATING
C2570 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n15 0 0.06fF $ **FLOATING
C2571 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n16 0 0.01fF $ **FLOATING
C2572 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n17 0 0.03fF $ **FLOATING
C2573 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n18 0 0.02fF $ **FLOATING
C2574 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n19 0 0.06fF $ **FLOATING
C2575 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n20 0 0.12fF $ **FLOATING
C2576 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n21 0 0.01fF $ **FLOATING
C2577 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n22 0 0.03fF $ **FLOATING
C2578 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n23 0 0.04fF $ **FLOATING
C2579 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n24 0 0.01fF $ **FLOATING
C2580 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n25 0 0.02fF $ **FLOATING
C2581 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n26 0 0.04fF $ **FLOATING
C2582 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t2 0 0.01fF $ **FLOATING
C2583 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n27 0 0.03fF $ **FLOATING
C2584 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n28 0 0.03fF $ **FLOATING
C2585 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t6 0 0.01fF $ **FLOATING
C2586 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n29 0 0.02fF $ **FLOATING
C2587 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n30 0 0.03fF $ **FLOATING
C2588 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n31 0 0.01fF $ **FLOATING
C2589 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n32 0 0.02fF $ **FLOATING
C2590 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n33 0 0.04fF $ **FLOATING
C2591 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n34 0 0.01fF $ **FLOATING
C2592 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n35 0 0.02fF $ **FLOATING
C2593 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n36 0 0.04fF $ **FLOATING
C2594 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t7 0 0.00fF $ **FLOATING
C2595 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t3 0 0.01fF $ **FLOATING
C2596 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n37 0 0.02fF $ **FLOATING
C2597 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n38 0 0.02fF $ **FLOATING
C2598 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n39 0 0.01fF $ **FLOATING
C2599 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n40 0 0.02fF $ **FLOATING
C2600 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n41 0 0.04fF $ **FLOATING
C2601 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n42 0 0.01fF $ **FLOATING
C2602 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n43 0 0.03fF $ **FLOATING
C2603 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n44 0 0.04fF $ **FLOATING
C2604 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n45 0 0.01fF $ **FLOATING
C2605 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n46 0 0.03fF $ **FLOATING
C2606 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n47 0 0.04fF $ **FLOATING
C2607 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n48 0 0.01fF $ **FLOATING
C2608 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n49 0 0.03fF $ **FLOATING
C2609 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n50 0 0.04fF $ **FLOATING
C2610 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t9 0 0.03fF $ **FLOATING
C2611 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n51 0 0.05fF $ **FLOATING
C2612 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n52 0 0.01fF $ **FLOATING
C2613 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n53 0 0.02fF $ **FLOATING
C2614 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n54 0 0.04fF $ **FLOATING
C2615 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n55 0 0.01fF $ **FLOATING
C2616 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n56 0 0.02fF $ **FLOATING
C2617 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n57 0 0.04fF $ **FLOATING
C2618 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t11 0 0.00fF $ **FLOATING
C2619 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.t10 0 0.01fF $ **FLOATING
C2620 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n58 0 0.02fF $ **FLOATING
C2621 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n59 0 0.03fF $ **FLOATING
C2622 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n60 0 0.01fF $ **FLOATING
C2623 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n61 0 0.02fF $ **FLOATING
C2624 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n62 0 0.04fF $ **FLOATING
C2625 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n63 0 0.01fF $ **FLOATING
C2626 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n64 0 0.02fF $ **FLOATING
C2627 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n65 0 0.04fF $ **FLOATING
C2628 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n66 0 0.04fF $ **FLOATING
C2629 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n67 0 0.04fF $ **FLOATING
C2630 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n68 0 0.04fF $ **FLOATING
C2631 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n69 0 0.04fF $ **FLOATING
C2632 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n70 0 0.04fF $ **FLOATING
C2633 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n71 0 0.04fF $ **FLOATING
C2634 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n72 0 0.07fF $ **FLOATING
C2635 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n73 0 0.01fF $ **FLOATING
C2636 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n74 0 0.02fF $ **FLOATING
C2637 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n75 0 0.04fF $ **FLOATING
C2638 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB.n76 0 0.01fF $ **FLOATING
C2639 sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0 0.07fF
C2640 sky130_fd_sc_hd__dfrbp_1_0[10]/D 0 1.76fF
C2641 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t8 0 0.01fF $ **FLOATING
C2642 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t5 0 0.01fF $ **FLOATING
C2643 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n0 0 0.03fF $ **FLOATING
C2644 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t0 0 0.01fF $ **FLOATING
C2645 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n1 0 0.01fF $ **FLOATING
C2646 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n2 0 0.03fF $ **FLOATING
C2647 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n3 0 0.01fF $ **FLOATING
C2648 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n4 0 0.03fF $ **FLOATING
C2649 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n5 0 0.01fF $ **FLOATING
C2650 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n6 0 0.03fF $ **FLOATING
C2651 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n7 0 0.01fF $ **FLOATING
C2652 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n8 0 0.02fF $ **FLOATING
C2653 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n9 0 0.04fF $ **FLOATING
C2654 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n10 0 0.01fF $ **FLOATING
C2655 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n11 0 0.03fF $ **FLOATING
C2656 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n12 0 0.01fF $ **FLOATING
C2657 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n13 0 0.03fF $ **FLOATING
C2658 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n14 0 0.01fF $ **FLOATING
C2659 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t4 0 0.01fF $ **FLOATING
C2660 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t1 0 0.00fF $ **FLOATING
C2661 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n15 0 0.06fF $ **FLOATING
C2662 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n16 0 0.01fF $ **FLOATING
C2663 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n17 0 0.03fF $ **FLOATING
C2664 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n18 0 0.02fF $ **FLOATING
C2665 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n19 0 0.06fF $ **FLOATING
C2666 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n20 0 0.12fF $ **FLOATING
C2667 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n21 0 0.01fF $ **FLOATING
C2668 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n22 0 0.03fF $ **FLOATING
C2669 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n23 0 0.04fF $ **FLOATING
C2670 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n24 0 0.01fF $ **FLOATING
C2671 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n25 0 0.02fF $ **FLOATING
C2672 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n26 0 0.04fF $ **FLOATING
C2673 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t2 0 0.01fF $ **FLOATING
C2674 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n27 0 0.03fF $ **FLOATING
C2675 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n28 0 0.03fF $ **FLOATING
C2676 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t6 0 0.01fF $ **FLOATING
C2677 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n29 0 0.02fF $ **FLOATING
C2678 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n30 0 0.03fF $ **FLOATING
C2679 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n31 0 0.01fF $ **FLOATING
C2680 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n32 0 0.02fF $ **FLOATING
C2681 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n33 0 0.04fF $ **FLOATING
C2682 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n34 0 0.01fF $ **FLOATING
C2683 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n35 0 0.02fF $ **FLOATING
C2684 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n36 0 0.04fF $ **FLOATING
C2685 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t7 0 0.00fF $ **FLOATING
C2686 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t3 0 0.01fF $ **FLOATING
C2687 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n37 0 0.02fF $ **FLOATING
C2688 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n38 0 0.02fF $ **FLOATING
C2689 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n39 0 0.01fF $ **FLOATING
C2690 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n40 0 0.02fF $ **FLOATING
C2691 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n41 0 0.04fF $ **FLOATING
C2692 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n42 0 0.01fF $ **FLOATING
C2693 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n43 0 0.03fF $ **FLOATING
C2694 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n44 0 0.04fF $ **FLOATING
C2695 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n45 0 0.01fF $ **FLOATING
C2696 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n46 0 0.03fF $ **FLOATING
C2697 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n47 0 0.04fF $ **FLOATING
C2698 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n48 0 0.01fF $ **FLOATING
C2699 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n49 0 0.03fF $ **FLOATING
C2700 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n50 0 0.04fF $ **FLOATING
C2701 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t9 0 0.03fF $ **FLOATING
C2702 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n51 0 0.05fF $ **FLOATING
C2703 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n52 0 0.01fF $ **FLOATING
C2704 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n53 0 0.02fF $ **FLOATING
C2705 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n54 0 0.04fF $ **FLOATING
C2706 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n55 0 0.01fF $ **FLOATING
C2707 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n56 0 0.02fF $ **FLOATING
C2708 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n57 0 0.04fF $ **FLOATING
C2709 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t11 0 0.00fF $ **FLOATING
C2710 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.t10 0 0.01fF $ **FLOATING
C2711 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n58 0 0.02fF $ **FLOATING
C2712 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n59 0 0.03fF $ **FLOATING
C2713 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n60 0 0.01fF $ **FLOATING
C2714 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n61 0 0.02fF $ **FLOATING
C2715 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n62 0 0.04fF $ **FLOATING
C2716 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n63 0 0.01fF $ **FLOATING
C2717 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n64 0 0.02fF $ **FLOATING
C2718 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n65 0 0.04fF $ **FLOATING
C2719 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n66 0 0.04fF $ **FLOATING
C2720 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n67 0 0.04fF $ **FLOATING
C2721 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n68 0 0.04fF $ **FLOATING
C2722 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n69 0 0.04fF $ **FLOATING
C2723 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n70 0 0.04fF $ **FLOATING
C2724 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n71 0 0.04fF $ **FLOATING
C2725 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n72 0 0.07fF $ **FLOATING
C2726 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n73 0 0.01fF $ **FLOATING
C2727 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n74 0 0.02fF $ **FLOATING
C2728 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n75 0 0.04fF $ **FLOATING
C2729 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB.n76 0 0.01fF $ **FLOATING
C2730 sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0 0.07fF
C2731 sky130_fd_sc_hd__dfrbp_1_0[9]/D 0 0.45fF
C2732 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t8 0 0.01fF $ **FLOATING
C2733 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t5 0 0.01fF $ **FLOATING
C2734 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n0 0 0.03fF $ **FLOATING
C2735 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t0 0 0.01fF $ **FLOATING
C2736 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n1 0 0.01fF $ **FLOATING
C2737 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n2 0 0.03fF $ **FLOATING
C2738 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n3 0 0.01fF $ **FLOATING
C2739 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n4 0 0.03fF $ **FLOATING
C2740 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n5 0 0.01fF $ **FLOATING
C2741 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n6 0 0.03fF $ **FLOATING
C2742 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n7 0 0.01fF $ **FLOATING
C2743 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n8 0 0.02fF $ **FLOATING
C2744 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n9 0 0.04fF $ **FLOATING
C2745 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n10 0 0.01fF $ **FLOATING
C2746 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n11 0 0.03fF $ **FLOATING
C2747 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n12 0 0.01fF $ **FLOATING
C2748 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n13 0 0.03fF $ **FLOATING
C2749 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n14 0 0.01fF $ **FLOATING
C2750 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t4 0 0.01fF $ **FLOATING
C2751 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t1 0 0.00fF $ **FLOATING
C2752 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n15 0 0.06fF $ **FLOATING
C2753 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n16 0 0.01fF $ **FLOATING
C2754 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n17 0 0.03fF $ **FLOATING
C2755 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n18 0 0.02fF $ **FLOATING
C2756 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n19 0 0.06fF $ **FLOATING
C2757 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n20 0 0.12fF $ **FLOATING
C2758 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n21 0 0.01fF $ **FLOATING
C2759 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n22 0 0.03fF $ **FLOATING
C2760 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n23 0 0.04fF $ **FLOATING
C2761 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n24 0 0.01fF $ **FLOATING
C2762 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n25 0 0.02fF $ **FLOATING
C2763 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n26 0 0.04fF $ **FLOATING
C2764 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t2 0 0.01fF $ **FLOATING
C2765 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n27 0 0.03fF $ **FLOATING
C2766 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n28 0 0.03fF $ **FLOATING
C2767 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t6 0 0.01fF $ **FLOATING
C2768 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n29 0 0.02fF $ **FLOATING
C2769 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n30 0 0.03fF $ **FLOATING
C2770 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n31 0 0.01fF $ **FLOATING
C2771 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n32 0 0.02fF $ **FLOATING
C2772 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n33 0 0.04fF $ **FLOATING
C2773 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n34 0 0.01fF $ **FLOATING
C2774 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n35 0 0.02fF $ **FLOATING
C2775 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n36 0 0.04fF $ **FLOATING
C2776 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t7 0 0.00fF $ **FLOATING
C2777 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t3 0 0.01fF $ **FLOATING
C2778 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n37 0 0.02fF $ **FLOATING
C2779 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n38 0 0.02fF $ **FLOATING
C2780 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n39 0 0.01fF $ **FLOATING
C2781 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n40 0 0.02fF $ **FLOATING
C2782 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n41 0 0.04fF $ **FLOATING
C2783 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n42 0 0.01fF $ **FLOATING
C2784 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n43 0 0.03fF $ **FLOATING
C2785 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n44 0 0.04fF $ **FLOATING
C2786 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n45 0 0.01fF $ **FLOATING
C2787 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n46 0 0.03fF $ **FLOATING
C2788 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n47 0 0.04fF $ **FLOATING
C2789 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n48 0 0.01fF $ **FLOATING
C2790 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n49 0 0.03fF $ **FLOATING
C2791 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n50 0 0.04fF $ **FLOATING
C2792 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t9 0 0.03fF $ **FLOATING
C2793 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n51 0 0.05fF $ **FLOATING
C2794 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n52 0 0.01fF $ **FLOATING
C2795 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n53 0 0.02fF $ **FLOATING
C2796 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n54 0 0.04fF $ **FLOATING
C2797 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n55 0 0.01fF $ **FLOATING
C2798 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n56 0 0.02fF $ **FLOATING
C2799 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n57 0 0.04fF $ **FLOATING
C2800 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t11 0 0.00fF $ **FLOATING
C2801 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.t10 0 0.01fF $ **FLOATING
C2802 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n58 0 0.02fF $ **FLOATING
C2803 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n59 0 0.03fF $ **FLOATING
C2804 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n60 0 0.01fF $ **FLOATING
C2805 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n61 0 0.02fF $ **FLOATING
C2806 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n62 0 0.04fF $ **FLOATING
C2807 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n63 0 0.01fF $ **FLOATING
C2808 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n64 0 0.02fF $ **FLOATING
C2809 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n65 0 0.04fF $ **FLOATING
C2810 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n66 0 0.04fF $ **FLOATING
C2811 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n67 0 0.04fF $ **FLOATING
C2812 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n68 0 0.04fF $ **FLOATING
C2813 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n69 0 0.04fF $ **FLOATING
C2814 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n70 0 0.04fF $ **FLOATING
C2815 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n71 0 0.04fF $ **FLOATING
C2816 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n72 0 0.07fF $ **FLOATING
C2817 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n73 0 0.01fF $ **FLOATING
C2818 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n74 0 0.02fF $ **FLOATING
C2819 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n75 0 0.04fF $ **FLOATING
C2820 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB.n76 0 0.01fF $ **FLOATING
C2821 sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0 0.07fF
C2822 sky130_fd_sc_hd__dfrbp_1_0[8]/D 0 1.76fF
C2823 VDD.t8 0 0.04fF
C2824 VDD.t5 0 0.02fF
C2825 VDD.n0 0 0.05fF $ **FLOATING
C2826 VDD.t0 0 0.02fF
C2827 VDD.n1 0 0.03fF $ **FLOATING
C2828 VDD.n2 0 0.05fF $ **FLOATING
C2829 VDD.n3 0 0.06fF $ **FLOATING
C2830 VDD.n4 0 0.04fF $ **FLOATING
C2831 VDD.n5 0 0.04fF $ **FLOATING
C2832 VDD.n6 0 0.04fF $ **FLOATING
C2833 VDD.n7 0 0.05fF $ **FLOATING
C2834 VDD.n8 0 0.03fF $ **FLOATING
C2835 VDD.n9 0 0.06fF $ **FLOATING
C2836 VDD.n10 0 0.05fF $ **FLOATING
C2837 VDD.n11 0 0.04fF $ **FLOATING
C2838 VDD.n12 0 0.05fF $ **FLOATING
C2839 VDD.n13 0 0.04fF $ **FLOATING
C2840 VDD.n14 0 0.05fF $ **FLOATING
C2841 VDD.t4 0 0.02fF
C2842 VDD.t1 0 0.01fF
C2843 VDD.n15 0 0.08fF $ **FLOATING
C2844 VDD.n16 0 0.08fF $ **FLOATING
C2845 VDD.n17 0 0.04fF $ **FLOATING
C2846 VDD.n18 0 0.05fF $ **FLOATING
C2847 VDD.n19 0 0.09fF $ **FLOATING
C2848 VDD.n20 0 0.19fF $ **FLOATING
C2849 VDD.n21 0 0.15fF $ **FLOATING
C2850 VDD.n22 0 0.04fF $ **FLOATING
C2851 VDD.n23 0 0.07fF $ **FLOATING
C2852 VDD.n24 0 0.06fF $ **FLOATING
C2853 VDD.n25 0 0.04fF $ **FLOATING
C2854 VDD.n26 0 0.06fF $ **FLOATING
C2855 VDD.t2 0 0.02fF
C2856 VDD.n27 0 0.08fF $ **FLOATING
C2857 VDD.n28 0 0.07fF $ **FLOATING
C2858 VDD.t6 0 0.02fF
C2859 VDD.n29 0 0.05fF $ **FLOATING
C2860 VDD.n30 0 0.05fF $ **FLOATING
C2861 VDD.n31 0 0.05fF $ **FLOATING
C2862 VDD.n32 0 0.04fF $ **FLOATING
C2863 VDD.n33 0 0.07fF $ **FLOATING
C2864 VDD.n34 0 0.06fF $ **FLOATING
C2865 VDD.n35 0 0.04fF $ **FLOATING
C2866 VDD.n36 0 0.06fF $ **FLOATING
C2867 VDD.t7 0 0.01fF
C2868 VDD.t3 0 0.02fF
C2869 VDD.n37 0 0.06fF $ **FLOATING
C2870 VDD.n38 0 0.05fF $ **FLOATING
C2871 VDD.n39 0 0.04fF $ **FLOATING
C2872 VDD.n40 0 0.03fF $ **FLOATING
C2873 VDD.n41 0 0.06fF $ **FLOATING
C2874 VDD.n42 0 0.06fF $ **FLOATING
C2875 VDD.n43 0 0.04fF $ **FLOATING
C2876 VDD.n44 0 0.07fF $ **FLOATING
C2877 VDD.n45 0 0.06fF $ **FLOATING
C2878 VDD.n46 0 0.04fF $ **FLOATING
C2879 VDD.n47 0 0.07fF $ **FLOATING
C2880 VDD.n48 0 0.06fF $ **FLOATING
C2881 VDD.n49 0 0.04fF $ **FLOATING
C2882 VDD.n50 0 0.07fF $ **FLOATING
C2883 VDD.t9 0 0.03fF
C2884 VDD.n51 0 0.10fF $ **FLOATING
C2885 VDD.n52 0 0.07fF $ **FLOATING
C2886 VDD.n53 0 0.03fF $ **FLOATING
C2887 VDD.n54 0 0.06fF $ **FLOATING
C2888 VDD.n55 0 0.06fF $ **FLOATING
C2889 VDD.n56 0 0.04fF $ **FLOATING
C2890 VDD.n57 0 0.06fF $ **FLOATING
C2891 VDD.t11 0 0.02fF
C2892 VDD.t10 0 0.02fF
C2893 VDD.n58 0 0.06fF $ **FLOATING
C2894 VDD.n59 0 0.05fF $ **FLOATING
C2895 VDD.n60 0 0.05fF $ **FLOATING
C2896 VDD.n61 0 0.04fF $ **FLOATING
C2897 VDD.n62 0 0.06fF $ **FLOATING
C2898 VDD.n63 0 0.06fF $ **FLOATING
C2899 VDD.n64 0 0.04fF $ **FLOATING
C2900 VDD.n65 0 0.06fF $ **FLOATING
C2901 VDD.n66 0 0.08fF $ **FLOATING
C2902 VDD.n67 0 0.05fF $ **FLOATING
C2903 VDD.n68 0 0.07fF $ **FLOATING
C2904 VDD.n69 0 0.08fF $ **FLOATING
C2905 VDD.n70 0 0.05fF $ **FLOATING
C2906 VDD.n71 0 0.07fF $ **FLOATING
C2907 VDD.n72 0 0.12fF $ **FLOATING
C2908 VDD.n73 0 0.03fF $ **FLOATING
C2909 VDD.n74 0 0.05fF $ **FLOATING
C2910 VDD.n75 0 0.08fF $ **FLOATING
C2911 VDD.n76 0 0.06fF $ **FLOATING
C2912 sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0 0.07fF
C2913 sky130_fd_sc_hd__dfrbp_1_0[7]/D 0 0.10fF
C2914 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t8 0 0.01fF $ **FLOATING
C2915 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t5 0 0.01fF $ **FLOATING
C2916 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n0 0 0.03fF $ **FLOATING
C2917 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t0 0 0.01fF $ **FLOATING
C2918 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n1 0 0.01fF $ **FLOATING
C2919 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n2 0 0.03fF $ **FLOATING
C2920 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n3 0 0.01fF $ **FLOATING
C2921 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n4 0 0.03fF $ **FLOATING
C2922 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n5 0 0.01fF $ **FLOATING
C2923 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n6 0 0.03fF $ **FLOATING
C2924 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n7 0 0.01fF $ **FLOATING
C2925 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n8 0 0.02fF $ **FLOATING
C2926 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n9 0 0.04fF $ **FLOATING
C2927 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n10 0 0.01fF $ **FLOATING
C2928 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n11 0 0.03fF $ **FLOATING
C2929 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n12 0 0.01fF $ **FLOATING
C2930 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n13 0 0.03fF $ **FLOATING
C2931 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n14 0 0.01fF $ **FLOATING
C2932 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t4 0 0.01fF $ **FLOATING
C2933 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t1 0 0.00fF $ **FLOATING
C2934 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n15 0 0.06fF $ **FLOATING
C2935 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n16 0 0.01fF $ **FLOATING
C2936 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n17 0 0.03fF $ **FLOATING
C2937 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n18 0 0.02fF $ **FLOATING
C2938 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n19 0 0.06fF $ **FLOATING
C2939 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n20 0 0.12fF $ **FLOATING
C2940 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n21 0 0.01fF $ **FLOATING
C2941 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n22 0 0.03fF $ **FLOATING
C2942 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n23 0 0.04fF $ **FLOATING
C2943 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n24 0 0.01fF $ **FLOATING
C2944 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n25 0 0.02fF $ **FLOATING
C2945 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n26 0 0.04fF $ **FLOATING
C2946 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t2 0 0.01fF $ **FLOATING
C2947 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n27 0 0.03fF $ **FLOATING
C2948 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n28 0 0.03fF $ **FLOATING
C2949 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t6 0 0.01fF $ **FLOATING
C2950 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n29 0 0.02fF $ **FLOATING
C2951 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n30 0 0.03fF $ **FLOATING
C2952 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n31 0 0.01fF $ **FLOATING
C2953 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n32 0 0.02fF $ **FLOATING
C2954 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n33 0 0.04fF $ **FLOATING
C2955 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n34 0 0.01fF $ **FLOATING
C2956 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n35 0 0.02fF $ **FLOATING
C2957 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n36 0 0.04fF $ **FLOATING
C2958 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t7 0 0.00fF $ **FLOATING
C2959 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t3 0 0.01fF $ **FLOATING
C2960 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n37 0 0.02fF $ **FLOATING
C2961 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n38 0 0.02fF $ **FLOATING
C2962 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n39 0 0.01fF $ **FLOATING
C2963 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n40 0 0.02fF $ **FLOATING
C2964 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n41 0 0.04fF $ **FLOATING
C2965 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n42 0 0.01fF $ **FLOATING
C2966 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n43 0 0.03fF $ **FLOATING
C2967 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n44 0 0.04fF $ **FLOATING
C2968 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n45 0 0.01fF $ **FLOATING
C2969 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n46 0 0.03fF $ **FLOATING
C2970 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n47 0 0.04fF $ **FLOATING
C2971 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n48 0 0.01fF $ **FLOATING
C2972 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n49 0 0.03fF $ **FLOATING
C2973 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n50 0 0.04fF $ **FLOATING
C2974 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t9 0 0.03fF $ **FLOATING
C2975 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n51 0 0.05fF $ **FLOATING
C2976 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n52 0 0.01fF $ **FLOATING
C2977 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n53 0 0.02fF $ **FLOATING
C2978 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n54 0 0.04fF $ **FLOATING
C2979 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n55 0 0.01fF $ **FLOATING
C2980 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n56 0 0.02fF $ **FLOATING
C2981 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n57 0 0.04fF $ **FLOATING
C2982 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t11 0 0.00fF $ **FLOATING
C2983 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.t10 0 0.01fF $ **FLOATING
C2984 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n58 0 0.02fF $ **FLOATING
C2985 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n59 0 0.03fF $ **FLOATING
C2986 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n60 0 0.01fF $ **FLOATING
C2987 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n61 0 0.02fF $ **FLOATING
C2988 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n62 0 0.04fF $ **FLOATING
C2989 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n63 0 0.01fF $ **FLOATING
C2990 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n64 0 0.02fF $ **FLOATING
C2991 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n65 0 0.04fF $ **FLOATING
C2992 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n66 0 0.04fF $ **FLOATING
C2993 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n67 0 0.04fF $ **FLOATING
C2994 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n68 0 0.04fF $ **FLOATING
C2995 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n69 0 0.04fF $ **FLOATING
C2996 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n70 0 0.04fF $ **FLOATING
C2997 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n71 0 0.04fF $ **FLOATING
C2998 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n72 0 0.07fF $ **FLOATING
C2999 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n73 0 0.01fF $ **FLOATING
C3000 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n74 0 0.02fF $ **FLOATING
C3001 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n75 0 0.04fF $ **FLOATING
C3002 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB.n76 0 0.01fF $ **FLOATING
C3003 sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0 0.07fF
C3004 sky130_fd_sc_hd__dfrbp_1_0[6]/D 0 1.59fF
C3005 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t8 0 0.01fF $ **FLOATING
C3006 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t5 0 0.01fF $ **FLOATING
C3007 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n0 0 0.03fF $ **FLOATING
C3008 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t0 0 0.01fF $ **FLOATING
C3009 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n1 0 0.01fF $ **FLOATING
C3010 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n2 0 0.03fF $ **FLOATING
C3011 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n3 0 0.01fF $ **FLOATING
C3012 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n4 0 0.03fF $ **FLOATING
C3013 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n5 0 0.01fF $ **FLOATING
C3014 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n6 0 0.03fF $ **FLOATING
C3015 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n7 0 0.01fF $ **FLOATING
C3016 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n8 0 0.02fF $ **FLOATING
C3017 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n9 0 0.04fF $ **FLOATING
C3018 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n10 0 0.01fF $ **FLOATING
C3019 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n11 0 0.03fF $ **FLOATING
C3020 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n12 0 0.01fF $ **FLOATING
C3021 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n13 0 0.03fF $ **FLOATING
C3022 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n14 0 0.01fF $ **FLOATING
C3023 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t4 0 0.01fF $ **FLOATING
C3024 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t1 0 0.00fF $ **FLOATING
C3025 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n15 0 0.06fF $ **FLOATING
C3026 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n16 0 0.01fF $ **FLOATING
C3027 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n17 0 0.03fF $ **FLOATING
C3028 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n18 0 0.02fF $ **FLOATING
C3029 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n19 0 0.06fF $ **FLOATING
C3030 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n20 0 0.12fF $ **FLOATING
C3031 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n21 0 0.01fF $ **FLOATING
C3032 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n22 0 0.03fF $ **FLOATING
C3033 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n23 0 0.04fF $ **FLOATING
C3034 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n24 0 0.01fF $ **FLOATING
C3035 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n25 0 0.02fF $ **FLOATING
C3036 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n26 0 0.04fF $ **FLOATING
C3037 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t2 0 0.01fF $ **FLOATING
C3038 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n27 0 0.03fF $ **FLOATING
C3039 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n28 0 0.03fF $ **FLOATING
C3040 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t6 0 0.01fF $ **FLOATING
C3041 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n29 0 0.02fF $ **FLOATING
C3042 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n30 0 0.03fF $ **FLOATING
C3043 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n31 0 0.01fF $ **FLOATING
C3044 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n32 0 0.02fF $ **FLOATING
C3045 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n33 0 0.04fF $ **FLOATING
C3046 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n34 0 0.01fF $ **FLOATING
C3047 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n35 0 0.02fF $ **FLOATING
C3048 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n36 0 0.04fF $ **FLOATING
C3049 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t7 0 0.00fF $ **FLOATING
C3050 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t3 0 0.01fF $ **FLOATING
C3051 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n37 0 0.02fF $ **FLOATING
C3052 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n38 0 0.02fF $ **FLOATING
C3053 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n39 0 0.01fF $ **FLOATING
C3054 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n40 0 0.02fF $ **FLOATING
C3055 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n41 0 0.04fF $ **FLOATING
C3056 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n42 0 0.01fF $ **FLOATING
C3057 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n43 0 0.03fF $ **FLOATING
C3058 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n44 0 0.04fF $ **FLOATING
C3059 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n45 0 0.01fF $ **FLOATING
C3060 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n46 0 0.03fF $ **FLOATING
C3061 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n47 0 0.04fF $ **FLOATING
C3062 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n48 0 0.01fF $ **FLOATING
C3063 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n49 0 0.03fF $ **FLOATING
C3064 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n50 0 0.04fF $ **FLOATING
C3065 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t9 0 0.03fF $ **FLOATING
C3066 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n51 0 0.05fF $ **FLOATING
C3067 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n52 0 0.01fF $ **FLOATING
C3068 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n53 0 0.02fF $ **FLOATING
C3069 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n54 0 0.04fF $ **FLOATING
C3070 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n55 0 0.01fF $ **FLOATING
C3071 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n56 0 0.02fF $ **FLOATING
C3072 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n57 0 0.04fF $ **FLOATING
C3073 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t11 0 0.00fF $ **FLOATING
C3074 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.t10 0 0.01fF $ **FLOATING
C3075 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n58 0 0.02fF $ **FLOATING
C3076 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n59 0 0.03fF $ **FLOATING
C3077 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n60 0 0.01fF $ **FLOATING
C3078 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n61 0 0.02fF $ **FLOATING
C3079 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n62 0 0.04fF $ **FLOATING
C3080 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n63 0 0.01fF $ **FLOATING
C3081 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n64 0 0.02fF $ **FLOATING
C3082 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n65 0 0.04fF $ **FLOATING
C3083 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n66 0 0.04fF $ **FLOATING
C3084 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n67 0 0.04fF $ **FLOATING
C3085 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n68 0 0.04fF $ **FLOATING
C3086 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n69 0 0.04fF $ **FLOATING
C3087 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n70 0 0.04fF $ **FLOATING
C3088 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n71 0 0.04fF $ **FLOATING
C3089 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n72 0 0.07fF $ **FLOATING
C3090 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n73 0 0.01fF $ **FLOATING
C3091 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n74 0 0.02fF $ **FLOATING
C3092 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n75 0 0.04fF $ **FLOATING
C3093 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB.n76 0 0.01fF $ **FLOATING
C3094 sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0 0.07fF
C3095 sky130_fd_sc_hd__dfrbp_1_0[5]/D 0 0.22fF
C3096 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t8 0 0.01fF $ **FLOATING
C3097 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t5 0 0.01fF $ **FLOATING
C3098 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n0 0 0.03fF $ **FLOATING
C3099 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t0 0 0.01fF $ **FLOATING
C3100 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n1 0 0.01fF $ **FLOATING
C3101 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n2 0 0.03fF $ **FLOATING
C3102 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n3 0 0.01fF $ **FLOATING
C3103 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n4 0 0.03fF $ **FLOATING
C3104 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n5 0 0.01fF $ **FLOATING
C3105 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n6 0 0.03fF $ **FLOATING
C3106 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n7 0 0.01fF $ **FLOATING
C3107 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n8 0 0.02fF $ **FLOATING
C3108 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n9 0 0.04fF $ **FLOATING
C3109 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n10 0 0.01fF $ **FLOATING
C3110 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n11 0 0.03fF $ **FLOATING
C3111 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n12 0 0.01fF $ **FLOATING
C3112 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n13 0 0.03fF $ **FLOATING
C3113 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n14 0 0.01fF $ **FLOATING
C3114 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t4 0 0.01fF $ **FLOATING
C3115 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t1 0 0.00fF $ **FLOATING
C3116 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n15 0 0.06fF $ **FLOATING
C3117 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n16 0 0.01fF $ **FLOATING
C3118 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n17 0 0.03fF $ **FLOATING
C3119 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n18 0 0.02fF $ **FLOATING
C3120 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n19 0 0.06fF $ **FLOATING
C3121 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n20 0 0.12fF $ **FLOATING
C3122 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n21 0 0.01fF $ **FLOATING
C3123 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n22 0 0.03fF $ **FLOATING
C3124 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n23 0 0.04fF $ **FLOATING
C3125 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n24 0 0.01fF $ **FLOATING
C3126 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n25 0 0.02fF $ **FLOATING
C3127 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n26 0 0.04fF $ **FLOATING
C3128 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t2 0 0.01fF $ **FLOATING
C3129 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n27 0 0.03fF $ **FLOATING
C3130 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n28 0 0.03fF $ **FLOATING
C3131 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t6 0 0.01fF $ **FLOATING
C3132 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n29 0 0.02fF $ **FLOATING
C3133 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n30 0 0.03fF $ **FLOATING
C3134 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n31 0 0.01fF $ **FLOATING
C3135 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n32 0 0.02fF $ **FLOATING
C3136 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n33 0 0.04fF $ **FLOATING
C3137 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n34 0 0.01fF $ **FLOATING
C3138 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n35 0 0.02fF $ **FLOATING
C3139 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n36 0 0.04fF $ **FLOATING
C3140 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t7 0 0.00fF $ **FLOATING
C3141 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t3 0 0.01fF $ **FLOATING
C3142 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n37 0 0.02fF $ **FLOATING
C3143 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n38 0 0.02fF $ **FLOATING
C3144 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n39 0 0.01fF $ **FLOATING
C3145 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n40 0 0.02fF $ **FLOATING
C3146 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n41 0 0.04fF $ **FLOATING
C3147 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n42 0 0.01fF $ **FLOATING
C3148 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n43 0 0.03fF $ **FLOATING
C3149 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n44 0 0.04fF $ **FLOATING
C3150 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n45 0 0.01fF $ **FLOATING
C3151 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n46 0 0.03fF $ **FLOATING
C3152 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n47 0 0.04fF $ **FLOATING
C3153 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n48 0 0.01fF $ **FLOATING
C3154 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n49 0 0.03fF $ **FLOATING
C3155 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n50 0 0.04fF $ **FLOATING
C3156 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t9 0 0.03fF $ **FLOATING
C3157 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n51 0 0.05fF $ **FLOATING
C3158 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n52 0 0.01fF $ **FLOATING
C3159 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n53 0 0.02fF $ **FLOATING
C3160 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n54 0 0.04fF $ **FLOATING
C3161 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n55 0 0.01fF $ **FLOATING
C3162 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n56 0 0.02fF $ **FLOATING
C3163 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n57 0 0.04fF $ **FLOATING
C3164 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t11 0 0.00fF $ **FLOATING
C3165 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.t10 0 0.01fF $ **FLOATING
C3166 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n58 0 0.02fF $ **FLOATING
C3167 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n59 0 0.03fF $ **FLOATING
C3168 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n60 0 0.01fF $ **FLOATING
C3169 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n61 0 0.02fF $ **FLOATING
C3170 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n62 0 0.04fF $ **FLOATING
C3171 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n63 0 0.01fF $ **FLOATING
C3172 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n64 0 0.02fF $ **FLOATING
C3173 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n65 0 0.04fF $ **FLOATING
C3174 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n66 0 0.04fF $ **FLOATING
C3175 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n67 0 0.04fF $ **FLOATING
C3176 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n68 0 0.04fF $ **FLOATING
C3177 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n69 0 0.04fF $ **FLOATING
C3178 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n70 0 0.04fF $ **FLOATING
C3179 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n71 0 0.04fF $ **FLOATING
C3180 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n72 0 0.07fF $ **FLOATING
C3181 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n73 0 0.01fF $ **FLOATING
C3182 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n74 0 0.02fF $ **FLOATING
C3183 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n75 0 0.04fF $ **FLOATING
C3184 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB.n76 0 0.01fF $ **FLOATING
C3185 sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0 0.07fF
C3186 sky130_fd_sc_hd__dfrbp_1_0[4]/D 0 2.14fF
C3187 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t8 0 0.01fF $ **FLOATING
C3188 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t5 0 0.01fF $ **FLOATING
C3189 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n0 0 0.03fF $ **FLOATING
C3190 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t0 0 0.01fF $ **FLOATING
C3191 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n1 0 0.01fF $ **FLOATING
C3192 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n2 0 0.03fF $ **FLOATING
C3193 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n3 0 0.01fF $ **FLOATING
C3194 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n4 0 0.03fF $ **FLOATING
C3195 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n5 0 0.01fF $ **FLOATING
C3196 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n6 0 0.03fF $ **FLOATING
C3197 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n7 0 0.01fF $ **FLOATING
C3198 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n8 0 0.02fF $ **FLOATING
C3199 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n9 0 0.04fF $ **FLOATING
C3200 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n10 0 0.01fF $ **FLOATING
C3201 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n11 0 0.03fF $ **FLOATING
C3202 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n12 0 0.01fF $ **FLOATING
C3203 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n13 0 0.03fF $ **FLOATING
C3204 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n14 0 0.01fF $ **FLOATING
C3205 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t4 0 0.01fF $ **FLOATING
C3206 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t1 0 0.00fF $ **FLOATING
C3207 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n15 0 0.06fF $ **FLOATING
C3208 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n16 0 0.01fF $ **FLOATING
C3209 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n17 0 0.03fF $ **FLOATING
C3210 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n18 0 0.02fF $ **FLOATING
C3211 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n19 0 0.06fF $ **FLOATING
C3212 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n20 0 0.12fF $ **FLOATING
C3213 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n21 0 0.01fF $ **FLOATING
C3214 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n22 0 0.03fF $ **FLOATING
C3215 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n23 0 0.04fF $ **FLOATING
C3216 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n24 0 0.01fF $ **FLOATING
C3217 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n25 0 0.02fF $ **FLOATING
C3218 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n26 0 0.04fF $ **FLOATING
C3219 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t2 0 0.01fF $ **FLOATING
C3220 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n27 0 0.03fF $ **FLOATING
C3221 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n28 0 0.03fF $ **FLOATING
C3222 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t6 0 0.01fF $ **FLOATING
C3223 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n29 0 0.02fF $ **FLOATING
C3224 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n30 0 0.03fF $ **FLOATING
C3225 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n31 0 0.01fF $ **FLOATING
C3226 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n32 0 0.02fF $ **FLOATING
C3227 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n33 0 0.04fF $ **FLOATING
C3228 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n34 0 0.01fF $ **FLOATING
C3229 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n35 0 0.02fF $ **FLOATING
C3230 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n36 0 0.04fF $ **FLOATING
C3231 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t7 0 0.00fF $ **FLOATING
C3232 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t3 0 0.01fF $ **FLOATING
C3233 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n37 0 0.02fF $ **FLOATING
C3234 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n38 0 0.02fF $ **FLOATING
C3235 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n39 0 0.01fF $ **FLOATING
C3236 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n40 0 0.02fF $ **FLOATING
C3237 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n41 0 0.04fF $ **FLOATING
C3238 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n42 0 0.01fF $ **FLOATING
C3239 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n43 0 0.03fF $ **FLOATING
C3240 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n44 0 0.04fF $ **FLOATING
C3241 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n45 0 0.01fF $ **FLOATING
C3242 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n46 0 0.03fF $ **FLOATING
C3243 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n47 0 0.04fF $ **FLOATING
C3244 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n48 0 0.01fF $ **FLOATING
C3245 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n49 0 0.03fF $ **FLOATING
C3246 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n50 0 0.04fF $ **FLOATING
C3247 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t9 0 0.03fF $ **FLOATING
C3248 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n51 0 0.05fF $ **FLOATING
C3249 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n52 0 0.01fF $ **FLOATING
C3250 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n53 0 0.02fF $ **FLOATING
C3251 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n54 0 0.04fF $ **FLOATING
C3252 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n55 0 0.01fF $ **FLOATING
C3253 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n56 0 0.02fF $ **FLOATING
C3254 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n57 0 0.04fF $ **FLOATING
C3255 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t11 0 0.00fF $ **FLOATING
C3256 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.t10 0 0.01fF $ **FLOATING
C3257 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n58 0 0.02fF $ **FLOATING
C3258 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n59 0 0.03fF $ **FLOATING
C3259 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n60 0 0.01fF $ **FLOATING
C3260 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n61 0 0.02fF $ **FLOATING
C3261 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n62 0 0.04fF $ **FLOATING
C3262 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n63 0 0.01fF $ **FLOATING
C3263 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n64 0 0.02fF $ **FLOATING
C3264 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n65 0 0.04fF $ **FLOATING
C3265 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n66 0 0.04fF $ **FLOATING
C3266 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n67 0 0.04fF $ **FLOATING
C3267 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n68 0 0.04fF $ **FLOATING
C3268 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n69 0 0.04fF $ **FLOATING
C3269 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n70 0 0.04fF $ **FLOATING
C3270 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n71 0 0.04fF $ **FLOATING
C3271 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n72 0 0.07fF $ **FLOATING
C3272 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n73 0 0.01fF $ **FLOATING
C3273 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n74 0 0.02fF $ **FLOATING
C3274 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n75 0 0.04fF $ **FLOATING
C3275 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB.n76 0 0.01fF $ **FLOATING
C3276 sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0 0.07fF
C3277 sky130_fd_sc_hd__dfrbp_1_0[3]/D 0 0.28fF
C3278 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t0 0 0.05fF
C3279 sky130_fd_sc_hd__dfrbp_1_0[4]/D.t1 0 0.06fF
C3280 sky130_fd_sc_hd__dfrbp_1_0[4]/D.n0 0 0.07fF $ **FLOATING
C3281 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t8 0 0.01fF $ **FLOATING
C3282 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t5 0 0.01fF $ **FLOATING
C3283 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n0 0 0.03fF $ **FLOATING
C3284 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t0 0 0.01fF $ **FLOATING
C3285 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n1 0 0.01fF $ **FLOATING
C3286 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n2 0 0.03fF $ **FLOATING
C3287 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n3 0 0.01fF $ **FLOATING
C3288 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n4 0 0.03fF $ **FLOATING
C3289 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n5 0 0.01fF $ **FLOATING
C3290 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n6 0 0.03fF $ **FLOATING
C3291 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n7 0 0.01fF $ **FLOATING
C3292 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n8 0 0.02fF $ **FLOATING
C3293 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n9 0 0.04fF $ **FLOATING
C3294 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n10 0 0.01fF $ **FLOATING
C3295 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n11 0 0.03fF $ **FLOATING
C3296 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n12 0 0.01fF $ **FLOATING
C3297 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n13 0 0.03fF $ **FLOATING
C3298 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n14 0 0.01fF $ **FLOATING
C3299 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t4 0 0.01fF $ **FLOATING
C3300 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t1 0 0.00fF $ **FLOATING
C3301 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n15 0 0.06fF $ **FLOATING
C3302 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n16 0 0.01fF $ **FLOATING
C3303 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n17 0 0.03fF $ **FLOATING
C3304 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n18 0 0.02fF $ **FLOATING
C3305 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n19 0 0.06fF $ **FLOATING
C3306 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n20 0 0.12fF $ **FLOATING
C3307 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n21 0 0.01fF $ **FLOATING
C3308 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n22 0 0.03fF $ **FLOATING
C3309 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n23 0 0.04fF $ **FLOATING
C3310 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n24 0 0.01fF $ **FLOATING
C3311 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n25 0 0.02fF $ **FLOATING
C3312 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n26 0 0.04fF $ **FLOATING
C3313 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t2 0 0.01fF $ **FLOATING
C3314 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n27 0 0.03fF $ **FLOATING
C3315 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n28 0 0.03fF $ **FLOATING
C3316 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t6 0 0.01fF $ **FLOATING
C3317 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n29 0 0.02fF $ **FLOATING
C3318 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n30 0 0.03fF $ **FLOATING
C3319 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n31 0 0.01fF $ **FLOATING
C3320 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n32 0 0.02fF $ **FLOATING
C3321 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n33 0 0.04fF $ **FLOATING
C3322 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n34 0 0.01fF $ **FLOATING
C3323 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n35 0 0.02fF $ **FLOATING
C3324 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n36 0 0.04fF $ **FLOATING
C3325 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t7 0 0.00fF $ **FLOATING
C3326 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t3 0 0.01fF $ **FLOATING
C3327 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n37 0 0.02fF $ **FLOATING
C3328 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n38 0 0.02fF $ **FLOATING
C3329 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n39 0 0.01fF $ **FLOATING
C3330 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n40 0 0.02fF $ **FLOATING
C3331 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n41 0 0.04fF $ **FLOATING
C3332 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n42 0 0.01fF $ **FLOATING
C3333 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n43 0 0.03fF $ **FLOATING
C3334 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n44 0 0.04fF $ **FLOATING
C3335 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n45 0 0.01fF $ **FLOATING
C3336 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n46 0 0.03fF $ **FLOATING
C3337 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n47 0 0.04fF $ **FLOATING
C3338 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n48 0 0.01fF $ **FLOATING
C3339 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n49 0 0.03fF $ **FLOATING
C3340 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n50 0 0.04fF $ **FLOATING
C3341 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t9 0 0.03fF $ **FLOATING
C3342 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n51 0 0.05fF $ **FLOATING
C3343 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n52 0 0.01fF $ **FLOATING
C3344 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n53 0 0.02fF $ **FLOATING
C3345 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n54 0 0.04fF $ **FLOATING
C3346 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n55 0 0.01fF $ **FLOATING
C3347 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n56 0 0.02fF $ **FLOATING
C3348 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n57 0 0.04fF $ **FLOATING
C3349 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t11 0 0.00fF $ **FLOATING
C3350 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.t10 0 0.01fF $ **FLOATING
C3351 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n58 0 0.02fF $ **FLOATING
C3352 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n59 0 0.03fF $ **FLOATING
C3353 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n60 0 0.01fF $ **FLOATING
C3354 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n61 0 0.02fF $ **FLOATING
C3355 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n62 0 0.04fF $ **FLOATING
C3356 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n63 0 0.01fF $ **FLOATING
C3357 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n64 0 0.02fF $ **FLOATING
C3358 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n65 0 0.04fF $ **FLOATING
C3359 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n66 0 0.04fF $ **FLOATING
C3360 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n67 0 0.04fF $ **FLOATING
C3361 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n68 0 0.04fF $ **FLOATING
C3362 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n69 0 0.04fF $ **FLOATING
C3363 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n70 0 0.04fF $ **FLOATING
C3364 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n71 0 0.04fF $ **FLOATING
C3365 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n72 0 0.07fF $ **FLOATING
C3366 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n73 0 0.01fF $ **FLOATING
C3367 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n74 0 0.02fF $ **FLOATING
C3368 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n75 0 0.04fF $ **FLOATING
C3369 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB.n76 0 0.01fF $ **FLOATING
C3370 sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0 0.07fF
C3371 sky130_fd_sc_hd__dfrbp_1_0[2]/D 0 1.77fF
C3372 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t8 0 0.01fF $ **FLOATING
C3373 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t5 0 0.01fF $ **FLOATING
C3374 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n0 0 0.03fF $ **FLOATING
C3375 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t0 0 0.01fF $ **FLOATING
C3376 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n1 0 0.01fF $ **FLOATING
C3377 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n2 0 0.03fF $ **FLOATING
C3378 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n3 0 0.01fF $ **FLOATING
C3379 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n4 0 0.03fF $ **FLOATING
C3380 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n5 0 0.01fF $ **FLOATING
C3381 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n6 0 0.03fF $ **FLOATING
C3382 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n7 0 0.01fF $ **FLOATING
C3383 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n8 0 0.02fF $ **FLOATING
C3384 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n9 0 0.04fF $ **FLOATING
C3385 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n10 0 0.01fF $ **FLOATING
C3386 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n11 0 0.03fF $ **FLOATING
C3387 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n12 0 0.01fF $ **FLOATING
C3388 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n13 0 0.03fF $ **FLOATING
C3389 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n14 0 0.01fF $ **FLOATING
C3390 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t4 0 0.01fF $ **FLOATING
C3391 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t1 0 0.00fF $ **FLOATING
C3392 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n15 0 0.06fF $ **FLOATING
C3393 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n16 0 0.01fF $ **FLOATING
C3394 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n17 0 0.03fF $ **FLOATING
C3395 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n18 0 0.02fF $ **FLOATING
C3396 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n19 0 0.06fF $ **FLOATING
C3397 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n20 0 0.12fF $ **FLOATING
C3398 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n21 0 0.01fF $ **FLOATING
C3399 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n22 0 0.03fF $ **FLOATING
C3400 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n23 0 0.04fF $ **FLOATING
C3401 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n24 0 0.01fF $ **FLOATING
C3402 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n25 0 0.02fF $ **FLOATING
C3403 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n26 0 0.04fF $ **FLOATING
C3404 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t2 0 0.01fF $ **FLOATING
C3405 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n27 0 0.03fF $ **FLOATING
C3406 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n28 0 0.03fF $ **FLOATING
C3407 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t6 0 0.01fF $ **FLOATING
C3408 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n29 0 0.02fF $ **FLOATING
C3409 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n30 0 0.03fF $ **FLOATING
C3410 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n31 0 0.01fF $ **FLOATING
C3411 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n32 0 0.02fF $ **FLOATING
C3412 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n33 0 0.04fF $ **FLOATING
C3413 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n34 0 0.01fF $ **FLOATING
C3414 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n35 0 0.02fF $ **FLOATING
C3415 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n36 0 0.04fF $ **FLOATING
C3416 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t7 0 0.00fF $ **FLOATING
C3417 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t3 0 0.01fF $ **FLOATING
C3418 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n37 0 0.02fF $ **FLOATING
C3419 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n38 0 0.02fF $ **FLOATING
C3420 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n39 0 0.01fF $ **FLOATING
C3421 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n40 0 0.02fF $ **FLOATING
C3422 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n41 0 0.04fF $ **FLOATING
C3423 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n42 0 0.01fF $ **FLOATING
C3424 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n43 0 0.03fF $ **FLOATING
C3425 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n44 0 0.04fF $ **FLOATING
C3426 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n45 0 0.01fF $ **FLOATING
C3427 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n46 0 0.03fF $ **FLOATING
C3428 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n47 0 0.04fF $ **FLOATING
C3429 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n48 0 0.01fF $ **FLOATING
C3430 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n49 0 0.03fF $ **FLOATING
C3431 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n50 0 0.04fF $ **FLOATING
C3432 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t9 0 0.03fF $ **FLOATING
C3433 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n51 0 0.05fF $ **FLOATING
C3434 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n52 0 0.01fF $ **FLOATING
C3435 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n53 0 0.02fF $ **FLOATING
C3436 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n54 0 0.04fF $ **FLOATING
C3437 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n55 0 0.01fF $ **FLOATING
C3438 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n56 0 0.02fF $ **FLOATING
C3439 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n57 0 0.04fF $ **FLOATING
C3440 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t11 0 0.00fF $ **FLOATING
C3441 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.t10 0 0.01fF $ **FLOATING
C3442 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n58 0 0.02fF $ **FLOATING
C3443 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n59 0 0.03fF $ **FLOATING
C3444 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n60 0 0.01fF $ **FLOATING
C3445 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n61 0 0.02fF $ **FLOATING
C3446 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n62 0 0.04fF $ **FLOATING
C3447 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n63 0 0.01fF $ **FLOATING
C3448 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n64 0 0.02fF $ **FLOATING
C3449 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n65 0 0.04fF $ **FLOATING
C3450 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n66 0 0.04fF $ **FLOATING
C3451 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n67 0 0.04fF $ **FLOATING
C3452 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n68 0 0.04fF $ **FLOATING
C3453 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n69 0 0.04fF $ **FLOATING
C3454 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n70 0 0.04fF $ **FLOATING
C3455 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n71 0 0.04fF $ **FLOATING
C3456 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n72 0 0.07fF $ **FLOATING
C3457 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n73 0 0.01fF $ **FLOATING
C3458 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n74 0 0.02fF $ **FLOATING
C3459 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n75 0 0.04fF $ **FLOATING
C3460 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB.n76 0 0.01fF $ **FLOATING
C3461 sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0 0.07fF
C3462 sky130_fd_sc_hd__dfrbp_1_0[1]/D 0 0.76fF
C3463 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t8 0 0.01fF $ **FLOATING
C3464 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t5 0 0.01fF $ **FLOATING
C3465 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n0 0 0.03fF $ **FLOATING
C3466 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t0 0 0.01fF $ **FLOATING
C3467 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n1 0 0.01fF $ **FLOATING
C3468 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n2 0 0.03fF $ **FLOATING
C3469 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n3 0 0.01fF $ **FLOATING
C3470 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n4 0 0.03fF $ **FLOATING
C3471 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n5 0 0.01fF $ **FLOATING
C3472 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n6 0 0.03fF $ **FLOATING
C3473 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n7 0 0.01fF $ **FLOATING
C3474 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n8 0 0.02fF $ **FLOATING
C3475 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n9 0 0.04fF $ **FLOATING
C3476 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n10 0 0.01fF $ **FLOATING
C3477 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n11 0 0.03fF $ **FLOATING
C3478 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n12 0 0.01fF $ **FLOATING
C3479 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n13 0 0.03fF $ **FLOATING
C3480 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n14 0 0.01fF $ **FLOATING
C3481 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t4 0 0.01fF $ **FLOATING
C3482 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t1 0 0.00fF $ **FLOATING
C3483 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n15 0 0.06fF $ **FLOATING
C3484 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n16 0 0.01fF $ **FLOATING
C3485 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n17 0 0.03fF $ **FLOATING
C3486 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n18 0 0.02fF $ **FLOATING
C3487 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n19 0 0.06fF $ **FLOATING
C3488 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n20 0 0.12fF $ **FLOATING
C3489 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n21 0 0.01fF $ **FLOATING
C3490 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n22 0 0.03fF $ **FLOATING
C3491 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n23 0 0.04fF $ **FLOATING
C3492 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n24 0 0.01fF $ **FLOATING
C3493 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n25 0 0.02fF $ **FLOATING
C3494 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n26 0 0.04fF $ **FLOATING
C3495 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t2 0 0.01fF $ **FLOATING
C3496 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n27 0 0.03fF $ **FLOATING
C3497 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n28 0 0.03fF $ **FLOATING
C3498 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t6 0 0.01fF $ **FLOATING
C3499 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n29 0 0.02fF $ **FLOATING
C3500 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n30 0 0.03fF $ **FLOATING
C3501 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n31 0 0.01fF $ **FLOATING
C3502 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n32 0 0.02fF $ **FLOATING
C3503 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n33 0 0.04fF $ **FLOATING
C3504 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n34 0 0.01fF $ **FLOATING
C3505 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n35 0 0.02fF $ **FLOATING
C3506 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n36 0 0.04fF $ **FLOATING
C3507 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t7 0 0.00fF $ **FLOATING
C3508 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t3 0 0.01fF $ **FLOATING
C3509 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n37 0 0.02fF $ **FLOATING
C3510 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n38 0 0.02fF $ **FLOATING
C3511 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n39 0 0.01fF $ **FLOATING
C3512 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n40 0 0.02fF $ **FLOATING
C3513 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n41 0 0.04fF $ **FLOATING
C3514 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n42 0 0.01fF $ **FLOATING
C3515 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n43 0 0.03fF $ **FLOATING
C3516 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n44 0 0.04fF $ **FLOATING
C3517 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n45 0 0.01fF $ **FLOATING
C3518 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n46 0 0.03fF $ **FLOATING
C3519 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n47 0 0.04fF $ **FLOATING
C3520 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n48 0 0.01fF $ **FLOATING
C3521 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n49 0 0.03fF $ **FLOATING
C3522 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n50 0 0.04fF $ **FLOATING
C3523 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t9 0 0.03fF $ **FLOATING
C3524 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n51 0 0.05fF $ **FLOATING
C3525 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n52 0 0.01fF $ **FLOATING
C3526 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n53 0 0.02fF $ **FLOATING
C3527 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n54 0 0.04fF $ **FLOATING
C3528 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n55 0 0.01fF $ **FLOATING
C3529 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n56 0 0.02fF $ **FLOATING
C3530 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n57 0 0.04fF $ **FLOATING
C3531 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t11 0 0.00fF $ **FLOATING
C3532 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.t10 0 0.01fF $ **FLOATING
C3533 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n58 0 0.02fF $ **FLOATING
C3534 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n59 0 0.03fF $ **FLOATING
C3535 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n60 0 0.01fF $ **FLOATING
C3536 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n61 0 0.02fF $ **FLOATING
C3537 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n62 0 0.04fF $ **FLOATING
C3538 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n63 0 0.01fF $ **FLOATING
C3539 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n64 0 0.02fF $ **FLOATING
C3540 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n65 0 0.04fF $ **FLOATING
C3541 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n66 0 0.04fF $ **FLOATING
C3542 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n67 0 0.04fF $ **FLOATING
C3543 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n68 0 0.04fF $ **FLOATING
C3544 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n69 0 0.04fF $ **FLOATING
C3545 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n70 0 0.04fF $ **FLOATING
C3546 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n71 0 0.04fF $ **FLOATING
C3547 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n72 0 0.07fF $ **FLOATING
C3548 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n73 0 0.01fF $ **FLOATING
C3549 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n74 0 0.02fF $ **FLOATING
C3550 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n75 0 0.04fF $ **FLOATING
C3551 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB.n76 0 0.01fF $ **FLOATING
C3552 sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0 0.07fF
C3553 sky130_fd_sc_hd__dfrbp_1_0[0]/D 0 2.23fF
C3554 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t8 0 0.01fF $ **FLOATING
C3555 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t5 0 0.01fF $ **FLOATING
C3556 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n0 0 0.03fF $ **FLOATING
C3557 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t0 0 0.01fF $ **FLOATING
C3558 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n1 0 0.01fF $ **FLOATING
C3559 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n2 0 0.03fF $ **FLOATING
C3560 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n3 0 0.01fF $ **FLOATING
C3561 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n4 0 0.03fF $ **FLOATING
C3562 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n5 0 0.01fF $ **FLOATING
C3563 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n6 0 0.03fF $ **FLOATING
C3564 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n7 0 0.01fF $ **FLOATING
C3565 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n8 0 0.02fF $ **FLOATING
C3566 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n9 0 0.04fF $ **FLOATING
C3567 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n10 0 0.01fF $ **FLOATING
C3568 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n11 0 0.03fF $ **FLOATING
C3569 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n12 0 0.01fF $ **FLOATING
C3570 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n13 0 0.03fF $ **FLOATING
C3571 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n14 0 0.01fF $ **FLOATING
C3572 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t4 0 0.01fF $ **FLOATING
C3573 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t1 0 0.00fF $ **FLOATING
C3574 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n15 0 0.06fF $ **FLOATING
C3575 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n16 0 0.01fF $ **FLOATING
C3576 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n17 0 0.03fF $ **FLOATING
C3577 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n18 0 0.02fF $ **FLOATING
C3578 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n19 0 0.06fF $ **FLOATING
C3579 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n20 0 0.12fF $ **FLOATING
C3580 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n21 0 0.01fF $ **FLOATING
C3581 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n22 0 0.03fF $ **FLOATING
C3582 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n23 0 0.04fF $ **FLOATING
C3583 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n24 0 0.01fF $ **FLOATING
C3584 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n25 0 0.02fF $ **FLOATING
C3585 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n26 0 0.04fF $ **FLOATING
C3586 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t2 0 0.01fF $ **FLOATING
C3587 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n27 0 0.03fF $ **FLOATING
C3588 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n28 0 0.03fF $ **FLOATING
C3589 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t6 0 0.01fF $ **FLOATING
C3590 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n29 0 0.02fF $ **FLOATING
C3591 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n30 0 0.03fF $ **FLOATING
C3592 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n31 0 0.01fF $ **FLOATING
C3593 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n32 0 0.02fF $ **FLOATING
C3594 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n33 0 0.04fF $ **FLOATING
C3595 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n34 0 0.01fF $ **FLOATING
C3596 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n35 0 0.02fF $ **FLOATING
C3597 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n36 0 0.04fF $ **FLOATING
C3598 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t7 0 0.00fF $ **FLOATING
C3599 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t3 0 0.01fF $ **FLOATING
C3600 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n37 0 0.02fF $ **FLOATING
C3601 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n38 0 0.02fF $ **FLOATING
C3602 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n39 0 0.01fF $ **FLOATING
C3603 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n40 0 0.02fF $ **FLOATING
C3604 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n41 0 0.04fF $ **FLOATING
C3605 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n42 0 0.01fF $ **FLOATING
C3606 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n43 0 0.03fF $ **FLOATING
C3607 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n44 0 0.04fF $ **FLOATING
C3608 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n45 0 0.01fF $ **FLOATING
C3609 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n46 0 0.03fF $ **FLOATING
C3610 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n47 0 0.04fF $ **FLOATING
C3611 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n48 0 0.01fF $ **FLOATING
C3612 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n49 0 0.03fF $ **FLOATING
C3613 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n50 0 0.04fF $ **FLOATING
C3614 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t9 0 0.03fF $ **FLOATING
C3615 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n51 0 0.05fF $ **FLOATING
C3616 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n52 0 0.01fF $ **FLOATING
C3617 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n53 0 0.02fF $ **FLOATING
C3618 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n54 0 0.04fF $ **FLOATING
C3619 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n55 0 0.01fF $ **FLOATING
C3620 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n56 0 0.02fF $ **FLOATING
C3621 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n57 0 0.04fF $ **FLOATING
C3622 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t11 0 0.00fF $ **FLOATING
C3623 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.t10 0 0.01fF $ **FLOATING
C3624 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n58 0 0.02fF $ **FLOATING
C3625 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n59 0 0.03fF $ **FLOATING
C3626 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n60 0 0.01fF $ **FLOATING
C3627 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n61 0 0.02fF $ **FLOATING
C3628 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n62 0 0.04fF $ **FLOATING
C3629 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n63 0 0.01fF $ **FLOATING
C3630 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n64 0 0.02fF $ **FLOATING
C3631 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n65 0 0.04fF $ **FLOATING
C3632 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n66 0 0.04fF $ **FLOATING
C3633 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n67 0 0.04fF $ **FLOATING
C3634 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n68 0 0.04fF $ **FLOATING
C3635 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n69 0 0.04fF $ **FLOATING
C3636 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n70 0 0.04fF $ **FLOATING
C3637 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n71 0 0.04fF $ **FLOATING
C3638 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n72 0 0.07fF $ **FLOATING
C3639 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n73 0 0.01fF $ **FLOATING
C3640 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n74 0 0.02fF $ **FLOATING
C3641 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n75 0 0.04fF $ **FLOATING
C3642 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB.n76 0 0.01fF $ **FLOATING
C3643 sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0 0.07fF
C3644 Vclk 0 0.33fF
C3645 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t0 0 0.05fF
C3646 sky130_fd_sc_hd__dfrbp_1_0[0]/D.t1 0 0.06fF
C3647 sky130_fd_sc_hd__dfrbp_1_0[0]/D.n0 0 0.07fF $ **FLOATING
C3648 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t8 0 0.01fF $ **FLOATING
C3649 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t5 0 0.01fF $ **FLOATING
C3650 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n0 0 0.03fF $ **FLOATING
C3651 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t0 0 0.01fF $ **FLOATING
C3652 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n1 0 0.01fF $ **FLOATING
C3653 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n2 0 0.03fF $ **FLOATING
C3654 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n3 0 0.01fF $ **FLOATING
C3655 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n4 0 0.03fF $ **FLOATING
C3656 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n5 0 0.01fF $ **FLOATING
C3657 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n6 0 0.03fF $ **FLOATING
C3658 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n7 0 0.01fF $ **FLOATING
C3659 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n8 0 0.02fF $ **FLOATING
C3660 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n9 0 0.04fF $ **FLOATING
C3661 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n10 0 0.01fF $ **FLOATING
C3662 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n11 0 0.03fF $ **FLOATING
C3663 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n12 0 0.01fF $ **FLOATING
C3664 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n13 0 0.03fF $ **FLOATING
C3665 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n14 0 0.01fF $ **FLOATING
C3666 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t4 0 0.01fF $ **FLOATING
C3667 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t1 0 0.00fF $ **FLOATING
C3668 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n15 0 0.06fF $ **FLOATING
C3669 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n16 0 0.01fF $ **FLOATING
C3670 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n17 0 0.03fF $ **FLOATING
C3671 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n18 0 0.02fF $ **FLOATING
C3672 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n19 0 0.06fF $ **FLOATING
C3673 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n20 0 0.12fF $ **FLOATING
C3674 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n21 0 0.01fF $ **FLOATING
C3675 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n22 0 0.03fF $ **FLOATING
C3676 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n23 0 0.04fF $ **FLOATING
C3677 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n24 0 0.01fF $ **FLOATING
C3678 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n25 0 0.02fF $ **FLOATING
C3679 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n26 0 0.04fF $ **FLOATING
C3680 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t2 0 0.01fF $ **FLOATING
C3681 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n27 0 0.03fF $ **FLOATING
C3682 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n28 0 0.03fF $ **FLOATING
C3683 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t6 0 0.01fF $ **FLOATING
C3684 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n29 0 0.02fF $ **FLOATING
C3685 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n30 0 0.03fF $ **FLOATING
C3686 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n31 0 0.01fF $ **FLOATING
C3687 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n32 0 0.02fF $ **FLOATING
C3688 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n33 0 0.04fF $ **FLOATING
C3689 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n34 0 0.01fF $ **FLOATING
C3690 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n35 0 0.02fF $ **FLOATING
C3691 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n36 0 0.04fF $ **FLOATING
C3692 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t7 0 0.00fF $ **FLOATING
C3693 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t3 0 0.01fF $ **FLOATING
C3694 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n37 0 0.02fF $ **FLOATING
C3695 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n38 0 0.02fF $ **FLOATING
C3696 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n39 0 0.01fF $ **FLOATING
C3697 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n40 0 0.02fF $ **FLOATING
C3698 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n41 0 0.04fF $ **FLOATING
C3699 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n42 0 0.01fF $ **FLOATING
C3700 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n43 0 0.03fF $ **FLOATING
C3701 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n44 0 0.04fF $ **FLOATING
C3702 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n45 0 0.01fF $ **FLOATING
C3703 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n46 0 0.03fF $ **FLOATING
C3704 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n47 0 0.04fF $ **FLOATING
C3705 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n48 0 0.01fF $ **FLOATING
C3706 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n49 0 0.03fF $ **FLOATING
C3707 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n50 0 0.04fF $ **FLOATING
C3708 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t9 0 0.03fF $ **FLOATING
C3709 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n51 0 0.05fF $ **FLOATING
C3710 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n52 0 0.01fF $ **FLOATING
C3711 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n53 0 0.02fF $ **FLOATING
C3712 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n54 0 0.04fF $ **FLOATING
C3713 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n55 0 0.01fF $ **FLOATING
C3714 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n56 0 0.02fF $ **FLOATING
C3715 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n57 0 0.04fF $ **FLOATING
C3716 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t11 0 0.00fF $ **FLOATING
C3717 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.t10 0 0.01fF $ **FLOATING
C3718 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n58 0 0.02fF $ **FLOATING
C3719 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n59 0 0.03fF $ **FLOATING
C3720 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n60 0 0.01fF $ **FLOATING
C3721 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n61 0 0.02fF $ **FLOATING
C3722 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n62 0 0.04fF $ **FLOATING
C3723 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n63 0 0.01fF $ **FLOATING
C3724 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n64 0 0.02fF $ **FLOATING
C3725 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n65 0 0.04fF $ **FLOATING
C3726 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n66 0 0.04fF $ **FLOATING
C3727 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n67 0 0.04fF $ **FLOATING
C3728 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n68 0 0.04fF $ **FLOATING
C3729 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n69 0 0.04fF $ **FLOATING
C3730 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n70 0 0.04fF $ **FLOATING
C3731 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n71 0 0.04fF $ **FLOATING
C3732 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n72 0 0.07fF $ **FLOATING
C3733 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n73 0 0.01fF $ **FLOATING
C3734 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n74 0 0.02fF $ **FLOATING
C3735 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n75 0 0.04fF $ **FLOATING
C3736 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB.n76 0 0.01fF $ **FLOATING
