* SPICE3 file created from extract.ext - technology: sky130A

X0 net2 GND GND sky130_fd_pr__res_xhigh_po_0p35 l=1.75e+09u
X1 net1 clkb_in net2 GND sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X2 net2 clk_in net1 VDD sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X3 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X4 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X5 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X6 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X7 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X8 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X9 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X10 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X11 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X12 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X13 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X14 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X15 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X16 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X17 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X18 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X19 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X20 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X21 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X22 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X23 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X24 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X25 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X26 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X27 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X28 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X29 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X30 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X31 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X32 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X33 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X34 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X35 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X36 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X37 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X38 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X39 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X40 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X41 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X42 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X43 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X44 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X45 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X46 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X47 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X48 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X49 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X50 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X51 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X52 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X53 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X54 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X55 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X56 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X57 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X58 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X59 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X60 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X61 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X62 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X63 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X64 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X65 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X66 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X67 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X68 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X69 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X70 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X71 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X72 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X73 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X74 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X75 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X76 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X77 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X78 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X79 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X80 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X81 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X82 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X83 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X84 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X85 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X86 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X87 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X88 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X89 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X90 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X91 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X92 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X93 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X94 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X95 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X96 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X97 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X98 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X99 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X100 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X101 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X102 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X103 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X104 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X105 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X106 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X107 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X108 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X109 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X110 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X111 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X112 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X113 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X114 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X115 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X116 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X117 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X118 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X119 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X120 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X121 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X122 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X123 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X124 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X125 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X126 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X127 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X128 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X129 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X130 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X131 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X132 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X133 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X134 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X135 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X136 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X137 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X138 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X139 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X140 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X141 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X142 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X143 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X144 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X145 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X146 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X147 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X148 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X149 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X150 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X151 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X152 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X153 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X154 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X155 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X156 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X157 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X158 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X159 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X160 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X161 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X162 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X163 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X164 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X165 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X166 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X167 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X168 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X169 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X170 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X171 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X172 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X173 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X174 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X175 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X176 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X177 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X178 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X179 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X180 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X181 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X182 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X183 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X184 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X185 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X186 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X187 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X188 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X189 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X190 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X191 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X192 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X193 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X194 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X195 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X196 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X197 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X198 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X199 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X200 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X201 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u
X202 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8 ad=1.06575e+12p pd=7.6545e+06u as=1.06575e+12p ps=7.6545e+06u w=7e+06u l=8e+06u

