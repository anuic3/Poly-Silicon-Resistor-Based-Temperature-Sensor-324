magic
tech sky130A
magscale 1 2
timestamp 1634815074
<< nwell >>
rect -6792 3168 11240 4900
rect -6792 3164 2184 3168
rect 2486 3164 11240 3168
rect 5476 3058 8626 3164
rect 9288 2992 10388 3164
<< nmos >>
rect -6492 2846 -6462 3046
rect -6276 2848 -6246 3048
rect -6058 2848 -6028 3048
rect -5836 2846 -5806 3046
rect -1306 2864 -1276 3064
rect -1090 2866 -1060 3066
rect -872 2866 -842 3066
rect -650 2864 -620 3064
rect 3870 2876 3900 3076
rect 4086 2878 4116 3078
rect 4304 2878 4334 3078
rect 4526 2876 4556 3076
rect 9526 2668 9556 2868
rect 9742 2670 9772 2870
rect 9960 2670 9990 2870
rect 10182 2668 10212 2868
<< pmos >>
rect -6516 3284 -6486 3684
rect -6284 3282 -6254 3682
rect -6056 3280 -6026 3680
rect -5838 3282 -5808 3682
rect -1330 3302 -1300 3702
rect -1098 3300 -1068 3700
rect -870 3298 -840 3698
rect -652 3300 -622 3700
rect 3846 3314 3876 3714
rect 4078 3312 4108 3712
rect 4306 3310 4336 3710
rect 4524 3312 4554 3712
rect 9502 3106 9532 3506
rect 9734 3104 9764 3504
rect 9962 3102 9992 3502
rect 10180 3104 10210 3504
<< pmoslvt >>
rect -4970 3562 -4770 4562
rect -4314 3570 -4114 4570
rect -4056 3570 -3856 4570
rect -3314 3570 -3114 4570
rect -3056 3570 -2856 4570
rect -2408 3574 -2208 4574
rect 966 3302 1166 4302
rect 1445 3294 1645 4294
rect 1703 3294 1903 4294
rect 2103 3296 2303 4296
rect 2361 3296 2561 4296
rect 2760 3276 2960 4276
rect 6240 3174 6440 4174
rect 6634 3156 7034 4156
rect 7206 3156 7606 4156
rect 7828 3186 8028 4186
<< nmoslvt >>
rect 1196 1930 1396 2330
rect 1454 1930 1654 2330
rect 1712 1930 1912 2330
rect 2210 1930 2410 2330
rect 2468 1930 2668 2330
rect 2726 1930 2926 2330
rect 1196 1374 1396 1774
rect 1454 1374 1654 1774
rect 1712 1374 1912 1774
rect 2210 1374 2410 1774
rect 2468 1374 2668 1774
rect 2726 1374 2926 1774
rect -4964 978 -4764 1178
rect -4488 980 -3688 1180
rect -3516 980 -2716 1180
rect -2430 978 -2230 1178
rect 1517 330 1917 530
rect 2112 330 2512 530
rect 5728 -1040 5928 1760
rect 6278 826 6478 1626
rect 6536 826 6736 1626
rect 6794 826 6994 1626
rect 7278 826 7478 1626
rect 7536 826 7736 1626
rect 7794 826 7994 1626
rect 6278 -130 6478 670
rect 6536 -130 6736 670
rect 6794 -130 6994 670
rect 7278 -130 7478 670
rect 7536 -130 7736 670
rect 7794 -130 7994 670
rect 6278 -1086 6478 -286
rect 6536 -1086 6736 -286
rect 6794 -1086 6994 -286
rect 7278 -1086 7478 -286
rect 7536 -1086 7736 -286
rect 7794 -1086 7994 -286
rect 8326 -1090 8526 1710
<< ndiff >>
rect -6550 2990 -6492 3046
rect -6550 2902 -6538 2990
rect -6504 2902 -6492 2990
rect -6550 2846 -6492 2902
rect -6462 2990 -6404 3046
rect -6462 2902 -6450 2990
rect -6416 2902 -6404 2990
rect -6462 2846 -6404 2902
rect -6334 2992 -6276 3048
rect -6334 2904 -6322 2992
rect -6288 2904 -6276 2992
rect -6334 2848 -6276 2904
rect -6246 2992 -6188 3048
rect -6246 2904 -6234 2992
rect -6200 2904 -6188 2992
rect -6246 2848 -6188 2904
rect -6116 2992 -6058 3048
rect -6116 2904 -6104 2992
rect -6070 2904 -6058 2992
rect -6116 2848 -6058 2904
rect -6028 2992 -5970 3048
rect -6028 2904 -6016 2992
rect -5982 2904 -5970 2992
rect -6028 2848 -5970 2904
rect -5894 2990 -5836 3046
rect -5894 2902 -5882 2990
rect -5848 2902 -5836 2990
rect -5894 2846 -5836 2902
rect -5806 2990 -5748 3046
rect -5806 2902 -5794 2990
rect -5760 2902 -5748 2990
rect -5806 2846 -5748 2902
rect -1364 3008 -1306 3064
rect -1364 2920 -1352 3008
rect -1318 2920 -1306 3008
rect -1364 2864 -1306 2920
rect -1276 3008 -1218 3064
rect -1276 2920 -1264 3008
rect -1230 2920 -1218 3008
rect -1276 2864 -1218 2920
rect -1148 3010 -1090 3066
rect -1148 2922 -1136 3010
rect -1102 2922 -1090 3010
rect -1148 2866 -1090 2922
rect -1060 3010 -1002 3066
rect -1060 2922 -1048 3010
rect -1014 2922 -1002 3010
rect -1060 2866 -1002 2922
rect -930 3010 -872 3066
rect -930 2922 -918 3010
rect -884 2922 -872 3010
rect -930 2866 -872 2922
rect -842 3010 -784 3066
rect -842 2922 -830 3010
rect -796 2922 -784 3010
rect -842 2866 -784 2922
rect -708 3008 -650 3064
rect -708 2920 -696 3008
rect -662 2920 -650 3008
rect -708 2864 -650 2920
rect -620 3008 -562 3064
rect -620 2920 -608 3008
rect -574 2920 -562 3008
rect -620 2864 -562 2920
rect 3812 3020 3870 3076
rect 3812 2932 3824 3020
rect 3858 2932 3870 3020
rect 3812 2876 3870 2932
rect 3900 3020 3958 3076
rect 3900 2932 3912 3020
rect 3946 2932 3958 3020
rect 3900 2876 3958 2932
rect 4028 3022 4086 3078
rect 4028 2934 4040 3022
rect 4074 2934 4086 3022
rect 4028 2878 4086 2934
rect 4116 3022 4174 3078
rect 4116 2934 4128 3022
rect 4162 2934 4174 3022
rect 4116 2878 4174 2934
rect 4246 3022 4304 3078
rect 4246 2934 4258 3022
rect 4292 2934 4304 3022
rect 4246 2878 4304 2934
rect 4334 3022 4392 3078
rect 4334 2934 4346 3022
rect 4380 2934 4392 3022
rect 4334 2878 4392 2934
rect 4468 3020 4526 3076
rect 4468 2932 4480 3020
rect 4514 2932 4526 3020
rect 4468 2876 4526 2932
rect 4556 3020 4614 3076
rect 4556 2932 4568 3020
rect 4602 2932 4614 3020
rect 4556 2876 4614 2932
rect 9468 2812 9526 2868
rect 9468 2724 9480 2812
rect 9514 2724 9526 2812
rect 9468 2668 9526 2724
rect 9556 2812 9614 2868
rect 9556 2724 9568 2812
rect 9602 2724 9614 2812
rect 9556 2668 9614 2724
rect 9684 2814 9742 2870
rect 9684 2726 9696 2814
rect 9730 2726 9742 2814
rect 9684 2670 9742 2726
rect 9772 2814 9830 2870
rect 9772 2726 9784 2814
rect 9818 2726 9830 2814
rect 9772 2670 9830 2726
rect 9902 2814 9960 2870
rect 9902 2726 9914 2814
rect 9948 2726 9960 2814
rect 9902 2670 9960 2726
rect 9990 2814 10048 2870
rect 9990 2726 10002 2814
rect 10036 2726 10048 2814
rect 9990 2670 10048 2726
rect 10124 2812 10182 2868
rect 10124 2724 10136 2812
rect 10170 2724 10182 2812
rect 10124 2668 10182 2724
rect 10212 2812 10270 2868
rect 10212 2724 10224 2812
rect 10258 2724 10270 2812
rect 10212 2668 10270 2724
rect 1138 2205 1196 2330
rect 1138 2055 1150 2205
rect 1184 2055 1196 2205
rect 1138 1930 1196 2055
rect 1396 2205 1454 2330
rect 1396 2055 1408 2205
rect 1442 2055 1454 2205
rect 1396 1930 1454 2055
rect 1654 2205 1712 2330
rect 1654 2055 1666 2205
rect 1700 2055 1712 2205
rect 1654 1930 1712 2055
rect 1912 2205 1970 2330
rect 1912 2055 1924 2205
rect 1958 2055 1970 2205
rect 1912 1930 1970 2055
rect 2152 2205 2210 2330
rect 2152 2055 2164 2205
rect 2198 2055 2210 2205
rect 2152 1930 2210 2055
rect 2410 2205 2468 2330
rect 2410 2055 2422 2205
rect 2456 2055 2468 2205
rect 2410 1930 2468 2055
rect 2668 2205 2726 2330
rect 2668 2055 2680 2205
rect 2714 2055 2726 2205
rect 2668 1930 2726 2055
rect 2926 2205 2984 2330
rect 2926 2055 2938 2205
rect 2972 2055 2984 2205
rect 2926 1930 2984 2055
rect 1138 1649 1196 1774
rect 1138 1499 1150 1649
rect 1184 1499 1196 1649
rect 1138 1374 1196 1499
rect 1396 1649 1454 1774
rect 1396 1499 1408 1649
rect 1442 1499 1454 1649
rect 1396 1374 1454 1499
rect 1654 1649 1712 1774
rect 1654 1499 1666 1649
rect 1700 1499 1712 1649
rect 1654 1374 1712 1499
rect 1912 1649 1970 1774
rect 1912 1499 1924 1649
rect 1958 1499 1970 1649
rect 1912 1374 1970 1499
rect 2152 1649 2210 1774
rect 2152 1499 2164 1649
rect 2198 1499 2210 1649
rect 2152 1374 2210 1499
rect 2410 1649 2468 1774
rect 2410 1499 2422 1649
rect 2456 1499 2468 1649
rect 2410 1374 2468 1499
rect 2668 1649 2726 1774
rect 2668 1499 2680 1649
rect 2714 1499 2726 1649
rect 2668 1374 2726 1499
rect 2926 1649 2984 1774
rect 2926 1499 2938 1649
rect 2972 1499 2984 1649
rect 2926 1374 2984 1499
rect -5022 1122 -4964 1178
rect -5022 1034 -5010 1122
rect -4976 1034 -4964 1122
rect -5022 978 -4964 1034
rect -4764 1122 -4706 1178
rect -4764 1034 -4752 1122
rect -4718 1034 -4706 1122
rect -4764 978 -4706 1034
rect -4546 1124 -4488 1180
rect -4546 1036 -4534 1124
rect -4500 1036 -4488 1124
rect -4546 980 -4488 1036
rect -3688 1124 -3630 1180
rect -3688 1036 -3676 1124
rect -3642 1036 -3630 1124
rect -3688 980 -3630 1036
rect -3574 1124 -3516 1180
rect -3574 1036 -3562 1124
rect -3528 1036 -3516 1124
rect -3574 980 -3516 1036
rect -2716 1124 -2658 1180
rect -2716 1036 -2704 1124
rect -2670 1036 -2658 1124
rect -2716 980 -2658 1036
rect -2488 1122 -2430 1178
rect -2488 1034 -2476 1122
rect -2442 1034 -2430 1122
rect -2488 978 -2430 1034
rect -2230 1122 -2172 1178
rect -2230 1034 -2218 1122
rect -2184 1034 -2172 1122
rect -2230 978 -2172 1034
rect 5670 1054 5728 1760
rect 1459 474 1517 530
rect 1459 386 1471 474
rect 1505 386 1517 474
rect 1459 330 1517 386
rect 1917 474 1975 530
rect 1917 386 1929 474
rect 1963 386 1975 474
rect 1917 330 1975 386
rect 2054 474 2112 530
rect 2054 386 2066 474
rect 2100 386 2112 474
rect 2054 330 2112 386
rect 2512 474 2570 530
rect 2512 386 2524 474
rect 2558 386 2570 474
rect 2512 330 2570 386
rect 5670 -334 5682 1054
rect 5716 -334 5728 1054
rect 5670 -1040 5728 -334
rect 5928 1054 5986 1760
rect 5928 -334 5940 1054
rect 5974 -334 5986 1054
rect 6220 1420 6278 1626
rect 6220 1032 6232 1420
rect 6266 1032 6278 1420
rect 6220 826 6278 1032
rect 6478 1420 6536 1626
rect 6478 1032 6490 1420
rect 6524 1032 6536 1420
rect 6478 826 6536 1032
rect 6736 1420 6794 1626
rect 6736 1032 6748 1420
rect 6782 1032 6794 1420
rect 6736 826 6794 1032
rect 6994 1420 7052 1626
rect 6994 1032 7006 1420
rect 7040 1032 7052 1420
rect 6994 826 7052 1032
rect 7220 1420 7278 1626
rect 7220 1032 7232 1420
rect 7266 1032 7278 1420
rect 7220 826 7278 1032
rect 7478 1420 7536 1626
rect 7478 1032 7490 1420
rect 7524 1032 7536 1420
rect 7478 826 7536 1032
rect 7736 1420 7794 1626
rect 7736 1032 7748 1420
rect 7782 1032 7794 1420
rect 7736 826 7794 1032
rect 7994 1420 8052 1626
rect 7994 1032 8006 1420
rect 8040 1032 8052 1420
rect 7994 826 8052 1032
rect 8268 1004 8326 1710
rect 6220 464 6278 670
rect 6220 76 6232 464
rect 6266 76 6278 464
rect 6220 -130 6278 76
rect 6478 464 6536 670
rect 6478 76 6490 464
rect 6524 76 6536 464
rect 6478 -130 6536 76
rect 6736 464 6794 670
rect 6736 76 6748 464
rect 6782 76 6794 464
rect 6736 -130 6794 76
rect 6994 464 7052 670
rect 6994 76 7006 464
rect 7040 76 7052 464
rect 6994 -130 7052 76
rect 7220 464 7278 670
rect 7220 76 7232 464
rect 7266 76 7278 464
rect 7220 -130 7278 76
rect 7478 464 7536 670
rect 7478 76 7490 464
rect 7524 76 7536 464
rect 7478 -130 7536 76
rect 7736 464 7794 670
rect 7736 76 7748 464
rect 7782 76 7794 464
rect 7736 -130 7794 76
rect 7994 464 8052 670
rect 7994 76 8006 464
rect 8040 76 8052 464
rect 7994 -130 8052 76
rect 5928 -1040 5986 -334
rect 6220 -492 6278 -286
rect 6220 -880 6232 -492
rect 6266 -880 6278 -492
rect 6220 -1086 6278 -880
rect 6478 -492 6536 -286
rect 6478 -880 6490 -492
rect 6524 -880 6536 -492
rect 6478 -1086 6536 -880
rect 6736 -492 6794 -286
rect 6736 -880 6748 -492
rect 6782 -880 6794 -492
rect 6736 -1086 6794 -880
rect 6994 -492 7052 -286
rect 6994 -880 7006 -492
rect 7040 -880 7052 -492
rect 6994 -1086 7052 -880
rect 7220 -492 7278 -286
rect 7220 -880 7232 -492
rect 7266 -880 7278 -492
rect 7220 -1086 7278 -880
rect 7478 -492 7536 -286
rect 7478 -880 7490 -492
rect 7524 -880 7536 -492
rect 7478 -1086 7536 -880
rect 7736 -492 7794 -286
rect 7736 -880 7748 -492
rect 7782 -880 7794 -492
rect 7736 -1086 7794 -880
rect 7994 -492 8052 -286
rect 7994 -880 8006 -492
rect 8040 -880 8052 -492
rect 7994 -1086 8052 -880
rect 8268 -384 8280 1004
rect 8314 -384 8326 1004
rect 8268 -1090 8326 -384
rect 8526 1004 8584 1710
rect 8526 -384 8538 1004
rect 8572 -384 8584 1004
rect 8526 -1090 8584 -384
<< pdiff >>
rect -5028 4306 -4970 4562
rect -5028 3818 -5016 4306
rect -4982 3818 -4970 4306
rect -6574 3578 -6516 3684
rect -6574 3390 -6562 3578
rect -6528 3390 -6516 3578
rect -6574 3284 -6516 3390
rect -6486 3578 -6428 3684
rect -6486 3390 -6474 3578
rect -6440 3390 -6428 3578
rect -6486 3284 -6428 3390
rect -6342 3576 -6284 3682
rect -6342 3388 -6330 3576
rect -6296 3388 -6284 3576
rect -6342 3282 -6284 3388
rect -6254 3576 -6196 3682
rect -6254 3388 -6242 3576
rect -6208 3388 -6196 3576
rect -6254 3282 -6196 3388
rect -6114 3574 -6056 3680
rect -6114 3386 -6102 3574
rect -6068 3386 -6056 3574
rect -6114 3280 -6056 3386
rect -6026 3574 -5968 3680
rect -6026 3386 -6014 3574
rect -5980 3386 -5968 3574
rect -6026 3280 -5968 3386
rect -5896 3576 -5838 3682
rect -5896 3388 -5884 3576
rect -5850 3388 -5838 3576
rect -5896 3282 -5838 3388
rect -5808 3576 -5750 3682
rect -5808 3388 -5796 3576
rect -5762 3388 -5750 3576
rect -5028 3562 -4970 3818
rect -4770 4306 -4712 4562
rect -4770 3818 -4758 4306
rect -4724 3818 -4712 4306
rect -4770 3562 -4712 3818
rect -4372 4314 -4314 4570
rect -4372 3826 -4360 4314
rect -4326 3826 -4314 4314
rect -4372 3570 -4314 3826
rect -4114 4314 -4056 4570
rect -4114 3826 -4102 4314
rect -4068 3826 -4056 4314
rect -4114 3570 -4056 3826
rect -3856 4314 -3798 4570
rect -3856 3826 -3844 4314
rect -3810 3826 -3798 4314
rect -3856 3570 -3798 3826
rect -3372 4314 -3314 4570
rect -3372 3826 -3360 4314
rect -3326 3826 -3314 4314
rect -3372 3570 -3314 3826
rect -3114 4314 -3056 4570
rect -3114 3826 -3102 4314
rect -3068 3826 -3056 4314
rect -3114 3570 -3056 3826
rect -2856 4314 -2798 4570
rect -2856 3826 -2844 4314
rect -2810 3826 -2798 4314
rect -2856 3570 -2798 3826
rect -2466 4318 -2408 4574
rect -2466 3830 -2454 4318
rect -2420 3830 -2408 4318
rect -2466 3574 -2408 3830
rect -2208 4318 -2150 4574
rect -2208 3830 -2196 4318
rect -2162 3830 -2150 4318
rect -2208 3574 -2150 3830
rect 908 4046 966 4302
rect -1388 3596 -1330 3702
rect -5808 3282 -5750 3388
rect -1388 3408 -1376 3596
rect -1342 3408 -1330 3596
rect -1388 3302 -1330 3408
rect -1300 3596 -1242 3702
rect -1300 3408 -1288 3596
rect -1254 3408 -1242 3596
rect -1300 3302 -1242 3408
rect -1156 3594 -1098 3700
rect -1156 3406 -1144 3594
rect -1110 3406 -1098 3594
rect -1156 3300 -1098 3406
rect -1068 3594 -1010 3700
rect -1068 3406 -1056 3594
rect -1022 3406 -1010 3594
rect -1068 3300 -1010 3406
rect -928 3592 -870 3698
rect -928 3404 -916 3592
rect -882 3404 -870 3592
rect -928 3298 -870 3404
rect -840 3592 -782 3698
rect -840 3404 -828 3592
rect -794 3404 -782 3592
rect -840 3298 -782 3404
rect -710 3594 -652 3700
rect -710 3406 -698 3594
rect -664 3406 -652 3594
rect -710 3300 -652 3406
rect -622 3594 -564 3700
rect -622 3406 -610 3594
rect -576 3406 -564 3594
rect -622 3300 -564 3406
rect 908 3558 920 4046
rect 954 3558 966 4046
rect 908 3302 966 3558
rect 1166 4046 1224 4302
rect 1166 3558 1178 4046
rect 1212 3558 1224 4046
rect 1166 3302 1224 3558
rect 1387 4038 1445 4294
rect 1387 3550 1399 4038
rect 1433 3550 1445 4038
rect 1387 3294 1445 3550
rect 1645 4038 1703 4294
rect 1645 3550 1657 4038
rect 1691 3550 1703 4038
rect 1645 3294 1703 3550
rect 1903 4038 1961 4294
rect 1903 3550 1915 4038
rect 1949 3550 1961 4038
rect 1903 3294 1961 3550
rect 2045 4040 2103 4296
rect 2045 3552 2057 4040
rect 2091 3552 2103 4040
rect 2045 3296 2103 3552
rect 2303 4040 2361 4296
rect 2303 3686 2315 4040
rect 2349 3686 2361 4040
rect 2303 3296 2361 3686
rect 2561 4040 2619 4296
rect 2561 3552 2573 4040
rect 2607 3552 2619 4040
rect 2561 3296 2619 3552
rect 2702 4020 2760 4276
rect 2702 3532 2714 4020
rect 2748 3532 2760 4020
rect 2702 3276 2760 3532
rect 2960 4020 3018 4276
rect 2960 3532 2972 4020
rect 3006 3532 3018 4020
rect 6182 3918 6240 4174
rect 2960 3276 3018 3532
rect 3788 3608 3846 3714
rect 3788 3420 3800 3608
rect 3834 3420 3846 3608
rect 3788 3314 3846 3420
rect 3876 3608 3934 3714
rect 3876 3420 3888 3608
rect 3922 3420 3934 3608
rect 3876 3314 3934 3420
rect 4020 3606 4078 3712
rect 4020 3418 4032 3606
rect 4066 3418 4078 3606
rect 4020 3312 4078 3418
rect 4108 3606 4166 3712
rect 4108 3418 4120 3606
rect 4154 3418 4166 3606
rect 4108 3312 4166 3418
rect 4248 3604 4306 3710
rect 4248 3416 4260 3604
rect 4294 3416 4306 3604
rect 4248 3310 4306 3416
rect 4336 3604 4394 3710
rect 4336 3416 4348 3604
rect 4382 3416 4394 3604
rect 4336 3310 4394 3416
rect 4466 3606 4524 3712
rect 4466 3418 4478 3606
rect 4512 3418 4524 3606
rect 4466 3312 4524 3418
rect 4554 3606 4612 3712
rect 4554 3418 4566 3606
rect 4600 3418 4612 3606
rect 4554 3312 4612 3418
rect 6182 3430 6194 3918
rect 6228 3430 6240 3918
rect 6182 3174 6240 3430
rect 6440 3918 6498 4174
rect 6440 3430 6452 3918
rect 6486 3430 6498 3918
rect 6440 3174 6498 3430
rect 6576 3900 6634 4156
rect 6576 3412 6588 3900
rect 6622 3412 6634 3900
rect 6576 3156 6634 3412
rect 7034 3900 7092 4156
rect 7034 3412 7046 3900
rect 7080 3412 7092 3900
rect 7034 3156 7092 3412
rect 7148 3900 7206 4156
rect 7148 3412 7160 3900
rect 7194 3412 7206 3900
rect 7148 3156 7206 3412
rect 7606 3900 7664 4156
rect 7606 3412 7618 3900
rect 7652 3412 7664 3900
rect 7606 3156 7664 3412
rect 7770 3930 7828 4186
rect 7770 3442 7782 3930
rect 7816 3442 7828 3930
rect 7770 3186 7828 3442
rect 8028 3930 8086 4186
rect 8028 3442 8040 3930
rect 8074 3442 8086 3930
rect 8028 3186 8086 3442
rect 9444 3400 9502 3506
rect 9444 3212 9456 3400
rect 9490 3212 9502 3400
rect 9444 3106 9502 3212
rect 9532 3400 9590 3506
rect 9532 3212 9544 3400
rect 9578 3212 9590 3400
rect 9532 3106 9590 3212
rect 9676 3398 9734 3504
rect 9676 3210 9688 3398
rect 9722 3210 9734 3398
rect 9676 3104 9734 3210
rect 9764 3398 9822 3504
rect 9764 3210 9776 3398
rect 9810 3210 9822 3398
rect 9764 3104 9822 3210
rect 9904 3396 9962 3502
rect 9904 3208 9916 3396
rect 9950 3208 9962 3396
rect 9904 3102 9962 3208
rect 9992 3396 10050 3502
rect 9992 3208 10004 3396
rect 10038 3208 10050 3396
rect 9992 3102 10050 3208
rect 10122 3398 10180 3504
rect 10122 3210 10134 3398
rect 10168 3210 10180 3398
rect 10122 3104 10180 3210
rect 10210 3398 10268 3504
rect 10210 3210 10222 3398
rect 10256 3210 10268 3398
rect 10210 3104 10268 3210
<< ndiffc >>
rect -6538 2902 -6504 2990
rect -6450 2902 -6416 2990
rect -6322 2904 -6288 2992
rect -6234 2904 -6200 2992
rect -6104 2904 -6070 2992
rect -6016 2904 -5982 2992
rect -5882 2902 -5848 2990
rect -5794 2902 -5760 2990
rect -1352 2920 -1318 3008
rect -1264 2920 -1230 3008
rect -1136 2922 -1102 3010
rect -1048 2922 -1014 3010
rect -918 2922 -884 3010
rect -830 2922 -796 3010
rect -696 2920 -662 3008
rect -608 2920 -574 3008
rect 3824 2932 3858 3020
rect 3912 2932 3946 3020
rect 4040 2934 4074 3022
rect 4128 2934 4162 3022
rect 4258 2934 4292 3022
rect 4346 2934 4380 3022
rect 4480 2932 4514 3020
rect 4568 2932 4602 3020
rect 9480 2724 9514 2812
rect 9568 2724 9602 2812
rect 9696 2726 9730 2814
rect 9784 2726 9818 2814
rect 9914 2726 9948 2814
rect 10002 2726 10036 2814
rect 10136 2724 10170 2812
rect 10224 2724 10258 2812
rect 1150 2055 1184 2205
rect 1408 2055 1442 2205
rect 1666 2055 1700 2205
rect 1924 2055 1958 2205
rect 2164 2055 2198 2205
rect 2422 2055 2456 2205
rect 2680 2055 2714 2205
rect 2938 2055 2972 2205
rect 1150 1499 1184 1649
rect 1408 1499 1442 1649
rect 1666 1499 1700 1649
rect 1924 1499 1958 1649
rect 2164 1499 2198 1649
rect 2422 1499 2456 1649
rect 2680 1499 2714 1649
rect 2938 1499 2972 1649
rect -5010 1034 -4976 1122
rect -4752 1034 -4718 1122
rect -4534 1036 -4500 1124
rect -3676 1036 -3642 1124
rect -3562 1036 -3528 1124
rect -2704 1036 -2670 1124
rect -2476 1034 -2442 1122
rect -2218 1034 -2184 1122
rect 1471 386 1505 474
rect 1929 386 1963 474
rect 2066 386 2100 474
rect 2524 386 2558 474
rect 5682 -334 5716 1054
rect 5940 -334 5974 1054
rect 6232 1032 6266 1420
rect 6490 1032 6524 1420
rect 6748 1032 6782 1420
rect 7006 1032 7040 1420
rect 7232 1032 7266 1420
rect 7490 1032 7524 1420
rect 7748 1032 7782 1420
rect 8006 1032 8040 1420
rect 6232 76 6266 464
rect 6490 76 6524 464
rect 6748 76 6782 464
rect 7006 76 7040 464
rect 7232 76 7266 464
rect 7490 76 7524 464
rect 7748 76 7782 464
rect 8006 76 8040 464
rect 6232 -880 6266 -492
rect 6490 -880 6524 -492
rect 6748 -880 6782 -492
rect 7006 -880 7040 -492
rect 7232 -880 7266 -492
rect 7490 -880 7524 -492
rect 7748 -880 7782 -492
rect 8006 -880 8040 -492
rect 8280 -384 8314 1004
rect 8538 -384 8572 1004
<< pdiffc >>
rect -5016 3818 -4982 4306
rect -6562 3390 -6528 3578
rect -6474 3390 -6440 3578
rect -6330 3388 -6296 3576
rect -6242 3388 -6208 3576
rect -6102 3386 -6068 3574
rect -6014 3386 -5980 3574
rect -5884 3388 -5850 3576
rect -5796 3388 -5762 3576
rect -4758 3818 -4724 4306
rect -4360 3826 -4326 4314
rect -4102 3826 -4068 4314
rect -3844 3826 -3810 4314
rect -3360 3826 -3326 4314
rect -3102 3826 -3068 4314
rect -2844 3826 -2810 4314
rect -2454 3830 -2420 4318
rect -2196 3830 -2162 4318
rect -1376 3408 -1342 3596
rect -1288 3408 -1254 3596
rect -1144 3406 -1110 3594
rect -1056 3406 -1022 3594
rect -916 3404 -882 3592
rect -828 3404 -794 3592
rect -698 3406 -664 3594
rect -610 3406 -576 3594
rect 920 3558 954 4046
rect 1178 3558 1212 4046
rect 1399 3550 1433 4038
rect 1657 3550 1691 4038
rect 1915 3550 1949 4038
rect 2057 3552 2091 4040
rect 2315 3686 2349 4040
rect 2573 3552 2607 4040
rect 2714 3532 2748 4020
rect 2972 3532 3006 4020
rect 3800 3420 3834 3608
rect 3888 3420 3922 3608
rect 4032 3418 4066 3606
rect 4120 3418 4154 3606
rect 4260 3416 4294 3604
rect 4348 3416 4382 3604
rect 4478 3418 4512 3606
rect 4566 3418 4600 3606
rect 6194 3430 6228 3918
rect 6452 3430 6486 3918
rect 6588 3412 6622 3900
rect 7046 3412 7080 3900
rect 7160 3412 7194 3900
rect 7618 3412 7652 3900
rect 7782 3442 7816 3930
rect 8040 3442 8074 3930
rect 9456 3212 9490 3400
rect 9544 3212 9578 3400
rect 9688 3210 9722 3398
rect 9776 3210 9810 3398
rect 9916 3208 9950 3396
rect 10004 3208 10038 3396
rect 10134 3210 10168 3398
rect 10222 3210 10256 3398
<< psubdiff >>
rect 10156 10714 11468 10908
rect 10156 10220 10364 10714
rect 11324 10220 11468 10714
rect 10156 10000 11468 10220
rect -4320 344 -3008 538
rect -4320 -150 -4112 344
rect -3152 -150 -3008 344
rect -4320 -370 -3008 -150
rect 3102 160 4414 354
rect 3102 -334 3310 160
rect 4270 -334 4414 160
rect 3102 -554 4414 -334
rect 9734 478 11046 672
rect 9734 -16 9942 478
rect 10902 -16 11046 478
rect 9734 -236 11046 -16
<< nsubdiff >>
rect -6356 4662 -5842 4758
rect -1468 4740 -954 4836
rect -6356 4422 -6262 4662
rect -5936 4422 -5842 4662
rect -6356 4324 -5842 4422
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect -1468 4402 -954 4500
rect 3844 4528 4358 4624
rect 3844 4288 3938 4528
rect 4264 4288 4358 4528
rect 3844 4190 4358 4288
rect 9280 4470 9794 4566
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
<< psubdiffcont >>
rect 10364 10220 11324 10714
rect -4112 -150 -3152 344
rect 3310 -334 4270 160
rect 9942 -16 10902 478
<< nsubdiffcont >>
rect -6262 4422 -5936 4662
rect -1374 4500 -1048 4740
rect 3938 4288 4264 4528
rect 9374 4230 9700 4470
<< poly >>
rect -4928 4643 -4812 4659
rect -4928 4626 -4912 4643
rect -4970 4609 -4912 4626
rect -4828 4626 -4812 4643
rect -4272 4651 -4156 4667
rect -4272 4634 -4256 4651
rect -4828 4609 -4770 4626
rect -4970 4562 -4770 4609
rect -4314 4617 -4256 4634
rect -4172 4634 -4156 4651
rect -4014 4651 -3898 4667
rect -4014 4634 -3998 4651
rect -4172 4617 -4114 4634
rect -4314 4570 -4114 4617
rect -4056 4617 -3998 4634
rect -3914 4634 -3898 4651
rect -3272 4651 -3156 4667
rect -3272 4634 -3256 4651
rect -3914 4617 -3856 4634
rect -4056 4570 -3856 4617
rect -3314 4617 -3256 4634
rect -3172 4634 -3156 4651
rect -3014 4651 -2898 4667
rect -3014 4634 -2998 4651
rect -3172 4617 -3114 4634
rect -3314 4570 -3114 4617
rect -3056 4617 -2998 4634
rect -2914 4634 -2898 4651
rect -2366 4655 -2250 4671
rect -2366 4638 -2350 4655
rect -2914 4617 -2856 4634
rect -3056 4570 -2856 4617
rect -2408 4621 -2350 4638
rect -2266 4638 -2250 4655
rect -2266 4621 -2208 4638
rect -2408 4574 -2208 4621
rect -6534 3765 -6468 3781
rect -6534 3731 -6518 3765
rect -6484 3731 -6468 3765
rect -6534 3715 -6468 3731
rect -6302 3763 -6236 3779
rect -6302 3729 -6286 3763
rect -6252 3729 -6236 3763
rect -6516 3684 -6486 3715
rect -6302 3713 -6236 3729
rect -6074 3761 -6008 3777
rect -6074 3727 -6058 3761
rect -6024 3727 -6008 3761
rect -6284 3682 -6254 3713
rect -6074 3711 -6008 3727
rect -5856 3763 -5790 3779
rect -5856 3729 -5840 3763
rect -5806 3729 -5790 3763
rect -5856 3713 -5790 3729
rect -6516 3253 -6486 3284
rect -6056 3680 -6026 3711
rect -5838 3682 -5808 3713
rect -6534 3237 -6468 3253
rect -6284 3251 -6254 3282
rect 1008 4383 1124 4399
rect 1008 4366 1024 4383
rect 966 4349 1024 4366
rect 1108 4366 1124 4383
rect 1487 4375 1603 4391
rect 1108 4349 1166 4366
rect 1487 4358 1503 4375
rect 966 4302 1166 4349
rect 1445 4341 1503 4358
rect 1587 4358 1603 4375
rect 1745 4375 1861 4391
rect 1745 4358 1761 4375
rect 1587 4341 1645 4358
rect -1348 3783 -1282 3799
rect -1348 3749 -1332 3783
rect -1298 3749 -1282 3783
rect -1348 3733 -1282 3749
rect -1116 3781 -1050 3797
rect -1116 3747 -1100 3781
rect -1066 3747 -1050 3781
rect -1330 3702 -1300 3733
rect -1116 3731 -1050 3747
rect -888 3779 -822 3795
rect -888 3745 -872 3779
rect -838 3745 -822 3779
rect -4970 3536 -4770 3562
rect -4314 3544 -4114 3570
rect -4056 3544 -3856 3570
rect -3314 3544 -3114 3570
rect -3056 3544 -2856 3570
rect -2408 3548 -2208 3574
rect -1098 3700 -1068 3731
rect -888 3729 -822 3745
rect -670 3781 -604 3797
rect -670 3747 -654 3781
rect -620 3747 -604 3781
rect -670 3731 -604 3747
rect -6534 3203 -6518 3237
rect -6484 3203 -6468 3237
rect -6534 3187 -6468 3203
rect -6302 3235 -6236 3251
rect -6056 3249 -6026 3280
rect -5838 3251 -5808 3282
rect -1330 3271 -1300 3302
rect -870 3698 -840 3729
rect -652 3700 -622 3731
rect -1348 3255 -1282 3271
rect -1098 3269 -1068 3300
rect 1445 4294 1645 4341
rect 1703 4341 1761 4358
rect 1845 4358 1861 4375
rect 2145 4377 2261 4393
rect 2145 4360 2161 4377
rect 1845 4341 1903 4358
rect 1703 4294 1903 4341
rect 2105 4343 2161 4360
rect 2245 4360 2261 4377
rect 2403 4377 2519 4393
rect 2403 4360 2419 4377
rect 2245 4343 2303 4360
rect 2105 4322 2303 4343
rect 2103 4296 2303 4322
rect 2361 4343 2419 4360
rect 2503 4360 2519 4377
rect 2503 4343 2561 4360
rect 2361 4296 2561 4343
rect 2802 4357 2918 4373
rect 2802 4340 2818 4357
rect 2760 4323 2818 4340
rect 2902 4340 2918 4357
rect 2902 4323 2960 4340
rect -6302 3201 -6286 3235
rect -6252 3201 -6236 3235
rect -6302 3185 -6236 3201
rect -6074 3233 -6008 3249
rect -6074 3199 -6058 3233
rect -6024 3199 -6008 3233
rect -6074 3183 -6008 3199
rect -5856 3235 -5790 3251
rect -5856 3201 -5840 3235
rect -5806 3201 -5790 3235
rect -1348 3221 -1332 3255
rect -1298 3221 -1282 3255
rect -1348 3205 -1282 3221
rect -1116 3253 -1050 3269
rect -870 3267 -840 3298
rect -652 3269 -622 3300
rect 966 3276 1166 3302
rect 2760 4276 2960 4323
rect -1116 3219 -1100 3253
rect -1066 3219 -1050 3253
rect -1116 3203 -1050 3219
rect -888 3251 -822 3267
rect -888 3217 -872 3251
rect -838 3217 -822 3251
rect -888 3201 -822 3217
rect -670 3253 -604 3269
rect 1445 3268 1645 3294
rect 1703 3268 1903 3294
rect 2103 3270 2303 3296
rect 2361 3270 2561 3296
rect 6282 4255 6398 4271
rect 6282 4238 6298 4255
rect 6240 4221 6298 4238
rect 6382 4238 6398 4255
rect 7870 4267 7986 4283
rect 6382 4221 6440 4238
rect 6240 4174 6440 4221
rect 6726 4237 6942 4253
rect 6726 4220 6742 4237
rect 6634 4203 6742 4220
rect 6926 4220 6942 4237
rect 7298 4237 7514 4253
rect 7870 4250 7886 4267
rect 7298 4220 7314 4237
rect 6926 4203 7034 4220
rect 3828 3795 3894 3811
rect 3828 3761 3844 3795
rect 3878 3761 3894 3795
rect 3828 3745 3894 3761
rect 4060 3793 4126 3809
rect 4060 3759 4076 3793
rect 4110 3759 4126 3793
rect 3846 3714 3876 3745
rect 4060 3743 4126 3759
rect 4288 3791 4354 3807
rect 4288 3757 4304 3791
rect 4338 3757 4354 3791
rect 4078 3712 4108 3743
rect 4288 3741 4354 3757
rect 4506 3793 4572 3809
rect 4506 3759 4522 3793
rect 4556 3759 4572 3793
rect 4506 3743 4572 3759
rect 3846 3283 3876 3314
rect 4306 3710 4336 3741
rect 4524 3712 4554 3743
rect -670 3219 -654 3253
rect -620 3219 -604 3253
rect 2760 3250 2960 3276
rect 3828 3267 3894 3283
rect 4078 3281 4108 3312
rect -670 3203 -604 3219
rect 3828 3233 3844 3267
rect 3878 3233 3894 3267
rect 3828 3217 3894 3233
rect 4060 3265 4126 3281
rect 4306 3279 4336 3310
rect 4524 3281 4554 3312
rect 4060 3231 4076 3265
rect 4110 3231 4126 3265
rect 4060 3215 4126 3231
rect 4288 3263 4354 3279
rect 4288 3229 4304 3263
rect 4338 3229 4354 3263
rect 4288 3213 4354 3229
rect 4506 3265 4572 3281
rect 4506 3231 4522 3265
rect 4556 3231 4572 3265
rect 4506 3215 4572 3231
rect -5856 3185 -5790 3201
rect 6634 4156 7034 4203
rect 7206 4203 7314 4220
rect 7498 4220 7514 4237
rect 7828 4233 7886 4250
rect 7970 4250 7986 4267
rect 7970 4233 8028 4250
rect 7498 4203 7606 4220
rect 7206 4156 7606 4203
rect 7828 4186 8028 4233
rect -1324 3136 -1258 3152
rect -6510 3118 -6444 3134
rect -6510 3084 -6494 3118
rect -6460 3084 -6444 3118
rect -6510 3068 -6444 3084
rect -6294 3120 -6228 3136
rect -6294 3086 -6278 3120
rect -6244 3086 -6228 3120
rect -6294 3070 -6228 3086
rect -6076 3120 -6010 3136
rect -6076 3086 -6060 3120
rect -6026 3086 -6010 3120
rect -6076 3070 -6010 3086
rect -5854 3118 -5788 3134
rect -5854 3084 -5838 3118
rect -5804 3084 -5788 3118
rect -1324 3102 -1308 3136
rect -1274 3102 -1258 3136
rect -1324 3086 -1258 3102
rect -1108 3138 -1042 3154
rect -1108 3104 -1092 3138
rect -1058 3104 -1042 3138
rect -1108 3088 -1042 3104
rect -890 3138 -824 3154
rect -890 3104 -874 3138
rect -840 3104 -824 3138
rect -890 3088 -824 3104
rect -668 3136 -602 3152
rect -668 3102 -652 3136
rect -618 3102 -602 3136
rect -6492 3046 -6462 3068
rect -6276 3048 -6246 3070
rect -6058 3048 -6028 3070
rect -5854 3068 -5788 3084
rect -5836 3046 -5806 3068
rect -1306 3064 -1276 3086
rect -1090 3066 -1060 3088
rect -872 3066 -842 3088
rect -668 3086 -602 3102
rect 3852 3148 3918 3164
rect 3852 3114 3868 3148
rect 3902 3114 3918 3148
rect 3852 3098 3918 3114
rect 4068 3150 4134 3166
rect 4068 3116 4084 3150
rect 4118 3116 4134 3150
rect 4068 3100 4134 3116
rect 4286 3150 4352 3166
rect 4286 3116 4302 3150
rect 4336 3116 4352 3150
rect 4286 3100 4352 3116
rect 4508 3148 4574 3164
rect 6240 3148 6440 3174
rect 9484 3587 9550 3603
rect 9484 3553 9500 3587
rect 9534 3553 9550 3587
rect 9484 3537 9550 3553
rect 9716 3585 9782 3601
rect 9716 3551 9732 3585
rect 9766 3551 9782 3585
rect 9502 3506 9532 3537
rect 9716 3535 9782 3551
rect 9944 3583 10010 3599
rect 9944 3549 9960 3583
rect 9994 3549 10010 3583
rect 7828 3160 8028 3186
rect 4508 3114 4524 3148
rect 4558 3114 4574 3148
rect 6634 3130 7034 3156
rect 7206 3130 7606 3156
rect -6492 2824 -6462 2846
rect -6276 2826 -6246 2848
rect -6058 2826 -6028 2848
rect -650 3064 -620 3086
rect 3870 3076 3900 3098
rect 4086 3078 4116 3100
rect 4304 3078 4334 3100
rect 4508 3098 4574 3114
rect 9734 3504 9764 3535
rect 9944 3533 10010 3549
rect 10162 3585 10228 3601
rect 10162 3551 10178 3585
rect 10212 3551 10228 3585
rect 10162 3535 10228 3551
rect -6510 2808 -6444 2824
rect -6510 2774 -6494 2808
rect -6460 2774 -6444 2808
rect -6510 2758 -6444 2774
rect -6294 2810 -6228 2826
rect -6294 2776 -6278 2810
rect -6244 2776 -6228 2810
rect -6294 2760 -6228 2776
rect -6076 2810 -6010 2826
rect -5836 2824 -5806 2846
rect -1306 2842 -1276 2864
rect -1090 2844 -1060 2866
rect -872 2844 -842 2866
rect 4526 3076 4556 3098
rect -1324 2826 -1258 2842
rect -6076 2776 -6060 2810
rect -6026 2776 -6010 2810
rect -6076 2760 -6010 2776
rect -5854 2808 -5788 2824
rect -5854 2774 -5838 2808
rect -5804 2774 -5788 2808
rect -1324 2792 -1308 2826
rect -1274 2792 -1258 2826
rect -1324 2776 -1258 2792
rect -1108 2828 -1042 2844
rect -1108 2794 -1092 2828
rect -1058 2794 -1042 2828
rect -1108 2778 -1042 2794
rect -890 2828 -824 2844
rect -650 2842 -620 2864
rect 3870 2854 3900 2876
rect 4086 2856 4116 2878
rect 4304 2856 4334 2878
rect 9502 3075 9532 3106
rect 9962 3502 9992 3533
rect 10180 3504 10210 3535
rect 9484 3059 9550 3075
rect 9734 3073 9764 3104
rect 9484 3025 9500 3059
rect 9534 3025 9550 3059
rect 9484 3009 9550 3025
rect 9716 3057 9782 3073
rect 9962 3071 9992 3102
rect 10180 3073 10210 3104
rect 9716 3023 9732 3057
rect 9766 3023 9782 3057
rect 9716 3007 9782 3023
rect 9944 3055 10010 3071
rect 9944 3021 9960 3055
rect 9994 3021 10010 3055
rect 9944 3005 10010 3021
rect 10162 3057 10228 3073
rect 10162 3023 10178 3057
rect 10212 3023 10228 3057
rect 10162 3007 10228 3023
rect 9508 2940 9574 2956
rect 9508 2906 9524 2940
rect 9558 2906 9574 2940
rect 9508 2890 9574 2906
rect 9724 2942 9790 2958
rect 9724 2908 9740 2942
rect 9774 2908 9790 2942
rect 9724 2892 9790 2908
rect 9942 2942 10008 2958
rect 9942 2908 9958 2942
rect 9992 2908 10008 2942
rect 9942 2892 10008 2908
rect 10164 2940 10230 2956
rect 10164 2906 10180 2940
rect 10214 2906 10230 2940
rect -890 2794 -874 2828
rect -840 2794 -824 2828
rect -890 2778 -824 2794
rect -668 2826 -602 2842
rect -668 2792 -652 2826
rect -618 2792 -602 2826
rect -668 2776 -602 2792
rect 3852 2838 3918 2854
rect 3852 2804 3868 2838
rect 3902 2804 3918 2838
rect 3852 2788 3918 2804
rect 4068 2840 4134 2856
rect 4068 2806 4084 2840
rect 4118 2806 4134 2840
rect 4068 2790 4134 2806
rect 4286 2840 4352 2856
rect 4526 2854 4556 2876
rect 9526 2868 9556 2890
rect 9742 2870 9772 2892
rect 9960 2870 9990 2892
rect 10164 2890 10230 2906
rect 4286 2806 4302 2840
rect 4336 2806 4352 2840
rect 4286 2790 4352 2806
rect 4508 2838 4574 2854
rect 4508 2804 4524 2838
rect 4558 2804 4574 2838
rect 4508 2788 4574 2804
rect -5854 2758 -5788 2774
rect 10182 2868 10212 2890
rect 9526 2646 9556 2668
rect 9742 2648 9772 2670
rect 9960 2648 9990 2670
rect 9508 2630 9574 2646
rect 9508 2596 9524 2630
rect 9558 2596 9574 2630
rect 9508 2580 9574 2596
rect 9724 2632 9790 2648
rect 9724 2598 9740 2632
rect 9774 2598 9790 2632
rect 9724 2582 9790 2598
rect 9942 2632 10008 2648
rect 10182 2646 10212 2668
rect 9942 2598 9958 2632
rect 9992 2598 10008 2632
rect 9942 2582 10008 2598
rect 10164 2630 10230 2646
rect 10164 2596 10180 2630
rect 10214 2596 10230 2630
rect 10164 2580 10230 2596
rect 1246 2402 1346 2418
rect 1246 2385 1262 2402
rect 1196 2368 1262 2385
rect 1330 2385 1346 2402
rect 1504 2402 1604 2418
rect 1504 2385 1520 2402
rect 1330 2368 1396 2385
rect 1196 2330 1396 2368
rect 1454 2368 1520 2385
rect 1588 2385 1604 2402
rect 1762 2402 1862 2418
rect 1762 2385 1778 2402
rect 1588 2368 1654 2385
rect 1454 2330 1654 2368
rect 1712 2368 1778 2385
rect 1846 2385 1862 2402
rect 2260 2402 2360 2418
rect 2260 2385 2276 2402
rect 1846 2368 1912 2385
rect 1712 2330 1912 2368
rect 2210 2368 2276 2385
rect 2344 2385 2360 2402
rect 2518 2402 2618 2418
rect 2518 2385 2534 2402
rect 2344 2368 2410 2385
rect 2210 2330 2410 2368
rect 2468 2368 2534 2385
rect 2602 2385 2618 2402
rect 2776 2402 2876 2418
rect 2776 2385 2792 2402
rect 2602 2368 2668 2385
rect 2468 2330 2668 2368
rect 2726 2368 2792 2385
rect 2860 2385 2876 2402
rect 2860 2368 2926 2385
rect 2726 2330 2926 2368
rect 1196 1904 1396 1930
rect 1454 1904 1654 1930
rect 1712 1904 1912 1930
rect 2210 1904 2410 1930
rect 2468 1904 2668 1930
rect 2726 1904 2926 1930
rect 1246 1846 1346 1862
rect 1246 1829 1262 1846
rect 1196 1812 1262 1829
rect 1330 1829 1346 1846
rect 1504 1846 1604 1862
rect 1504 1829 1520 1846
rect 1330 1812 1396 1829
rect 1196 1774 1396 1812
rect 1454 1812 1520 1829
rect 1588 1829 1604 1846
rect 1762 1846 1862 1862
rect 1762 1829 1778 1846
rect 1588 1812 1654 1829
rect 1454 1774 1654 1812
rect 1712 1812 1778 1829
rect 1846 1829 1862 1846
rect 2260 1846 2360 1862
rect 2260 1829 2276 1846
rect 1846 1812 1912 1829
rect 1712 1774 1912 1812
rect 2210 1812 2276 1829
rect 2344 1829 2360 1846
rect 2518 1846 2618 1862
rect 2518 1829 2534 1846
rect 2344 1812 2410 1829
rect 2210 1774 2410 1812
rect 2468 1812 2534 1829
rect 2602 1829 2618 1846
rect 2776 1846 2876 1862
rect 2776 1829 2792 1846
rect 2602 1812 2668 1829
rect 2468 1774 2668 1812
rect 2726 1812 2792 1829
rect 2860 1829 2876 1846
rect 5770 1832 5886 1848
rect 2860 1812 2926 1829
rect 5770 1815 5786 1832
rect 2726 1774 2926 1812
rect 5728 1798 5786 1815
rect 5870 1815 5886 1832
rect 5870 1798 5928 1815
rect 5728 1760 5928 1798
rect 8368 1782 8484 1798
rect 8368 1765 8384 1782
rect 1196 1348 1396 1374
rect 1454 1348 1654 1374
rect 1712 1348 1912 1374
rect 2210 1348 2410 1374
rect 2468 1348 2668 1374
rect 2726 1348 2926 1374
rect -4922 1250 -4806 1266
rect -4922 1233 -4906 1250
rect -4964 1216 -4906 1233
rect -4822 1233 -4806 1250
rect -4296 1252 -3880 1268
rect -4296 1235 -4280 1252
rect -4822 1216 -4764 1233
rect -4964 1178 -4764 1216
rect -4488 1218 -4280 1235
rect -3896 1235 -3880 1252
rect -3324 1252 -2908 1268
rect -3324 1235 -3308 1252
rect -3896 1218 -3688 1235
rect -4488 1180 -3688 1218
rect -3516 1218 -3308 1235
rect -2924 1235 -2908 1252
rect -2388 1250 -2272 1266
rect -2924 1218 -2716 1235
rect -2388 1233 -2372 1250
rect -3516 1180 -2716 1218
rect -2430 1216 -2372 1233
rect -2288 1233 -2272 1250
rect -2288 1216 -2230 1233
rect -2430 1178 -2230 1216
rect -4964 952 -4764 978
rect -4488 954 -3688 980
rect -3516 954 -2716 980
rect -2430 952 -2230 978
rect 1609 602 1825 618
rect 1609 585 1625 602
rect 1517 568 1625 585
rect 1809 585 1825 602
rect 2204 602 2420 618
rect 2204 585 2220 602
rect 1809 568 1917 585
rect 1517 530 1917 568
rect 2112 568 2220 585
rect 2404 585 2420 602
rect 2404 568 2512 585
rect 2112 530 2512 568
rect 1517 304 1917 330
rect 2112 304 2512 330
rect 8326 1748 8384 1765
rect 8468 1765 8484 1782
rect 8468 1748 8526 1765
rect 6320 1698 6436 1714
rect 6320 1681 6336 1698
rect 6278 1664 6336 1681
rect 6420 1681 6436 1698
rect 6578 1698 6694 1714
rect 6578 1681 6594 1698
rect 6420 1664 6478 1681
rect 6278 1626 6478 1664
rect 6536 1664 6594 1681
rect 6678 1681 6694 1698
rect 6836 1698 6952 1714
rect 6836 1681 6852 1698
rect 6678 1664 6736 1681
rect 6536 1626 6736 1664
rect 6794 1664 6852 1681
rect 6936 1681 6952 1698
rect 7320 1698 7436 1714
rect 7320 1681 7336 1698
rect 6936 1664 6994 1681
rect 6794 1626 6994 1664
rect 7278 1664 7336 1681
rect 7420 1681 7436 1698
rect 7578 1698 7694 1714
rect 7578 1681 7594 1698
rect 7420 1664 7478 1681
rect 7278 1626 7478 1664
rect 7536 1664 7594 1681
rect 7678 1681 7694 1698
rect 7836 1698 7952 1714
rect 8326 1710 8526 1748
rect 7836 1681 7852 1698
rect 7678 1664 7736 1681
rect 7536 1626 7736 1664
rect 7794 1664 7852 1681
rect 7936 1681 7952 1698
rect 7936 1664 7994 1681
rect 7794 1626 7994 1664
rect 6278 800 6478 826
rect 6536 800 6736 826
rect 6794 800 6994 826
rect 7278 800 7478 826
rect 7536 800 7736 826
rect 7794 800 7994 826
rect 6320 742 6436 758
rect 6320 725 6336 742
rect 6278 708 6336 725
rect 6420 725 6436 742
rect 6578 742 6694 758
rect 6578 725 6594 742
rect 6420 708 6478 725
rect 6278 670 6478 708
rect 6536 708 6594 725
rect 6678 725 6694 742
rect 6836 742 6952 758
rect 6836 725 6852 742
rect 6678 708 6736 725
rect 6536 670 6736 708
rect 6794 708 6852 725
rect 6936 725 6952 742
rect 7320 742 7436 758
rect 7320 725 7336 742
rect 6936 708 6994 725
rect 6794 670 6994 708
rect 7278 708 7336 725
rect 7420 725 7436 742
rect 7578 742 7694 758
rect 7578 725 7594 742
rect 7420 708 7478 725
rect 7278 670 7478 708
rect 7536 708 7594 725
rect 7678 725 7694 742
rect 7836 742 7952 758
rect 7836 725 7852 742
rect 7678 708 7736 725
rect 7536 670 7736 708
rect 7794 708 7852 725
rect 7936 725 7952 742
rect 7936 708 7994 725
rect 7794 670 7994 708
rect 6278 -156 6478 -130
rect 6536 -156 6736 -130
rect 6794 -156 6994 -130
rect 7278 -156 7478 -130
rect 7536 -156 7736 -130
rect 7794 -156 7994 -130
rect 6320 -214 6436 -198
rect 6320 -231 6336 -214
rect 6278 -248 6336 -231
rect 6420 -231 6436 -214
rect 6578 -214 6694 -198
rect 6578 -231 6594 -214
rect 6420 -248 6478 -231
rect 6278 -286 6478 -248
rect 6536 -248 6594 -231
rect 6678 -231 6694 -214
rect 6836 -214 6952 -198
rect 6836 -231 6852 -214
rect 6678 -248 6736 -231
rect 6536 -286 6736 -248
rect 6794 -248 6852 -231
rect 6936 -231 6952 -214
rect 7320 -214 7436 -198
rect 7320 -231 7336 -214
rect 6936 -248 6994 -231
rect 6794 -286 6994 -248
rect 7278 -248 7336 -231
rect 7420 -231 7436 -214
rect 7578 -214 7694 -198
rect 7578 -231 7594 -214
rect 7420 -248 7478 -231
rect 7278 -286 7478 -248
rect 7536 -248 7594 -231
rect 7678 -231 7694 -214
rect 7836 -214 7952 -198
rect 7836 -231 7852 -214
rect 7678 -248 7736 -231
rect 7536 -286 7736 -248
rect 7794 -248 7852 -231
rect 7936 -231 7952 -214
rect 7936 -248 7994 -231
rect 7794 -286 7994 -248
rect 5728 -1066 5928 -1040
rect 6278 -1112 6478 -1086
rect 6536 -1112 6736 -1086
rect 6794 -1112 6994 -1086
rect 7278 -1112 7478 -1086
rect 7536 -1112 7736 -1086
rect 7794 -1112 7994 -1086
rect 8326 -1116 8526 -1090
<< polycont >>
rect -4912 4609 -4828 4643
rect -4256 4617 -4172 4651
rect -3998 4617 -3914 4651
rect -3256 4617 -3172 4651
rect -2998 4617 -2914 4651
rect -2350 4621 -2266 4655
rect -6518 3731 -6484 3765
rect -6286 3729 -6252 3763
rect -6058 3727 -6024 3761
rect -5840 3729 -5806 3763
rect 1024 4349 1108 4383
rect 1503 4341 1587 4375
rect -1332 3749 -1298 3783
rect -1100 3747 -1066 3781
rect -872 3745 -838 3779
rect -654 3747 -620 3781
rect -6518 3203 -6484 3237
rect 1761 4341 1845 4375
rect 2161 4343 2245 4377
rect 2419 4343 2503 4377
rect 2818 4323 2902 4357
rect -6286 3201 -6252 3235
rect -6058 3199 -6024 3233
rect -5840 3201 -5806 3235
rect -1332 3221 -1298 3255
rect -1100 3219 -1066 3253
rect -872 3217 -838 3251
rect 6298 4221 6382 4255
rect 6742 4203 6926 4237
rect 3844 3761 3878 3795
rect 4076 3759 4110 3793
rect 4304 3757 4338 3791
rect 4522 3759 4556 3793
rect -654 3219 -620 3253
rect 3844 3233 3878 3267
rect 4076 3231 4110 3265
rect 4304 3229 4338 3263
rect 4522 3231 4556 3265
rect 7314 4203 7498 4237
rect 7886 4233 7970 4267
rect -6494 3084 -6460 3118
rect -6278 3086 -6244 3120
rect -6060 3086 -6026 3120
rect -5838 3084 -5804 3118
rect -1308 3102 -1274 3136
rect -1092 3104 -1058 3138
rect -874 3104 -840 3138
rect -652 3102 -618 3136
rect 3868 3114 3902 3148
rect 4084 3116 4118 3150
rect 4302 3116 4336 3150
rect 9500 3553 9534 3587
rect 9732 3551 9766 3585
rect 9960 3549 9994 3583
rect 4524 3114 4558 3148
rect 10178 3551 10212 3585
rect -6494 2774 -6460 2808
rect -6278 2776 -6244 2810
rect -6060 2776 -6026 2810
rect -5838 2774 -5804 2808
rect -1308 2792 -1274 2826
rect -1092 2794 -1058 2828
rect 9500 3025 9534 3059
rect 9732 3023 9766 3057
rect 9960 3021 9994 3055
rect 10178 3023 10212 3057
rect 9524 2906 9558 2940
rect 9740 2908 9774 2942
rect 9958 2908 9992 2942
rect 10180 2906 10214 2940
rect -874 2794 -840 2828
rect -652 2792 -618 2826
rect 3868 2804 3902 2838
rect 4084 2806 4118 2840
rect 4302 2806 4336 2840
rect 4524 2804 4558 2838
rect 9524 2596 9558 2630
rect 9740 2598 9774 2632
rect 9958 2598 9992 2632
rect 10180 2596 10214 2630
rect 1262 2368 1330 2402
rect 1520 2368 1588 2402
rect 1778 2368 1846 2402
rect 2276 2368 2344 2402
rect 2534 2368 2602 2402
rect 2792 2368 2860 2402
rect 1262 1812 1330 1846
rect 1520 1812 1588 1846
rect 1778 1812 1846 1846
rect 2276 1812 2344 1846
rect 2534 1812 2602 1846
rect 2792 1812 2860 1846
rect 5786 1798 5870 1832
rect -4906 1216 -4822 1250
rect -4280 1218 -3896 1252
rect -3308 1218 -2924 1252
rect -2372 1216 -2288 1250
rect 1625 568 1809 602
rect 2220 568 2404 602
rect 8384 1748 8468 1782
rect 6336 1664 6420 1698
rect 6594 1664 6678 1698
rect 6852 1664 6936 1698
rect 7336 1664 7420 1698
rect 7594 1664 7678 1698
rect 7852 1664 7936 1698
rect 6336 708 6420 742
rect 6594 708 6678 742
rect 6852 708 6936 742
rect 7336 708 7420 742
rect 7594 708 7678 742
rect 7852 708 7936 742
rect 6336 -248 6420 -214
rect 6594 -248 6678 -214
rect 6852 -248 6936 -214
rect 7336 -248 7420 -214
rect 7594 -248 7678 -214
rect 7852 -248 7936 -214
<< xpolycontact >>
rect -7512 9378 -7080 9448
rect -3230 9378 -2798 9448
rect -2282 9378 -1850 9448
rect 2000 9378 2432 9448
rect 2948 9378 3380 9448
rect 7230 9378 7662 9448
rect 8178 9378 8610 9448
rect 12460 9378 12892 9448
rect -7512 9058 -7080 9128
rect -3230 9058 -2798 9128
rect -2282 9058 -1850 9128
rect 2000 9058 2432 9128
rect 2948 9058 3380 9128
rect 7230 9058 7662 9128
rect 8178 9058 8610 9128
rect 12460 9058 12892 9128
rect -7512 8738 -7080 8808
rect -3230 8738 -2798 8808
rect -2268 8716 -1836 8786
rect 2014 8716 2446 8786
rect 2928 8718 3360 8788
rect 7210 8718 7642 8788
rect 8178 8738 8610 8808
rect 12460 8738 12892 8808
rect -7512 8418 -7080 8488
rect -3230 8418 -2798 8488
rect -2268 8398 -1836 8468
rect 2014 8398 2446 8468
rect 2928 8400 3360 8470
rect 7210 8400 7642 8470
rect 8178 8418 8610 8488
rect 12460 8418 12892 8488
rect -7512 8098 -7080 8168
rect -3230 8098 -2798 8168
rect -2268 8080 -1836 8150
rect 2014 8080 2446 8150
rect 2928 8082 3360 8152
rect 7210 8082 7642 8152
rect 8178 8098 8610 8168
rect 12460 8098 12892 8168
rect -7512 7778 -7080 7848
rect -3230 7778 -2798 7848
rect -2268 7762 -1836 7832
rect 2014 7762 2446 7832
rect 2928 7764 3360 7834
rect 7210 7764 7642 7834
rect 8178 7778 8610 7848
rect 12460 7778 12892 7848
rect -7512 7458 -7080 7528
rect -3230 7458 -2798 7528
rect -2268 7444 -1836 7514
rect 2014 7444 2446 7514
rect 2928 7446 3360 7516
rect 7210 7446 7642 7516
rect 8178 7458 8610 7528
rect 12460 7458 12892 7528
rect -7512 7138 -7080 7208
rect -3230 7138 -2798 7208
rect -2268 7126 -1836 7196
rect 2014 7126 2446 7196
rect 2928 7128 3360 7198
rect 7210 7128 7642 7198
rect 8178 7138 8610 7208
rect 12460 7138 12892 7208
rect -7512 6818 -7080 6888
rect -3230 6818 -2798 6888
rect -2268 6808 -1836 6878
rect 2014 6808 2446 6878
rect 2928 6810 3360 6880
rect 7210 6810 7642 6880
rect 8178 6818 8610 6888
rect 12460 6818 12892 6888
rect -7512 6498 -7080 6568
rect -3230 6498 -2798 6568
rect -2268 6490 -1836 6560
rect 2014 6490 2446 6560
rect 2928 6492 3360 6562
rect 7210 6492 7642 6562
rect 8178 6498 8610 6568
rect 12460 6498 12892 6568
rect -7512 6178 -7080 6248
rect -3230 6178 -2798 6248
rect -2268 6172 -1836 6242
rect 2014 6172 2446 6242
rect 2928 6174 3360 6244
rect 7210 6174 7642 6244
rect 8178 6178 8610 6248
rect 12460 6178 12892 6248
rect -7512 5858 -7080 5928
rect -3230 5858 -2798 5928
rect -2248 5826 -1816 5896
rect 2034 5826 2466 5896
rect 2948 5856 3380 5926
rect 7230 5856 7662 5926
rect 8178 5858 8610 5928
rect 12460 5858 12892 5928
rect -7512 5538 -7080 5608
rect -3230 5538 -2798 5608
rect -2248 5506 -1816 5576
rect 2034 5506 2466 5576
rect 2948 5538 3380 5608
rect 7230 5538 7662 5608
rect 8178 5538 8610 5608
rect 12460 5538 12892 5608
<< xpolyres >>
rect -7080 9378 -3230 9448
rect -1850 9378 2000 9448
rect 3380 9378 7230 9448
rect 8610 9378 12460 9448
rect -7080 9058 -3230 9128
rect -1850 9058 2000 9128
rect 3380 9058 7230 9128
rect 8610 9058 12460 9128
rect -7080 8738 -3230 8808
rect -1836 8716 2014 8786
rect 3360 8718 7210 8788
rect 8610 8738 12460 8808
rect -7080 8418 -3230 8488
rect -1836 8398 2014 8468
rect 3360 8400 7210 8470
rect 8610 8418 12460 8488
rect -7080 8098 -3230 8168
rect -1836 8080 2014 8150
rect 3360 8082 7210 8152
rect 8610 8098 12460 8168
rect -7080 7778 -3230 7848
rect -1836 7762 2014 7832
rect 3360 7764 7210 7834
rect 8610 7778 12460 7848
rect -7080 7458 -3230 7528
rect -1836 7444 2014 7514
rect 3360 7446 7210 7516
rect 8610 7458 12460 7528
rect -7080 7138 -3230 7208
rect -1836 7126 2014 7196
rect 3360 7128 7210 7198
rect 8610 7138 12460 7208
rect -7080 6818 -3230 6888
rect -1836 6808 2014 6878
rect 3360 6810 7210 6880
rect 8610 6818 12460 6888
rect -7080 6498 -3230 6568
rect -1836 6490 2014 6560
rect 3360 6492 7210 6562
rect 8610 6498 12460 6568
rect -7080 6178 -3230 6248
rect -1836 6172 2014 6242
rect 3360 6174 7210 6244
rect 8610 6178 12460 6248
rect -7080 5858 -3230 5928
rect -1816 5826 2034 5896
rect 3380 5856 7230 5926
rect 8610 5858 12460 5928
rect -7080 5538 -3230 5608
rect -1816 5506 2034 5576
rect 3380 5538 7230 5608
rect 8610 5538 12460 5608
<< locali >>
rect 10156 10714 11468 10908
rect 10156 10220 10364 10714
rect 11324 10220 11468 10714
rect 10156 10000 11468 10220
rect -7520 9448 -7076 9458
rect -2290 9448 -1846 9458
rect 2940 9448 3384 9458
rect 8170 9448 8614 9458
rect -7520 9378 -7512 9448
rect -7080 9378 -7076 9448
rect -2290 9378 -2282 9448
rect -1850 9378 -1846 9448
rect 2940 9378 2948 9448
rect 3380 9378 3384 9448
rect 8170 9378 8178 9448
rect 8610 9378 8614 9448
rect -7520 9366 -7076 9378
rect -2290 9366 -1846 9378
rect 2940 9366 3384 9378
rect 8170 9366 8614 9378
rect -7520 9128 -7076 9138
rect -2290 9128 -1846 9138
rect 2940 9128 3384 9138
rect 8170 9128 8614 9138
rect -7520 9058 -7512 9128
rect -7080 9058 -7076 9128
rect -2290 9058 -2282 9128
rect -1850 9058 -1846 9128
rect 2940 9058 2948 9128
rect 3380 9058 3384 9128
rect 8170 9058 8178 9128
rect 8610 9058 8614 9128
rect -7520 9046 -7076 9058
rect -2290 9046 -1846 9058
rect 2940 9046 3384 9058
rect 8170 9046 8614 9058
rect -7520 8808 -7076 8818
rect 8170 8808 8614 8818
rect -7520 8738 -7512 8808
rect -7080 8738 -7076 8808
rect -7520 8726 -7076 8738
rect 8170 8738 8178 8808
rect 8610 8738 8614 8808
rect 8170 8726 8614 8738
rect -7520 8488 -7076 8498
rect 8170 8488 8614 8498
rect -7520 8418 -7512 8488
rect -7080 8418 -7076 8488
rect -7520 8406 -7076 8418
rect 8170 8418 8178 8488
rect 8610 8418 8614 8488
rect 8170 8406 8614 8418
rect -7520 8168 -7076 8178
rect 8170 8168 8614 8178
rect -7520 8098 -7512 8168
rect -7080 8098 -7076 8168
rect -7520 8086 -7076 8098
rect 8170 8098 8178 8168
rect 8610 8098 8614 8168
rect 8170 8086 8614 8098
rect -7520 7848 -7076 7858
rect 8170 7848 8614 7858
rect -7520 7778 -7512 7848
rect -7080 7778 -7076 7848
rect -7520 7766 -7076 7778
rect 8170 7778 8178 7848
rect 8610 7778 8614 7848
rect 8170 7766 8614 7778
rect -7520 7528 -7076 7538
rect 8170 7528 8614 7538
rect -7520 7458 -7512 7528
rect -7080 7458 -7076 7528
rect -7520 7446 -7076 7458
rect 8170 7458 8178 7528
rect 8610 7458 8614 7528
rect 8170 7446 8614 7458
rect -7520 7208 -7076 7218
rect 8170 7208 8614 7218
rect -7520 7138 -7512 7208
rect -7080 7138 -7076 7208
rect -7520 7126 -7076 7138
rect 8170 7138 8178 7208
rect 8610 7138 8614 7208
rect 8170 7126 8614 7138
rect -7520 6888 -7076 6898
rect 8170 6888 8614 6898
rect -7520 6818 -7512 6888
rect -7080 6818 -7076 6888
rect -7520 6806 -7076 6818
rect 8170 6818 8178 6888
rect 8610 6818 8614 6888
rect 8170 6806 8614 6818
rect -7520 6568 -7076 6578
rect 8170 6568 8614 6578
rect -7520 6498 -7512 6568
rect -7080 6498 -7076 6568
rect -7520 6486 -7076 6498
rect 8170 6498 8178 6568
rect 8610 6498 8614 6568
rect 8170 6486 8614 6498
rect -7520 6248 -7076 6258
rect 8170 6248 8614 6258
rect -7520 6178 -7512 6248
rect -7080 6178 -7076 6248
rect -7520 6166 -7076 6178
rect 8170 6178 8178 6248
rect 8610 6178 8614 6248
rect 8170 6166 8614 6178
rect -7520 5928 -7076 5938
rect -7520 5858 -7512 5928
rect -7080 5858 -7076 5928
rect 2940 5926 3384 5936
rect 8170 5928 8614 5938
rect -2256 5896 -1812 5906
rect -7520 5846 -7076 5858
rect -2256 5826 -2248 5896
rect -1816 5826 -1812 5896
rect 2940 5856 2948 5926
rect 3380 5856 3384 5926
rect 8170 5858 8178 5928
rect 8610 5858 8614 5928
rect 2940 5844 3384 5856
rect 8170 5846 8614 5858
rect -2256 5814 -1812 5826
rect -7520 5608 -7076 5618
rect 2940 5608 3384 5618
rect 8170 5608 8614 5618
rect -7520 5538 -7512 5608
rect -7080 5538 -7076 5608
rect -2256 5576 -1812 5586
rect -7520 5526 -7076 5538
rect -2256 5506 -2248 5576
rect -1816 5506 -1812 5576
rect 2940 5538 2948 5608
rect 3380 5538 3384 5608
rect 8170 5538 8178 5608
rect 8610 5538 8614 5608
rect 2940 5526 3384 5538
rect 8170 5526 8614 5538
rect -2256 5494 -1812 5506
rect -1802 5088 -312 5094
rect -4124 5052 -312 5088
rect -4124 5050 -1748 5052
rect -6356 4662 -5842 4758
rect -4116 4680 -4078 5050
rect -1770 5012 -1726 5014
rect -3102 4974 -1726 5012
rect 2662 5098 2780 5124
rect -18 5052 58 5072
rect -3102 4680 -3064 4974
rect -6356 4422 -6262 4662
rect -5936 4422 -5842 4662
rect -4286 4651 -3876 4680
rect -4928 4609 -4912 4643
rect -4828 4609 -4812 4643
rect -4286 4617 -4256 4651
rect -4172 4617 -3998 4651
rect -3914 4617 -3876 4651
rect -3278 4651 -2868 4680
rect -4286 4606 -3876 4617
rect -3278 4617 -3256 4651
rect -3172 4617 -2998 4651
rect -2914 4617 -2868 4651
rect -2366 4621 -2350 4655
rect -2266 4621 -2250 4655
rect -3278 4606 -2868 4617
rect -3678 4522 -3610 4554
rect -6356 4324 -5842 4422
rect -4494 4478 -4066 4480
rect -4494 4414 -4064 4478
rect -5016 4306 -4982 4322
rect -6710 3834 -6482 3846
rect -6710 3810 -6018 3834
rect -6518 3800 -6018 3810
rect -5016 3802 -4982 3818
rect -4758 4306 -4724 4322
rect -4758 3802 -4724 3818
rect -6518 3765 -6462 3800
rect -6534 3731 -6518 3765
rect -6484 3760 -6462 3765
rect -6072 3782 -6018 3800
rect -6484 3731 -6468 3760
rect -6302 3729 -6286 3763
rect -6252 3729 -6236 3763
rect -6072 3761 -6008 3782
rect -6074 3727 -6058 3761
rect -6024 3727 -6008 3761
rect -5856 3729 -5840 3763
rect -5806 3729 -5790 3763
rect -6062 3724 -6020 3727
rect -6526 3237 -6478 3240
rect -6534 3203 -6518 3237
rect -6484 3203 -6468 3237
rect -6390 3235 -6246 3242
rect -6168 3240 -6106 3242
rect -6526 3172 -6478 3203
rect -6390 3202 -6286 3235
rect -6706 3124 -6436 3126
rect -6390 3124 -6354 3202
rect -6302 3201 -6286 3202
rect -6252 3201 -6236 3235
rect -6168 3233 -6018 3240
rect -5942 3235 -5804 3238
rect -6706 3118 -6354 3124
rect -6168 3199 -6058 3233
rect -6024 3199 -6008 3233
rect -5942 3201 -5840 3235
rect -5806 3201 -5790 3235
rect -5942 3200 -5804 3201
rect -6168 3190 -6018 3199
rect -6168 3176 -6106 3190
rect -6168 3120 -6130 3176
rect -5942 3120 -5906 3200
rect -6706 3084 -6494 3118
rect -6460 3084 -6354 3118
rect -6294 3086 -6278 3120
rect -6244 3086 -6130 3120
rect -6076 3086 -6060 3120
rect -6026 3086 -5906 3120
rect -5854 3084 -5838 3118
rect -5804 3084 -5788 3118
rect -6706 3080 -6436 3084
rect -4492 3004 -4450 4414
rect -4108 4402 -4064 4414
rect -4106 4380 -4064 4402
rect -3676 4402 -3610 4522
rect -4360 4314 -4326 4330
rect -4370 3826 -4360 3884
rect -4106 4314 -4062 4380
rect -4106 4290 -4102 4314
rect -4326 3826 -4318 3884
rect -4370 3694 -4318 3826
rect -4068 4290 -4062 4314
rect -3844 4314 -3810 4330
rect -4102 3810 -4068 3826
rect -3852 3826 -3844 3880
rect -3810 3826 -3800 3880
rect -3852 3706 -3800 3826
rect -3676 3706 -3614 4402
rect -3108 4378 -2670 4478
rect -3360 4314 -3326 4330
rect -4038 3694 -3614 3706
rect -4370 3686 -3614 3694
rect -3366 3826 -3360 3848
rect -3106 4314 -3062 4378
rect -3106 4292 -3102 4314
rect -3326 3826 -3320 3848
rect -3366 3716 -3320 3826
rect -3068 4292 -3062 4314
rect -2844 4314 -2810 4330
rect -3102 3810 -3068 3826
rect -2850 3826 -2844 3860
rect -2810 3826 -2804 3860
rect -2850 3716 -2804 3826
rect -3366 3686 -2804 3716
rect -4370 3622 -2804 3686
rect -4370 3620 -3798 3622
rect -3692 3620 -2804 3622
rect -4122 3618 -4048 3620
rect -3852 3618 -3800 3620
rect -3366 3618 -2804 3620
rect -3362 3610 -2804 3618
rect -2708 3340 -2670 4378
rect -2454 4318 -2420 4334
rect -2454 3814 -2420 3830
rect -2196 4318 -2162 4334
rect -2196 3814 -2162 3830
rect -2734 3304 -2668 3340
rect -4492 2966 -3642 3004
rect -6240 2814 -6150 2818
rect -6494 2808 -6458 2812
rect -6240 2810 -6210 2814
rect -6510 2774 -6494 2808
rect -6460 2774 -6444 2808
rect -6294 2776 -6278 2810
rect -6244 2776 -6210 2810
rect -6170 2776 -6150 2814
rect -6076 2810 -6010 2812
rect -6076 2776 -6060 2810
rect -6026 2776 -6010 2810
rect -5942 2810 -5854 2818
rect -5942 2776 -5932 2810
rect -5898 2808 -5854 2810
rect -5898 2776 -5838 2808
rect -6494 2738 -6458 2774
rect -6240 2772 -6150 2776
rect -6058 2738 -6024 2776
rect -5942 2774 -5838 2776
rect -5804 2774 -5788 2808
rect -5942 2772 -5854 2774
rect -5942 2766 -5886 2772
rect -6494 2698 -6024 2738
rect -3686 2828 -3646 2966
rect -3774 2780 -3640 2828
rect -3686 2082 -3646 2780
rect -2712 2550 -2668 3304
rect -1770 2672 -1726 4974
rect -18 4952 -6 5052
rect 46 4952 58 5052
rect -18 4932 58 4952
rect 158 5048 244 5072
rect 158 4964 174 5048
rect 226 4964 244 5048
rect 158 4940 244 4964
rect 886 5070 986 5090
rect 886 4972 898 5070
rect 976 4972 986 5070
rect 886 4940 986 4972
rect 2662 4966 2676 5098
rect 2764 4966 2780 5098
rect 2662 4946 2780 4966
rect -1468 4740 -954 4836
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect -1468 4402 -954 4500
rect -1508 3852 -1286 3860
rect -1508 3824 -832 3852
rect -1332 3818 -832 3824
rect -1332 3783 -1276 3818
rect -1348 3749 -1332 3783
rect -1298 3778 -1276 3783
rect -886 3800 -832 3818
rect -1298 3749 -1282 3778
rect -1116 3747 -1100 3781
rect -1066 3747 -1050 3781
rect -886 3779 -822 3800
rect -888 3745 -872 3779
rect -838 3745 -822 3779
rect -670 3747 -654 3781
rect -620 3747 -604 3781
rect -876 3742 -834 3745
rect -1340 3255 -1292 3258
rect -1348 3221 -1332 3255
rect -1298 3221 -1282 3255
rect -1204 3253 -1060 3260
rect -982 3258 -920 3260
rect -1340 3190 -1292 3221
rect -1204 3220 -1100 3253
rect -1204 3144 -1168 3220
rect -1116 3219 -1100 3220
rect -1066 3219 -1050 3253
rect -982 3251 -832 3258
rect -756 3253 -618 3256
rect -1498 3136 -1168 3144
rect -982 3217 -872 3251
rect -838 3217 -822 3251
rect -756 3219 -654 3253
rect -620 3219 -604 3253
rect -756 3218 -618 3219
rect -982 3208 -832 3217
rect -982 3194 -920 3208
rect -982 3138 -944 3194
rect -756 3138 -720 3218
rect -1498 3102 -1308 3136
rect -1274 3102 -1168 3136
rect -1108 3104 -1092 3138
rect -1058 3104 -944 3138
rect -890 3104 -874 3138
rect -840 3104 -720 3138
rect -668 3102 -652 3136
rect -618 3102 -602 3136
rect -1498 3098 -1196 3102
rect -1054 2832 -964 2836
rect -1308 2826 -1272 2830
rect -1054 2828 -1024 2832
rect -1324 2792 -1308 2826
rect -1274 2792 -1258 2826
rect -1108 2794 -1092 2828
rect -1058 2794 -1024 2828
rect -984 2794 -964 2832
rect -890 2828 -824 2830
rect -890 2794 -874 2828
rect -840 2794 -824 2828
rect -756 2828 -668 2836
rect -756 2794 -746 2828
rect -712 2826 -668 2828
rect -712 2794 -652 2826
rect -1308 2756 -1272 2792
rect -1054 2790 -964 2794
rect -872 2756 -838 2794
rect -756 2792 -652 2794
rect -618 2792 -602 2826
rect -756 2790 -668 2792
rect -756 2784 -700 2790
rect -1308 2716 -838 2756
rect -1770 2602 -1726 2604
rect -2760 2502 -2662 2550
rect -3688 2034 -3644 2082
rect -2712 2064 -2668 2502
rect -3686 1482 -3646 2034
rect -2714 2004 -2666 2064
rect -2712 1482 -2668 2004
rect -3686 1396 -3638 1482
rect -2712 1444 -2664 1482
rect -3682 1366 -3638 1396
rect -4922 1216 -4906 1250
rect -4822 1216 -4806 1250
rect -4296 1218 -4280 1252
rect -3896 1218 -3880 1252
rect -5010 1122 -4976 1138
rect -5010 1018 -4976 1034
rect -4752 1122 -4718 1138
rect -4752 1018 -4718 1034
rect -4534 1124 -4500 1140
rect -4534 1020 -4500 1036
rect -3678 1124 -3640 1366
rect -2706 1362 -2664 1444
rect -3324 1218 -3308 1252
rect -2924 1218 -2908 1252
rect -3678 1036 -3676 1124
rect -3642 1036 -3640 1124
rect -3678 1010 -3640 1036
rect -3562 1124 -3528 1140
rect -3562 1020 -3528 1036
rect -2704 1124 -2666 1362
rect -2388 1216 -2372 1250
rect -2288 1216 -2272 1250
rect -2670 1036 -2666 1124
rect -2704 1016 -2666 1036
rect -2476 1122 -2442 1138
rect -2476 1018 -2442 1034
rect -2218 1122 -2184 1138
rect -2218 1018 -2184 1034
rect -4320 344 -3008 538
rect -4320 -150 -4112 344
rect -3152 -150 -3008 344
rect 0 40 44 4932
rect 176 276 218 4940
rect 908 4498 976 4940
rect 908 4046 968 4498
rect 1648 4404 1702 4574
rect 2094 4406 2164 4408
rect 2312 4406 2370 4634
rect 2692 4524 2760 4946
rect 5128 4838 5236 4850
rect 5128 4752 5142 4838
rect 5224 4752 5236 4838
rect 5128 4734 5236 4752
rect 6560 4820 6658 4826
rect 6560 4766 6582 4820
rect 6642 4766 6658 4820
rect 6560 4750 6658 4766
rect 7032 4750 7096 4760
rect 3844 4528 4358 4624
rect 1008 4349 1024 4383
rect 1108 4349 1124 4383
rect 1497 4375 1972 4404
rect 1487 4341 1503 4375
rect 1587 4341 1761 4375
rect 1845 4341 1972 4375
rect 1497 4332 1972 4341
rect 2094 4377 2652 4406
rect 2094 4343 2161 4377
rect 2245 4343 2419 4377
rect 2503 4343 2652 4377
rect 2094 4336 2652 4343
rect 2155 4334 2652 4336
rect 908 3558 920 4046
rect 954 3558 968 4046
rect 908 3546 968 3558
rect 1162 4046 1218 4066
rect 1661 4054 1695 4110
rect 1162 3558 1178 4046
rect 1212 3558 1218 4046
rect 920 3542 954 3546
rect 1162 3230 1218 3558
rect 1657 4038 1695 4054
rect 1915 4052 1949 4054
rect 1654 3550 1657 3626
rect 1691 3744 1695 4038
rect 1911 4038 1953 4052
rect 1691 3550 1700 3626
rect 1399 3534 1433 3540
rect 1654 3204 1700 3550
rect 1911 3544 1915 4038
rect 1949 3544 1953 4038
rect 2319 4056 2353 4082
rect 2315 4040 2353 4056
rect 2309 3686 2315 3810
rect 2349 3810 2353 4040
rect 2573 4040 2607 4056
rect 2349 3686 2355 3810
rect 2309 3656 2355 3686
rect 1911 3304 1953 3544
rect 2057 3536 2091 3546
rect 1906 3024 1954 3304
rect 2312 3192 2352 3656
rect 2566 3546 2573 3610
rect 2566 3536 2607 3546
rect 2698 4020 2750 4524
rect 2802 4323 2818 4357
rect 2902 4323 2918 4357
rect 3844 4288 3938 4528
rect 4264 4288 4358 4528
rect 3844 4190 4358 4288
rect 2972 4034 3006 4036
rect 2566 3264 2605 3536
rect 2698 3532 2714 4020
rect 2748 3532 2750 4020
rect 2698 3524 2750 3532
rect 2962 4020 3014 4034
rect 2962 3532 2972 4020
rect 3006 3532 3014 4020
rect 3298 3938 3474 3970
rect 3298 3862 3328 3938
rect 3438 3862 3474 3938
rect 3298 3820 3474 3862
rect 3772 3830 4344 3864
rect 2714 3516 2748 3524
rect 2566 3262 2608 3264
rect 1896 2914 1954 3024
rect 1896 2644 1948 2914
rect 878 2604 1948 2644
rect 882 2586 1948 2604
rect 2308 2646 2356 3192
rect 2564 3012 2610 3262
rect 2962 3162 3014 3532
rect 3346 3536 3386 3820
rect 3844 3795 3900 3830
rect 3828 3761 3844 3795
rect 3878 3790 3900 3795
rect 4290 3812 4344 3830
rect 3878 3761 3894 3790
rect 4060 3759 4076 3793
rect 4110 3759 4126 3793
rect 4290 3791 4354 3812
rect 4288 3757 4304 3791
rect 4338 3757 4354 3791
rect 4506 3759 4522 3793
rect 4556 3759 4572 3793
rect 4300 3754 4342 3757
rect 3346 3496 3754 3536
rect 2608 2972 2610 3012
rect 2960 2910 3014 3162
rect 3544 3222 3660 3236
rect 3544 3152 3562 3222
rect 3638 3152 3660 3222
rect 3544 3134 3660 3152
rect 2308 2608 2612 2646
rect 882 2560 940 2586
rect 2308 2578 2878 2608
rect 2308 2576 2356 2578
rect 878 2546 940 2560
rect 2564 2554 2878 2578
rect 878 2429 948 2546
rect 1518 2430 1596 2438
rect 2532 2430 2610 2438
rect 859 2411 972 2429
rect 1518 2428 1604 2430
rect 2012 2428 2048 2430
rect 2532 2428 2618 2430
rect 859 2310 869 2411
rect 969 2310 972 2411
rect 1250 2402 2056 2428
rect 2264 2416 3016 2428
rect 3076 2416 3252 2432
rect 2264 2414 3252 2416
rect 2264 2402 3102 2414
rect 1246 2368 1262 2402
rect 1330 2368 1520 2402
rect 1588 2368 1778 2402
rect 1846 2368 2056 2402
rect 2260 2368 2276 2402
rect 2344 2368 2534 2402
rect 2602 2368 2792 2402
rect 2860 2368 3102 2402
rect 859 2291 972 2310
rect 1250 2362 2056 2368
rect 2264 2362 3102 2368
rect 3226 2362 3252 2414
rect 888 1226 942 2291
rect 1139 2205 1191 2242
rect 1139 2055 1150 2205
rect 1184 2055 1191 2205
rect 1139 1950 1191 2055
rect 1146 1660 1190 1950
rect 1250 1846 1336 2362
rect 1408 2220 1442 2221
rect 1518 1846 1604 2362
rect 1246 1812 1262 1846
rect 1330 1812 1346 1846
rect 1504 1812 1520 1846
rect 1588 1812 1604 1846
rect 1250 1798 1336 1812
rect 1518 1808 1604 1812
rect 1660 2205 1704 2230
rect 1660 2055 1666 2205
rect 1700 2055 1704 2205
rect 1142 1649 1190 1660
rect 1142 1499 1150 1649
rect 1184 1499 1190 1649
rect 1142 1480 1190 1499
rect 1660 1649 1704 2055
rect 1776 1846 1862 2362
rect 1924 2039 1958 2044
rect 1762 1812 1778 1846
rect 1846 1812 1862 1846
rect 1776 1806 1862 1812
rect 1660 1624 1666 1649
rect 1656 1499 1666 1624
rect 1700 1499 1704 1649
rect 1656 1490 1704 1499
rect 1142 1392 1186 1480
rect 1656 1392 1700 1490
rect 1924 1483 1958 1488
rect 1140 1314 1704 1392
rect 888 1214 954 1226
rect 888 1174 902 1214
rect 944 1174 954 1214
rect 888 1162 954 1174
rect 1534 1036 1574 1314
rect 2012 1246 2048 2362
rect 2153 2205 2205 2242
rect 2153 2055 2164 2205
rect 2198 2055 2205 2205
rect 2153 1950 2205 2055
rect 2160 1660 2204 1950
rect 2264 1846 2350 2362
rect 2422 2220 2456 2221
rect 2532 1846 2618 2362
rect 2260 1812 2276 1846
rect 2344 1812 2360 1846
rect 2518 1812 2534 1846
rect 2602 1812 2618 1846
rect 2264 1798 2350 1812
rect 2532 1808 2618 1812
rect 2674 2205 2718 2230
rect 2674 2055 2680 2205
rect 2714 2055 2718 2205
rect 2156 1649 2204 1660
rect 2156 1499 2164 1649
rect 2198 1499 2204 1649
rect 2156 1480 2204 1499
rect 2674 1649 2718 2055
rect 2790 1846 2876 2362
rect 3076 2344 3252 2362
rect 2938 2039 2972 2044
rect 2776 1812 2792 1846
rect 2860 1812 2876 1846
rect 2790 1806 2876 1812
rect 2674 1624 2680 1649
rect 2670 1499 2680 1624
rect 2714 1499 2718 1649
rect 2670 1490 2718 1499
rect 2156 1392 2200 1480
rect 2670 1392 2714 1490
rect 2938 1483 2972 1488
rect 2154 1326 2718 1392
rect 2154 1314 2808 1326
rect 2548 1290 2808 1314
rect 2764 1158 2808 1290
rect 2764 1156 3188 1158
rect 2764 1114 3316 1156
rect 3136 1112 3316 1114
rect 3558 1036 3594 3134
rect 1534 998 3594 1036
rect 3696 1984 3730 3496
rect 3836 3267 3884 3270
rect 3828 3233 3844 3267
rect 3878 3233 3894 3267
rect 3972 3265 4116 3272
rect 4194 3270 4256 3272
rect 3836 3202 3884 3233
rect 3972 3232 4076 3265
rect 3972 3154 4008 3232
rect 4060 3231 4076 3232
rect 4110 3231 4126 3265
rect 4194 3263 4344 3270
rect 4420 3265 4558 3268
rect 3780 3148 4008 3154
rect 4194 3229 4304 3263
rect 4338 3229 4354 3263
rect 4420 3231 4522 3265
rect 4556 3231 4572 3265
rect 4420 3230 4558 3231
rect 4194 3220 4344 3229
rect 4194 3206 4256 3220
rect 4194 3150 4232 3206
rect 4420 3150 4456 3230
rect 3780 3114 3868 3148
rect 3902 3114 4008 3148
rect 4068 3116 4084 3150
rect 4118 3116 4232 3150
rect 4286 3116 4302 3150
rect 4336 3116 4456 3150
rect 4508 3114 4524 3148
rect 4558 3114 4574 3148
rect 3780 3108 3922 3114
rect 4122 2844 4212 2848
rect 3868 2838 3904 2842
rect 4122 2840 4152 2844
rect 3852 2804 3868 2838
rect 3902 2804 3918 2838
rect 4068 2806 4084 2840
rect 4118 2806 4152 2840
rect 4192 2806 4212 2844
rect 4286 2840 4352 2842
rect 4286 2806 4302 2840
rect 4336 2806 4352 2840
rect 4420 2840 4508 2848
rect 4420 2806 4430 2840
rect 4464 2838 4508 2840
rect 4464 2806 4524 2838
rect 3868 2768 3904 2804
rect 4122 2802 4212 2806
rect 4304 2768 4338 2806
rect 4420 2804 4524 2806
rect 4558 2804 4574 2838
rect 4420 2802 4508 2804
rect 4420 2796 4476 2802
rect 3868 2728 4338 2768
rect 3696 1938 5050 1984
rect 3696 936 3730 1938
rect 1918 888 3730 936
rect 1918 632 1974 888
rect 3126 820 4672 828
rect 2522 774 4672 820
rect 2522 632 2576 774
rect 3126 772 4672 774
rect 1599 623 1884 625
rect 1508 606 1884 623
rect 1508 566 1612 606
rect 1810 566 1884 606
rect 1508 561 1884 566
rect 1599 555 1884 561
rect 1918 542 1972 632
rect 2205 604 2426 625
rect 2205 602 2223 604
rect 2204 568 2220 602
rect 2205 566 2223 568
rect 2205 555 2426 566
rect 1471 487 1505 490
rect 1459 479 1505 487
rect 1459 474 1509 479
rect 1459 386 1471 474
rect 1505 386 1509 474
rect 1459 360 1509 386
rect 1926 474 1971 542
rect 1926 386 1929 474
rect 1963 386 1971 474
rect 1926 379 1971 386
rect 2049 480 2101 493
rect 2527 490 2567 632
rect 2049 474 2112 480
rect 2049 386 2066 474
rect 2100 386 2112 474
rect 1929 370 1963 379
rect 1470 276 1509 360
rect 2049 369 2112 386
rect 2524 474 2567 490
rect 2558 386 2567 474
rect 2524 384 2567 386
rect 2524 370 2558 384
rect 2049 276 2101 369
rect 176 230 1512 276
rect 1470 226 1509 230
rect 2050 40 2100 276
rect 0 0 2100 40
rect 3102 160 4414 354
rect -4320 -370 -3008 -150
rect 3102 -334 3310 160
rect 4270 -334 4414 160
rect 3102 -554 4414 -334
rect 5164 -1308 5206 4734
rect 6282 4221 6298 4255
rect 6382 4221 6398 4255
rect 6580 4030 6630 4750
rect 7026 4716 8618 4750
rect 6726 4203 6742 4237
rect 6926 4203 6942 4237
rect 6194 3918 6228 3934
rect 6194 3414 6228 3430
rect 6452 3918 6486 3934
rect 6580 3900 6628 4030
rect 6580 3860 6588 3900
rect 6452 3414 6486 3430
rect 6622 3860 6628 3900
rect 7032 3900 7096 4716
rect 7654 4644 8708 4648
rect 7602 4608 8708 4644
rect 7150 3998 7200 4430
rect 7298 4203 7314 4237
rect 7498 4203 7514 4237
rect 7032 3862 7046 3900
rect 6588 3396 6622 3412
rect 7014 3412 7046 3470
rect 7080 3862 7096 3900
rect 7152 3900 7200 3998
rect 7152 3862 7160 3900
rect 7080 3412 7100 3470
rect 7014 3048 7100 3412
rect 7194 3862 7200 3900
rect 7602 3900 7666 4608
rect 9280 4470 9794 4566
rect 7870 4233 7886 4267
rect 7970 4233 7986 4267
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
rect 7602 3872 7618 3900
rect 7160 3396 7194 3412
rect 7588 3412 7618 3450
rect 7652 3872 7666 3900
rect 7782 3930 7816 3946
rect 7652 3412 7690 3450
rect 7782 3426 7816 3442
rect 8040 3930 8074 3946
rect 9400 3656 9538 3662
rect 9400 3626 10000 3656
rect 9500 3622 10000 3626
rect 9500 3587 9556 3622
rect 9484 3553 9500 3587
rect 9534 3582 9556 3587
rect 9946 3604 10000 3622
rect 9534 3553 9550 3582
rect 9716 3551 9732 3585
rect 9766 3551 9782 3585
rect 9946 3583 10010 3604
rect 9944 3549 9960 3583
rect 9994 3549 10010 3583
rect 10162 3551 10178 3585
rect 10212 3551 10228 3585
rect 9956 3546 9998 3549
rect 8040 3426 8074 3442
rect 7588 3058 7690 3412
rect 9492 3059 9540 3062
rect 7014 3040 7076 3048
rect 6988 2704 7076 3040
rect 7588 3036 7672 3058
rect 6982 2590 7082 2704
rect 7586 2694 7672 3036
rect 9484 3025 9500 3059
rect 9534 3025 9550 3059
rect 9628 3057 9772 3064
rect 9850 3062 9912 3064
rect 9492 2994 9540 3025
rect 9628 3024 9732 3057
rect 9628 2946 9664 3024
rect 9716 3023 9732 3024
rect 9766 3023 9782 3057
rect 9850 3055 10000 3062
rect 10076 3057 10214 3060
rect 9340 2940 9664 2946
rect 9850 3021 9960 3055
rect 9994 3021 10010 3055
rect 10076 3023 10178 3057
rect 10212 3023 10228 3057
rect 10076 3022 10214 3023
rect 9850 3012 10000 3021
rect 9850 2998 9912 3012
rect 9850 2942 9888 2998
rect 10076 2942 10112 3022
rect 9340 2906 9524 2940
rect 9558 2906 9664 2940
rect 9724 2908 9740 2942
rect 9774 2908 9888 2942
rect 9942 2908 9958 2942
rect 9992 2908 10112 2942
rect 10164 2906 10180 2940
rect 10214 2906 10230 2940
rect 7578 2604 7696 2694
rect 9778 2636 9868 2640
rect 9524 2630 9560 2634
rect 9778 2632 9808 2636
rect 6988 2002 7076 2590
rect 6992 2000 7076 2002
rect 7586 2036 7672 2604
rect 9508 2596 9524 2630
rect 9558 2596 9574 2630
rect 9724 2598 9740 2632
rect 9774 2598 9808 2632
rect 9848 2598 9868 2636
rect 9942 2632 10008 2634
rect 9942 2598 9958 2632
rect 9992 2598 10008 2632
rect 10076 2632 10164 2640
rect 10076 2598 10086 2632
rect 10120 2630 10164 2632
rect 10120 2598 10180 2630
rect 9524 2560 9560 2596
rect 9778 2594 9868 2598
rect 9960 2560 9994 2598
rect 10076 2596 10180 2598
rect 10214 2596 10230 2630
rect 10076 2594 10164 2596
rect 10076 2588 10132 2594
rect 9524 2520 9994 2560
rect 5770 1798 5786 1832
rect 5870 1798 5886 1832
rect 6320 1664 6336 1698
rect 6420 1664 6436 1698
rect 6578 1664 6594 1698
rect 6678 1664 6694 1698
rect 6836 1664 6852 1698
rect 6936 1664 6952 1698
rect 6992 1624 7078 2000
rect 7586 1998 7668 2036
rect 7586 1950 8052 1998
rect 7996 1846 8052 1950
rect 7320 1664 7336 1698
rect 7420 1664 7436 1698
rect 7578 1664 7594 1698
rect 7678 1664 7694 1698
rect 7836 1664 7852 1698
rect 7936 1664 7952 1698
rect 6480 1554 7078 1624
rect 8006 1620 8050 1846
rect 8368 1748 8384 1782
rect 8468 1748 8484 1782
rect 7478 1618 7556 1620
rect 7680 1618 8052 1620
rect 6222 1420 6278 1446
rect 5682 1054 5716 1070
rect 5682 -350 5716 -334
rect 5940 1054 5974 1070
rect 5940 -350 5974 -334
rect 6222 1032 6232 1420
rect 6266 1032 6278 1420
rect 6222 464 6278 1032
rect 6480 1420 6536 1554
rect 6480 1032 6490 1420
rect 6524 1032 6536 1420
rect 6748 1420 6782 1436
rect 6320 708 6336 742
rect 6420 708 6436 742
rect 6222 76 6232 464
rect 6266 76 6278 464
rect 6222 -492 6278 76
rect 6480 464 6536 1032
rect 6740 1032 6748 1418
rect 6996 1420 7052 1554
rect 7478 1550 8052 1618
rect 7232 1426 7266 1436
rect 7484 1430 7534 1550
rect 7998 1544 8050 1550
rect 7748 1434 7782 1436
rect 6782 1032 6796 1418
rect 6996 1364 7006 1420
rect 6578 708 6594 742
rect 6678 708 6694 742
rect 6480 76 6490 464
rect 6524 76 6536 464
rect 6320 -248 6336 -214
rect 6420 -248 6436 -214
rect 6222 -854 6232 -492
rect 6218 -880 6232 -854
rect 6266 -880 6278 -492
rect 6218 -886 6278 -880
rect 6480 -492 6536 76
rect 6740 464 6796 1032
rect 6998 1032 7006 1364
rect 7040 1414 7052 1420
rect 7220 1420 7276 1426
rect 7040 1032 7054 1414
rect 6836 708 6852 742
rect 6936 708 6952 742
rect 6740 76 6748 464
rect 6782 76 6796 464
rect 6578 -248 6594 -214
rect 6678 -248 6694 -214
rect 6480 -880 6490 -492
rect 6524 -880 6536 -492
rect 6218 -982 6276 -886
rect 6480 -918 6536 -880
rect 6740 -492 6796 76
rect 6998 464 7054 1032
rect 6998 76 7006 464
rect 7040 76 7054 464
rect 6836 -248 6852 -214
rect 6936 -248 6952 -214
rect 6740 -880 6748 -492
rect 6782 -848 6796 -492
rect 6998 -492 7054 76
rect 6782 -880 6798 -848
rect 6740 -982 6798 -880
rect 6998 -880 7006 -492
rect 7040 -880 7054 -492
rect 6998 -918 7054 -880
rect 7220 1032 7232 1420
rect 7266 1032 7276 1420
rect 7220 464 7276 1032
rect 7482 1420 7538 1430
rect 7482 1032 7490 1420
rect 7524 1032 7538 1420
rect 7320 708 7336 742
rect 7420 708 7436 742
rect 7220 76 7232 464
rect 7266 76 7276 464
rect 7220 -492 7276 76
rect 7482 464 7538 1032
rect 7734 1420 7790 1434
rect 7998 1430 8048 1544
rect 7734 1032 7748 1420
rect 7782 1032 7790 1420
rect 7578 708 7594 742
rect 7678 708 7694 742
rect 7482 76 7490 464
rect 7524 76 7538 464
rect 7320 -248 7336 -214
rect 7420 -248 7436 -214
rect 7220 -880 7232 -492
rect 7266 -858 7276 -492
rect 7482 -492 7538 76
rect 7734 464 7790 1032
rect 7992 1420 8048 1430
rect 7992 1032 8006 1420
rect 8040 1032 8048 1420
rect 7836 708 7852 742
rect 7936 708 7952 742
rect 7734 76 7748 464
rect 7782 76 7790 464
rect 7578 -248 7594 -214
rect 7678 -248 7694 -214
rect 7266 -880 7280 -858
rect 7220 -906 7280 -880
rect 7482 -880 7490 -492
rect 7524 -880 7538 -492
rect 7482 -902 7538 -880
rect 7734 -492 7790 76
rect 7992 464 8048 1032
rect 7992 76 8006 464
rect 8040 76 8048 464
rect 7836 -248 7852 -214
rect 7936 -248 7952 -214
rect 7734 -880 7748 -492
rect 7782 -858 7790 -492
rect 7992 -492 8048 76
rect 8280 1004 8314 1020
rect 8280 -400 8314 -384
rect 8538 1004 8572 1020
rect 9734 478 11046 672
rect 9734 -16 9942 478
rect 10902 -16 11046 478
rect 9734 -236 11046 -16
rect 8538 -400 8572 -384
rect 7782 -880 7796 -858
rect 7734 -898 7796 -880
rect 7222 -982 7280 -906
rect 7738 -982 7796 -898
rect 7992 -880 8006 -492
rect 8040 -880 8048 -492
rect 7992 -902 8048 -880
rect 6214 -1090 7796 -982
rect 7092 -1308 7132 -1090
rect 5164 -1352 7132 -1308
rect 5164 -1354 7130 -1352
<< viali >>
rect 10364 10220 11324 10714
rect -7494 9394 -7097 9432
rect -3213 9394 -2816 9432
rect -2264 9394 -1867 9432
rect 2017 9394 2414 9432
rect 2966 9394 3363 9432
rect 7247 9394 7644 9432
rect 8196 9394 8593 9432
rect 12477 9394 12874 9432
rect -7494 9074 -7097 9112
rect -3213 9074 -2816 9112
rect -2264 9074 -1867 9112
rect 2017 9074 2414 9112
rect 2966 9074 3363 9112
rect 7247 9074 7644 9112
rect 8196 9074 8593 9112
rect 12477 9074 12874 9112
rect -7494 8754 -7097 8792
rect -3213 8754 -2816 8792
rect -2250 8732 -1853 8770
rect 2031 8732 2428 8770
rect 2946 8734 3343 8772
rect 7227 8734 7624 8772
rect 8196 8754 8593 8792
rect 12477 8754 12874 8792
rect -7494 8434 -7097 8472
rect -3213 8434 -2816 8472
rect -2250 8414 -1853 8452
rect 2031 8414 2428 8452
rect 2946 8416 3343 8454
rect 7227 8416 7624 8454
rect 8196 8434 8593 8472
rect 12477 8434 12874 8472
rect -7494 8114 -7097 8152
rect -3213 8114 -2816 8152
rect -2250 8096 -1853 8134
rect 2031 8096 2428 8134
rect 2946 8098 3343 8136
rect 7227 8098 7624 8136
rect 8196 8114 8593 8152
rect 12477 8114 12874 8152
rect -7494 7794 -7097 7832
rect -3213 7794 -2816 7832
rect -2250 7778 -1853 7816
rect 2031 7778 2428 7816
rect 2946 7780 3343 7818
rect 7227 7780 7624 7818
rect 8196 7794 8593 7832
rect 12477 7794 12874 7832
rect -7494 7474 -7097 7512
rect -3213 7474 -2816 7512
rect -2250 7460 -1853 7498
rect 2031 7460 2428 7498
rect 2946 7462 3343 7500
rect 7227 7462 7624 7500
rect 8196 7474 8593 7512
rect 12477 7474 12874 7512
rect -7494 7154 -7097 7192
rect -3213 7154 -2816 7192
rect -2250 7142 -1853 7180
rect 2031 7142 2428 7180
rect 2946 7144 3343 7182
rect 7227 7144 7624 7182
rect 8196 7154 8593 7192
rect 12477 7154 12874 7192
rect -7494 6834 -7097 6872
rect -3213 6834 -2816 6872
rect -2250 6824 -1853 6862
rect 2031 6824 2428 6862
rect 2946 6826 3343 6864
rect 7227 6826 7624 6864
rect 8196 6834 8593 6872
rect 12477 6834 12874 6872
rect -7494 6514 -7097 6552
rect -3213 6514 -2816 6552
rect -2250 6506 -1853 6544
rect 2031 6506 2428 6544
rect 2946 6508 3343 6546
rect 7227 6508 7624 6546
rect 8196 6514 8593 6552
rect 12477 6514 12874 6552
rect -7494 6194 -7097 6232
rect -3213 6194 -2816 6232
rect -2250 6188 -1853 6226
rect 2031 6188 2428 6226
rect 2946 6190 3343 6228
rect 7227 6190 7624 6228
rect 8196 6194 8593 6232
rect 12477 6194 12874 6232
rect -7494 5874 -7097 5912
rect -3213 5874 -2816 5912
rect -2230 5842 -1833 5880
rect 2051 5842 2448 5880
rect 2966 5872 3363 5910
rect 7247 5872 7644 5910
rect 8196 5874 8593 5912
rect 12477 5874 12874 5912
rect -7494 5554 -7097 5592
rect -3213 5554 -2816 5592
rect -2230 5522 -1833 5560
rect 2051 5522 2448 5560
rect 2966 5554 3363 5592
rect 7247 5554 7644 5592
rect 8196 5554 8593 5592
rect 12477 5554 12874 5592
rect -312 5002 -172 5126
rect -6262 4422 -5936 4662
rect -4912 4609 -4828 4643
rect -3710 4554 -3586 4646
rect -2350 4621 -2266 4655
rect -5016 3818 -4982 4306
rect -4758 3818 -4724 4306
rect -6562 3578 -6528 3672
rect -6562 3390 -6528 3578
rect -6562 3296 -6528 3390
rect -6474 3578 -6440 3672
rect -6474 3390 -6440 3578
rect -6474 3296 -6440 3390
rect -6330 3576 -6296 3670
rect -6330 3388 -6296 3576
rect -6330 3294 -6296 3388
rect -6242 3576 -6208 3670
rect -6242 3388 -6208 3576
rect -6242 3294 -6208 3388
rect -6102 3574 -6068 3668
rect -6102 3386 -6068 3574
rect -6102 3292 -6068 3386
rect -6014 3574 -5980 3668
rect -6014 3386 -5980 3574
rect -6014 3292 -5980 3386
rect -5884 3576 -5850 3670
rect -5884 3388 -5850 3576
rect -5884 3294 -5850 3388
rect -5796 3576 -5762 3670
rect -5796 3388 -5762 3576
rect -5796 3294 -5762 3388
rect -6538 2990 -6504 3034
rect -6538 2902 -6504 2990
rect -6538 2858 -6504 2902
rect -6450 2990 -6416 3034
rect -6450 2902 -6416 2990
rect -6450 2858 -6416 2902
rect -6322 2992 -6288 3036
rect -6322 2904 -6288 2992
rect -6322 2860 -6288 2904
rect -6234 2992 -6200 3036
rect -6234 2904 -6200 2992
rect -6234 2860 -6200 2904
rect -6104 2992 -6070 3036
rect -6104 2904 -6070 2992
rect -6104 2860 -6070 2904
rect -6016 2992 -5982 3036
rect -6016 2904 -5982 2992
rect -6016 2860 -5982 2904
rect -5882 2990 -5848 3034
rect -5882 2902 -5848 2990
rect -5882 2858 -5848 2902
rect -5794 2990 -5760 3034
rect -5794 2902 -5760 2990
rect -2454 3830 -2420 4318
rect -2196 3830 -2162 4318
rect -5794 2858 -5760 2902
rect -6210 2776 -6170 2814
rect -5932 2776 -5898 2810
rect -3968 2716 -3774 2892
rect -2954 2436 -2760 2612
rect -6 4952 46 5052
rect 174 4964 226 5048
rect 898 4972 976 5070
rect 2676 4966 2764 5098
rect -1374 4500 -1048 4740
rect -1376 3596 -1342 3690
rect -1376 3408 -1342 3596
rect -1376 3314 -1342 3408
rect -1288 3596 -1254 3690
rect -1288 3408 -1254 3596
rect -1288 3314 -1254 3408
rect -1144 3594 -1110 3688
rect -1144 3406 -1110 3594
rect -1144 3312 -1110 3406
rect -1056 3594 -1022 3688
rect -1056 3406 -1022 3594
rect -1056 3312 -1022 3406
rect -916 3592 -882 3686
rect -916 3404 -882 3592
rect -916 3310 -882 3404
rect -828 3592 -794 3686
rect -828 3404 -794 3592
rect -828 3310 -794 3404
rect -698 3594 -664 3688
rect -698 3406 -664 3594
rect -698 3312 -664 3406
rect -610 3594 -576 3688
rect -610 3406 -576 3594
rect -610 3312 -576 3406
rect -1352 3008 -1318 3052
rect -1352 2920 -1318 3008
rect -1352 2876 -1318 2920
rect -1264 3008 -1230 3052
rect -1264 2920 -1230 3008
rect -1264 2876 -1230 2920
rect -1136 3010 -1102 3054
rect -1136 2922 -1102 3010
rect -1136 2878 -1102 2922
rect -1048 3010 -1014 3054
rect -1048 2922 -1014 3010
rect -1048 2878 -1014 2922
rect -918 3010 -884 3054
rect -918 2922 -884 3010
rect -918 2878 -884 2922
rect -830 3010 -796 3054
rect -830 2922 -796 3010
rect -830 2878 -796 2922
rect -696 3008 -662 3052
rect -696 2920 -662 3008
rect -696 2876 -662 2920
rect -608 3008 -574 3052
rect -608 2920 -574 3008
rect -608 2876 -574 2920
rect -1024 2794 -984 2832
rect -746 2794 -712 2828
rect -1782 2604 -1720 2672
rect -4906 1216 -4822 1250
rect -4280 1218 -3896 1252
rect -5010 1034 -4976 1122
rect -4752 1034 -4718 1122
rect -4534 1036 -4500 1124
rect -3308 1218 -2924 1252
rect -3562 1036 -3528 1124
rect -2372 1216 -2288 1250
rect -2476 1034 -2442 1122
rect -2218 1034 -2184 1122
rect -4112 -150 -3152 344
rect 1610 4574 1742 4658
rect 2266 4634 2422 4744
rect 5142 4752 5224 4838
rect 6582 4766 6642 4820
rect 1024 4349 1108 4383
rect 920 3558 954 4046
rect 1178 3558 1212 4046
rect 1386 4038 1444 4054
rect 1386 3550 1399 4038
rect 1399 3550 1433 4038
rect 1433 3550 1444 4038
rect 1386 3540 1444 3550
rect 1915 3550 1949 4032
rect 1915 3544 1949 3550
rect 2055 4040 2095 4070
rect 2055 3552 2057 4040
rect 2057 3552 2091 4040
rect 2091 3552 2095 4040
rect 2055 3546 2095 3552
rect 1612 3116 1746 3204
rect 2573 3552 2607 4034
rect 2573 3546 2607 3552
rect 2818 4323 2902 4357
rect 3938 4288 4264 4528
rect 2714 3532 2748 4020
rect 2972 3532 3006 4020
rect 3328 3862 3438 3938
rect 3800 3608 3834 3702
rect 2564 2944 2608 3012
rect 3562 3152 3638 3222
rect 2878 2788 3080 2910
rect 2878 2490 3084 2622
rect 869 2310 969 2411
rect 3102 2362 3226 2414
rect 1392 2205 1452 2220
rect 1392 2055 1408 2205
rect 1408 2055 1442 2205
rect 1442 2055 1452 2205
rect 1392 2028 1452 2055
rect 1396 1649 1456 1674
rect 1396 1499 1408 1649
rect 1408 1499 1442 1649
rect 1442 1499 1456 1649
rect 1918 2205 1978 2236
rect 1918 2055 1924 2205
rect 1924 2055 1958 2205
rect 1958 2055 1978 2205
rect 1918 2044 1978 2055
rect 1396 1482 1456 1499
rect 1920 1649 1976 1680
rect 1920 1499 1924 1649
rect 1924 1499 1958 1649
rect 1958 1499 1976 1649
rect 1920 1488 1976 1499
rect 902 1174 944 1214
rect 2406 2205 2466 2220
rect 2406 2055 2422 2205
rect 2422 2055 2456 2205
rect 2456 2055 2466 2205
rect 2406 2028 2466 2055
rect 2410 1649 2470 1674
rect 2410 1499 2422 1649
rect 2422 1499 2456 1649
rect 2456 1499 2470 1649
rect 2932 2205 2992 2236
rect 2932 2055 2938 2205
rect 2938 2055 2972 2205
rect 2972 2055 2992 2205
rect 2932 2044 2992 2055
rect 2410 1482 2470 1499
rect 2934 1649 2990 1680
rect 2934 1499 2938 1649
rect 2938 1499 2972 1649
rect 2972 1499 2990 1649
rect 2934 1488 2990 1499
rect 1980 1110 2100 1246
rect 3316 1098 3436 1190
rect 3800 3420 3834 3608
rect 3800 3326 3834 3420
rect 3888 3608 3922 3702
rect 3888 3420 3922 3608
rect 3888 3326 3922 3420
rect 4032 3606 4066 3700
rect 4032 3418 4066 3606
rect 4032 3324 4066 3418
rect 4120 3606 4154 3700
rect 4120 3418 4154 3606
rect 4120 3324 4154 3418
rect 4260 3604 4294 3698
rect 4260 3416 4294 3604
rect 4260 3322 4294 3416
rect 4348 3604 4382 3698
rect 4348 3416 4382 3604
rect 4348 3322 4382 3416
rect 4478 3606 4512 3700
rect 4478 3418 4512 3606
rect 4478 3324 4512 3418
rect 4566 3606 4600 3700
rect 4566 3418 4600 3606
rect 4566 3324 4600 3418
rect 3824 3020 3858 3064
rect 3824 2932 3858 3020
rect 3824 2888 3858 2932
rect 3912 3020 3946 3064
rect 3912 2932 3946 3020
rect 3912 2888 3946 2932
rect 4040 3022 4074 3066
rect 4040 2934 4074 3022
rect 4040 2890 4074 2934
rect 4128 3022 4162 3066
rect 4128 2934 4162 3022
rect 4128 2890 4162 2934
rect 4258 3022 4292 3066
rect 4258 2934 4292 3022
rect 4258 2890 4292 2934
rect 4346 3022 4380 3066
rect 4346 2934 4380 3022
rect 4346 2890 4380 2934
rect 4480 3020 4514 3064
rect 4480 2932 4514 3020
rect 4480 2888 4514 2932
rect 4568 3020 4602 3064
rect 4568 2932 4602 3020
rect 4568 2888 4602 2932
rect 4152 2806 4192 2844
rect 4430 2806 4464 2840
rect 5050 1918 5110 2022
rect 4672 742 4816 874
rect 1612 602 1810 606
rect 1612 568 1625 602
rect 1625 568 1809 602
rect 1809 568 1810 602
rect 1612 566 1810 568
rect 2223 602 2427 604
rect 2223 568 2404 602
rect 2404 568 2427 602
rect 2223 566 2427 568
rect 3310 -334 4270 160
rect 6298 4221 6382 4255
rect 6742 4237 6926 4240
rect 6742 4203 6926 4237
rect 6742 4202 6926 4203
rect 6194 3430 6228 3918
rect 6452 3430 6486 3918
rect 8618 4706 8812 4770
rect 7146 4430 7206 4532
rect 7314 4237 7498 4242
rect 7314 4204 7498 4237
rect 8708 4600 8842 4650
rect 7886 4233 7970 4267
rect 9374 4230 9700 4470
rect 7782 3442 7816 3930
rect 8040 3442 8074 3930
rect 9456 3400 9490 3494
rect 9456 3212 9490 3400
rect 9456 3118 9490 3212
rect 9544 3400 9578 3494
rect 9544 3212 9578 3400
rect 9544 3118 9578 3212
rect 9688 3398 9722 3492
rect 9688 3210 9722 3398
rect 9688 3116 9722 3210
rect 9776 3398 9810 3492
rect 9776 3210 9810 3398
rect 9776 3116 9810 3210
rect 9916 3396 9950 3490
rect 9916 3208 9950 3396
rect 9916 3114 9950 3208
rect 10004 3396 10038 3490
rect 10004 3208 10038 3396
rect 10004 3114 10038 3208
rect 10134 3398 10168 3492
rect 10134 3210 10168 3398
rect 10134 3116 10168 3210
rect 10222 3398 10256 3492
rect 10222 3210 10256 3398
rect 10222 3116 10256 3210
rect 9480 2812 9514 2856
rect 9480 2724 9514 2812
rect 9480 2680 9514 2724
rect 9568 2812 9602 2856
rect 9568 2724 9602 2812
rect 9568 2680 9602 2724
rect 9696 2814 9730 2858
rect 9696 2726 9730 2814
rect 9696 2682 9730 2726
rect 9784 2814 9818 2858
rect 9784 2726 9818 2814
rect 9784 2682 9818 2726
rect 9914 2814 9948 2858
rect 9914 2726 9948 2814
rect 9914 2682 9948 2726
rect 10002 2814 10036 2858
rect 10002 2726 10036 2814
rect 10002 2682 10036 2726
rect 10136 2812 10170 2856
rect 10136 2724 10170 2812
rect 10136 2680 10170 2724
rect 10224 2812 10258 2856
rect 10224 2724 10258 2812
rect 10224 2680 10258 2724
rect 9808 2598 9848 2636
rect 10086 2598 10120 2632
rect 5786 1798 5870 1832
rect 6336 1664 6420 1698
rect 6594 1664 6678 1698
rect 6852 1664 6936 1698
rect 7336 1664 7420 1698
rect 7594 1664 7678 1698
rect 7852 1664 7936 1698
rect 8384 1748 8468 1782
rect 5682 -334 5716 1054
rect 5940 -334 5974 1054
rect 6336 708 6420 742
rect 6594 708 6678 742
rect 6336 -248 6420 -214
rect 6852 708 6936 742
rect 6594 -248 6678 -214
rect 6852 -248 6936 -214
rect 7336 708 7420 742
rect 7594 708 7678 742
rect 7336 -248 7420 -214
rect 7852 708 7936 742
rect 7594 -248 7678 -214
rect 7852 -248 7936 -214
rect 8280 -384 8314 1004
rect 8538 -384 8572 1004
rect 9942 -16 10902 478
<< metal1 >>
rect 10156 10714 11468 10908
rect 10156 10220 10364 10714
rect 11324 10220 11468 10714
rect 10156 10000 11468 10220
rect -7636 9530 8190 9562
rect 10482 9530 10542 10000
rect -7636 9432 12994 9530
rect -7636 9394 -7494 9432
rect -7097 9394 -3213 9432
rect -2816 9394 -2264 9432
rect -1867 9394 2017 9432
rect 2414 9394 2966 9432
rect 3363 9394 7247 9432
rect 7644 9394 8196 9432
rect 8593 9394 12477 9432
rect 12874 9394 12994 9432
rect -7636 9112 12994 9394
rect -7636 9074 -7494 9112
rect -7097 9074 -3213 9112
rect -2816 9074 -2264 9112
rect -1867 9074 2017 9112
rect 2414 9074 2966 9112
rect 3363 9074 7247 9112
rect 7644 9074 8196 9112
rect 8593 9074 12477 9112
rect 12874 9074 12994 9112
rect -7636 8946 12994 9074
rect -7636 8792 -2632 8946
rect -7636 8754 -7494 8792
rect -7097 8754 -3213 8792
rect -2816 8754 -2632 8792
rect -7636 8472 -2632 8754
rect -7636 8434 -7494 8472
rect -7097 8434 -3213 8472
rect -2816 8434 -2632 8472
rect -7636 8152 -2632 8434
rect -2282 8786 -1832 8800
rect -2282 8716 -2268 8786
rect -1836 8716 -1832 8786
rect -2282 8468 -1832 8716
rect 2008 8786 2462 8804
rect 2008 8716 2014 8786
rect 2446 8716 2462 8786
rect 2008 8698 2462 8716
rect 2916 8790 3366 8800
rect 2916 8716 2928 8790
rect 3362 8716 3366 8790
rect -2282 8398 -2268 8468
rect -1836 8398 -1832 8468
rect -2282 8388 -1832 8398
rect 2006 8468 2462 8482
rect 2006 8398 2014 8468
rect 2446 8398 2462 8468
rect -7636 8114 -7494 8152
rect -7097 8114 -3213 8152
rect -2816 8114 -2632 8152
rect -7636 7832 -2632 8114
rect -2280 8150 -1826 8170
rect -2280 8080 -2268 8150
rect -1836 8080 -1826 8150
rect -2280 8064 -1826 8080
rect 2006 8150 2462 8398
rect 2916 8470 3366 8716
rect 2916 8396 2928 8470
rect 3362 8396 3366 8470
rect 2916 8384 3366 8396
rect 7198 8788 7656 8800
rect 7198 8718 7210 8788
rect 7638 8718 7656 8788
rect 7198 8468 7656 8718
rect 7198 8398 7212 8468
rect 7640 8398 7656 8468
rect 2006 8080 2014 8150
rect 2446 8080 2462 8150
rect 2006 8066 2462 8080
rect 2916 8156 3370 8166
rect 2916 8082 2926 8156
rect 3360 8082 3370 8156
rect 2916 8072 3370 8082
rect 7198 8152 7656 8398
rect 7198 8082 7212 8152
rect 7640 8082 7656 8152
rect 7198 8062 7656 8082
rect 7990 8792 12994 8946
rect 7990 8754 8196 8792
rect 8593 8754 12477 8792
rect 12874 8754 12994 8792
rect 7990 8472 12994 8754
rect 7990 8434 8196 8472
rect 8593 8434 12477 8472
rect 12874 8434 12994 8472
rect 7990 8152 12994 8434
rect 7990 8114 8196 8152
rect 8593 8114 12477 8152
rect 12874 8114 12994 8152
rect -7636 7794 -7494 7832
rect -7097 7794 -3213 7832
rect -2816 7794 -2632 7832
rect -7636 7512 -2632 7794
rect -7636 7474 -7494 7512
rect -7097 7474 -3213 7512
rect -2816 7474 -2632 7512
rect -7636 7192 -2632 7474
rect -2274 7832 -1830 7840
rect -2274 7758 -2268 7832
rect -1834 7758 -1830 7832
rect -2274 7516 -1830 7758
rect -2274 7442 -2270 7516
rect -1836 7442 -1830 7516
rect -2274 7432 -1830 7442
rect 2000 7834 2456 7852
rect 2000 7762 2014 7834
rect 2446 7762 2456 7834
rect 2000 7516 2456 7762
rect 2000 7444 2014 7516
rect 2446 7444 2456 7516
rect -7636 7154 -7494 7192
rect -7097 7154 -3213 7192
rect -2816 7154 -2632 7192
rect -7636 6872 -2632 7154
rect -2276 7196 -1828 7206
rect -2276 7126 -2268 7196
rect -1836 7126 -1828 7196
rect -2276 7114 -1828 7126
rect 2000 7198 2456 7444
rect 2918 7834 3364 7846
rect 2918 7764 2928 7834
rect 3360 7764 3364 7834
rect 2918 7516 3364 7764
rect 7206 7834 7654 7844
rect 7206 7764 7210 7834
rect 7642 7764 7654 7834
rect 7206 7754 7654 7764
rect 7990 7832 12994 8114
rect 7990 7794 8196 7832
rect 8593 7794 12477 7832
rect 12874 7794 12994 7832
rect 2918 7446 2928 7516
rect 3360 7446 3364 7516
rect 2918 7434 3364 7446
rect 7206 7516 7652 7528
rect 7206 7446 7210 7516
rect 7642 7446 7652 7516
rect 2000 7124 2014 7198
rect 2446 7124 2456 7198
rect 2000 7112 2456 7124
rect 2918 7198 3366 7208
rect 2918 7128 2928 7198
rect 3360 7128 3366 7198
rect 2918 7118 3366 7128
rect 7206 7198 7652 7446
rect 7206 7128 7210 7198
rect 7642 7128 7652 7198
rect 7206 7116 7652 7128
rect 7990 7512 12994 7794
rect 7990 7474 8196 7512
rect 8593 7474 12477 7512
rect 12874 7474 12994 7512
rect 7990 7192 12994 7474
rect 7990 7154 8196 7192
rect 8593 7154 12477 7192
rect 12874 7154 12994 7192
rect -7636 6834 -7494 6872
rect -7097 6834 -3213 6872
rect -2816 6834 -2632 6872
rect -7636 6552 -2632 6834
rect -7636 6514 -7494 6552
rect -7097 6514 -3213 6552
rect -2816 6514 -2632 6552
rect -7636 6232 -2632 6514
rect -2282 6882 -1832 6890
rect -2282 6880 -1830 6882
rect -2282 6808 -2268 6880
rect -1842 6808 -1830 6880
rect -2282 6562 -1830 6808
rect -2282 6490 -2268 6562
rect -1842 6490 -1830 6562
rect -2282 6488 -1830 6490
rect 2010 6878 2456 6896
rect 2010 6806 2014 6878
rect 2446 6806 2456 6878
rect 2010 6562 2456 6806
rect 2920 6882 3374 6892
rect 2920 6808 2926 6882
rect 3364 6808 3374 6882
rect 2920 6798 3374 6808
rect 7200 6880 7654 6892
rect 7200 6810 7210 6880
rect 7642 6810 7654 6880
rect 7200 6798 7654 6810
rect 7990 6872 12994 7154
rect 7990 6834 8196 6872
rect 8593 6834 12477 6872
rect 12874 6834 12994 6872
rect 2010 6490 2014 6562
rect 2446 6490 2456 6562
rect -2282 6478 -1832 6488
rect 2010 6478 2456 6490
rect 2916 6564 3370 6580
rect 2916 6494 2926 6564
rect 3362 6494 3370 6564
rect -7636 6194 -7494 6232
rect -7097 6194 -3213 6232
rect -2816 6194 -2632 6232
rect -7636 6056 -2632 6194
rect -2276 6244 -1828 6256
rect -2276 6172 -2268 6244
rect -1836 6172 -1828 6244
rect -2276 6162 -1828 6172
rect 2010 6244 2458 6254
rect 2010 6172 2016 6244
rect 2444 6172 2458 6244
rect 2010 6160 2458 6172
rect 2916 6244 3370 6494
rect 2916 6174 2926 6244
rect 3362 6174 3370 6244
rect 2916 6154 3370 6174
rect 7202 6562 7658 6576
rect 7202 6492 7210 6562
rect 7646 6492 7658 6562
rect 7202 6244 7658 6492
rect 7202 6174 7210 6244
rect 7646 6174 7658 6244
rect 7202 6158 7658 6174
rect 7990 6552 12994 6834
rect 7990 6514 8196 6552
rect 8593 6514 12477 6552
rect 12874 6514 12994 6552
rect 7990 6232 12994 6514
rect 7990 6194 8196 6232
rect 8593 6194 12477 6232
rect 12874 6194 12994 6232
rect 7990 6056 12994 6194
rect -7636 5912 12994 6056
rect -7636 5874 -7494 5912
rect -7097 5874 -3213 5912
rect -2816 5910 8196 5912
rect -2816 5880 2966 5910
rect -2816 5874 -2230 5880
rect -7636 5842 -2230 5874
rect -1833 5842 2051 5880
rect 2448 5872 2966 5880
rect 3363 5872 7247 5910
rect 7644 5874 8196 5910
rect 8593 5874 12477 5912
rect 12874 5874 12994 5912
rect 7644 5872 12994 5874
rect 2448 5842 12994 5872
rect -7636 5592 12994 5842
rect -7636 5554 -7494 5592
rect -7097 5554 -3213 5592
rect -2816 5560 2966 5592
rect -2816 5554 -2230 5560
rect -7636 5522 -2230 5554
rect -1833 5522 2051 5560
rect 2448 5554 2966 5560
rect 3363 5554 7247 5592
rect 7644 5554 8196 5592
rect 8593 5554 12477 5592
rect 12874 5554 12994 5592
rect 2448 5522 12994 5554
rect -7636 5454 12994 5522
rect -3058 5424 12994 5454
rect 7990 5422 12994 5424
rect -3726 5250 -3558 5280
rect -3726 5172 -3704 5250
rect -3584 5172 -3558 5250
rect -3726 5138 -3558 5172
rect -6356 4662 -5842 4758
rect -6356 4422 -6262 4662
rect -5936 4546 -5842 4662
rect -5036 4643 -4704 4692
rect -3666 4682 -3626 5138
rect -344 5126 -134 5158
rect -344 5002 -312 5126
rect -172 5002 -134 5126
rect 2662 5098 2780 5124
rect -344 4972 -134 5002
rect -18 5052 58 5072
rect -1468 4740 -954 4836
rect -5036 4609 -4912 4643
rect -4828 4609 -4704 4643
rect -5036 4546 -4704 4609
rect -5936 4504 -4704 4546
rect -3750 4646 -3536 4682
rect -3750 4554 -3710 4646
rect -3586 4554 -3536 4646
rect -3750 4510 -3536 4554
rect -2472 4655 -2140 4696
rect -2472 4621 -2350 4655
rect -2266 4621 -2140 4655
rect -5936 4422 -5842 4504
rect -6356 4324 -5842 4422
rect -5036 4306 -4704 4504
rect -6444 3886 -5856 3888
rect -6444 3852 -5380 3886
rect -6444 3848 -5856 3852
rect -6444 3686 -6390 3848
rect -5906 3846 -5856 3848
rect -6666 3672 -6522 3686
rect -6476 3684 -6390 3686
rect -6666 3526 -6562 3672
rect -6666 3462 -6648 3526
rect -6588 3462 -6562 3526
rect -6666 3296 -6562 3462
rect -6528 3296 -6522 3672
rect -6666 3284 -6522 3296
rect -6480 3672 -6390 3684
rect -6334 3784 -5966 3818
rect -6334 3682 -6302 3784
rect -6016 3782 -5966 3784
rect -6006 3686 -5966 3782
rect -6480 3296 -6474 3672
rect -6440 3296 -6390 3672
rect -6480 3286 -6390 3296
rect -6336 3670 -6290 3682
rect -6336 3294 -6330 3670
rect -6296 3294 -6290 3670
rect -6480 3284 -6426 3286
rect -6578 3178 -6534 3284
rect -6336 3282 -6290 3294
rect -6252 3670 -6180 3682
rect -6252 3508 -6242 3670
rect -6208 3508 -6180 3670
rect -6252 3444 -6250 3508
rect -6186 3444 -6180 3508
rect -6252 3294 -6242 3444
rect -6208 3294 -6180 3444
rect -6252 3282 -6180 3294
rect -6152 3668 -6062 3686
rect -6006 3680 -5944 3686
rect -5896 3682 -5856 3846
rect -5800 3682 -5724 3684
rect -5896 3680 -5844 3682
rect -6020 3678 -5944 3680
rect -6152 3620 -6102 3668
rect -6068 3620 -6062 3668
rect -6152 3550 -6144 3620
rect -6066 3550 -6062 3620
rect -6152 3292 -6102 3550
rect -6068 3292 -6062 3550
rect -6028 3668 -5944 3678
rect -6028 3516 -6014 3668
rect -6020 3448 -6014 3516
rect -6330 3182 -6302 3282
rect -6152 3280 -6062 3292
rect -6028 3410 -6014 3448
rect -5980 3410 -5944 3668
rect -6028 3344 -6020 3410
rect -5948 3344 -5944 3410
rect -6028 3292 -6014 3344
rect -5980 3292 -5944 3344
rect -6028 3282 -5944 3292
rect -5890 3670 -5844 3680
rect -5890 3294 -5884 3670
rect -5850 3294 -5844 3670
rect -5890 3282 -5844 3294
rect -5802 3670 -5724 3682
rect -5802 3624 -5796 3670
rect -5762 3624 -5724 3670
rect -5802 3558 -5800 3624
rect -5728 3558 -5724 3624
rect -5802 3294 -5796 3558
rect -5762 3294 -5724 3558
rect -5802 3282 -5724 3294
rect -6578 3150 -6390 3178
rect -6330 3154 -6174 3182
rect -6418 3046 -6390 3150
rect -6210 3050 -6174 3154
rect -6116 3180 -6078 3280
rect -6028 3278 -5952 3282
rect -6116 3152 -5958 3180
rect -6210 3048 -6126 3050
rect -5994 3048 -5958 3152
rect -5890 3178 -5856 3282
rect -5890 3150 -5730 3178
rect -6328 3046 -6282 3048
rect -6544 3036 -6498 3046
rect -6582 3034 -6498 3036
rect -6582 2970 -6538 3034
rect -6582 2912 -6568 2970
rect -6582 2858 -6538 2912
rect -6504 2858 -6498 3034
rect -6582 2848 -6498 2858
rect -6544 2846 -6498 2848
rect -6456 3036 -6282 3046
rect -6456 3034 -6322 3036
rect -6456 2858 -6450 3034
rect -6416 2860 -6322 3034
rect -6288 2860 -6282 3036
rect -6416 2858 -6282 2860
rect -6456 2848 -6282 2858
rect -6240 3046 -6064 3048
rect -6022 3046 -5888 3048
rect -5770 3046 -5730 3150
rect -6240 3036 -6062 3046
rect -6240 2860 -6234 3036
rect -6200 2860 -6104 3036
rect -6070 2860 -6062 3036
rect -6240 2852 -6062 2860
rect -6022 3036 -5842 3046
rect -6022 2860 -6016 3036
rect -5982 3034 -5842 3036
rect -5982 2860 -5882 3034
rect -6022 2858 -5882 2860
rect -5848 2858 -5842 3034
rect -6240 2850 -6064 2852
rect -6240 2848 -6194 2850
rect -6128 2848 -6064 2850
rect -6022 2850 -5842 2858
rect -6022 2848 -5976 2850
rect -6456 2846 -6296 2848
rect -6128 2846 -6088 2848
rect -5888 2846 -5842 2850
rect -5800 3034 -5722 3046
rect -5800 2858 -5794 3034
rect -5760 2968 -5722 3034
rect -5734 2910 -5722 2968
rect -5760 2858 -5722 2910
rect -5800 2852 -5722 2858
rect -5800 2846 -5754 2852
rect -6216 2818 -6164 2820
rect -5416 2818 -5380 3852
rect -5036 3818 -5016 4306
rect -4982 3818 -4758 4306
rect -4724 3818 -4704 4306
rect -5036 3694 -4704 3818
rect -2472 4318 -2140 4621
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect -1468 4402 -954 4500
rect -2472 3830 -2454 4318
rect -2420 3830 -2196 4318
rect -2162 3830 -2140 4318
rect -2472 3694 -2140 3830
rect -1258 3866 -670 3906
rect -1258 3704 -1204 3866
rect -720 3864 -670 3866
rect -5036 3646 -2140 3694
rect -5036 3520 -4704 3646
rect -2472 3524 -2140 3646
rect -1480 3690 -1336 3704
rect -1290 3702 -1204 3704
rect -1480 3544 -1376 3690
rect -1480 3480 -1462 3544
rect -1402 3480 -1376 3544
rect -1480 3314 -1376 3480
rect -1342 3314 -1336 3690
rect -1480 3302 -1336 3314
rect -1294 3690 -1204 3702
rect -1148 3802 -780 3836
rect -1148 3700 -1116 3802
rect -830 3800 -780 3802
rect -820 3704 -780 3800
rect -1294 3314 -1288 3690
rect -1254 3314 -1204 3690
rect -1294 3304 -1204 3314
rect -1150 3688 -1104 3700
rect -1150 3312 -1144 3688
rect -1110 3312 -1104 3688
rect -1294 3302 -1240 3304
rect -1392 3196 -1348 3302
rect -1150 3300 -1104 3312
rect -1066 3688 -994 3700
rect -1066 3526 -1056 3688
rect -1022 3526 -994 3688
rect -1066 3462 -1064 3526
rect -1000 3462 -994 3526
rect -1066 3312 -1056 3462
rect -1022 3312 -994 3462
rect -1066 3300 -994 3312
rect -966 3686 -876 3704
rect -820 3698 -758 3704
rect -710 3700 -670 3864
rect -614 3700 -538 3702
rect -710 3698 -658 3700
rect -834 3696 -758 3698
rect -966 3638 -916 3686
rect -882 3638 -876 3686
rect -966 3568 -958 3638
rect -880 3568 -876 3638
rect -966 3310 -916 3568
rect -882 3310 -876 3568
rect -842 3686 -758 3696
rect -842 3534 -828 3686
rect -834 3466 -828 3534
rect -1144 3200 -1116 3300
rect -966 3298 -876 3310
rect -842 3428 -828 3466
rect -794 3428 -758 3686
rect -842 3362 -834 3428
rect -762 3362 -758 3428
rect -842 3310 -828 3362
rect -794 3310 -758 3362
rect -842 3300 -758 3310
rect -704 3688 -658 3698
rect -704 3312 -698 3688
rect -664 3312 -658 3688
rect -704 3300 -658 3312
rect -616 3688 -538 3700
rect -616 3642 -610 3688
rect -576 3642 -538 3688
rect -616 3576 -614 3642
rect -542 3636 -538 3642
rect -276 3640 -236 4972
rect -18 4952 -6 5052
rect 46 4952 58 5052
rect -18 4932 58 4952
rect 158 5048 244 5072
rect 158 4964 174 5048
rect 226 4964 244 5048
rect 158 4940 244 4964
rect 886 5070 986 5090
rect 886 4972 898 5070
rect 976 4972 986 5070
rect 886 4940 986 4972
rect 2662 4966 2676 5098
rect 2764 4966 2780 5098
rect 2662 4946 2780 4966
rect 7140 4882 7238 4900
rect 5128 4838 5236 4850
rect 258 4764 490 4788
rect 258 4712 282 4764
rect 458 4752 490 4764
rect 2246 4752 2444 4776
rect 458 4744 2444 4752
rect 458 4712 2266 4744
rect 258 4692 490 4712
rect -196 4668 -56 4686
rect -196 4582 -180 4668
rect -72 4640 -56 4668
rect 1584 4658 1770 4684
rect 1584 4640 1610 4658
rect -72 4592 1610 4640
rect -72 4590 346 4592
rect -72 4582 -56 4590
rect -196 4562 -56 4582
rect 1584 4574 1610 4592
rect 1742 4574 1770 4658
rect 2246 4634 2266 4712
rect 2422 4634 2444 4744
rect 5128 4752 5142 4838
rect 5224 4752 5236 4838
rect 5128 4734 5236 4752
rect 6560 4820 6658 4826
rect 6560 4766 6582 4820
rect 6642 4766 6658 4820
rect 7140 4822 7158 4882
rect 7220 4822 7238 4882
rect 6560 4750 6658 4766
rect 6830 4760 6882 4812
rect 7140 4804 7238 4822
rect 2246 4598 2444 4634
rect 1584 4546 1770 4574
rect 2802 4510 2918 4550
rect 3844 4528 4358 4624
rect 1196 4504 2918 4510
rect 3068 4504 3174 4524
rect 1196 4464 3174 4504
rect 1196 4460 2918 4464
rect 1198 4392 1236 4460
rect 1016 4389 1236 4392
rect 1012 4383 1236 4389
rect 1012 4349 1024 4383
rect 1108 4349 1236 4383
rect 2802 4358 2918 4460
rect 3068 4454 3174 4464
rect 1012 4343 1236 4349
rect 1016 4342 1236 4343
rect 2794 4357 3272 4358
rect 2794 4323 2818 4357
rect 2902 4323 3272 4357
rect 2794 4310 3272 4323
rect 3844 4288 3938 4528
rect 4264 4288 4358 4528
rect 3844 4190 4358 4288
rect 6144 4255 6532 4288
rect 6144 4221 6298 4255
rect 6382 4221 6532 4255
rect 6832 4250 6880 4760
rect 7164 4578 7204 4804
rect 8586 4770 8844 4788
rect 8586 4706 8618 4770
rect 8812 4752 8844 4770
rect 8812 4714 10626 4752
rect 8812 4706 8844 4714
rect 8586 4688 8844 4706
rect 8696 4650 8866 4656
rect 8696 4600 8708 4650
rect 8842 4600 8866 4650
rect 8696 4592 8866 4600
rect 7124 4532 7238 4578
rect 7124 4430 7146 4532
rect 7206 4430 7238 4532
rect 7124 4378 7238 4430
rect 7734 4267 8122 4316
rect 4090 4134 4130 4190
rect 6144 4134 6532 4221
rect 6720 4242 7520 4250
rect 6720 4240 7314 4242
rect 6720 4202 6742 4240
rect 6926 4204 7314 4240
rect 7498 4204 7520 4242
rect 6926 4202 7520 4204
rect 6720 4190 7520 4202
rect 7734 4233 7886 4267
rect 7970 4233 8122 4267
rect 4090 4106 6532 4134
rect 4098 4098 6532 4106
rect 1366 4070 1449 4090
rect 2025 4072 2107 4092
rect 2025 4070 2651 4072
rect 1174 4058 1226 4064
rect 914 4046 960 4058
rect -276 3636 242 3640
rect -542 3596 242 3636
rect -542 3592 -236 3596
rect -542 3576 -538 3592
rect -616 3312 -610 3576
rect -576 3312 -538 3576
rect -616 3300 -538 3312
rect -1392 3168 -1204 3196
rect -1144 3172 -988 3200
rect -1232 3064 -1204 3168
rect -1024 3068 -988 3172
rect -930 3198 -892 3298
rect -842 3296 -766 3300
rect -930 3170 -772 3198
rect -1024 3066 -940 3068
rect -808 3066 -772 3170
rect -704 3196 -670 3300
rect 198 3206 238 3596
rect 914 3558 920 4046
rect 954 3558 960 4046
rect 914 3546 960 3558
rect 1172 4046 1226 4058
rect 1172 3558 1178 4046
rect 1212 3558 1226 4046
rect 1366 4054 1993 4070
rect 1366 3962 1386 4054
rect 1172 3546 1226 3558
rect 198 3200 534 3206
rect 1174 3200 1226 3546
rect 1367 3540 1386 3962
rect 1444 4032 1993 4054
rect 1444 3544 1915 4032
rect 1949 3544 1993 4032
rect 1444 3540 1993 3544
rect 1367 3512 1993 3540
rect 2025 3546 2055 4070
rect 2095 4034 2651 4070
rect 2095 3546 2573 4034
rect 2607 3546 2651 4034
rect 2025 3514 2651 3546
rect 2708 4020 2754 4032
rect 2708 3532 2714 4020
rect 2748 3532 2754 4020
rect 2708 3520 2754 3532
rect 2966 4020 3012 4032
rect 2966 3532 2972 4020
rect 3006 3532 3012 4020
rect 3298 3938 3474 3970
rect 3298 3862 3328 3938
rect 3438 3910 3474 3938
rect 6144 3918 6532 4098
rect 3918 3910 4506 3918
rect 3438 3878 4506 3910
rect 3438 3868 3972 3878
rect 4456 3876 4506 3878
rect 3438 3862 3474 3868
rect 3298 3820 3474 3862
rect 3918 3716 3972 3868
rect 2966 3520 3012 3532
rect 3696 3702 3840 3716
rect 3886 3714 3972 3716
rect 3696 3556 3800 3702
rect 3696 3492 3714 3556
rect 3774 3492 3800 3556
rect 3696 3326 3800 3492
rect 3834 3326 3840 3702
rect 3696 3314 3840 3326
rect 3882 3702 3972 3714
rect 4028 3814 4396 3848
rect 4028 3712 4060 3814
rect 4346 3812 4396 3814
rect 4356 3716 4396 3812
rect 3882 3326 3888 3702
rect 3922 3326 3972 3702
rect 3882 3316 3972 3326
rect 4026 3700 4072 3712
rect 4026 3324 4032 3700
rect 4066 3324 4072 3700
rect 3882 3314 3936 3316
rect -704 3168 -544 3196
rect -584 3134 -544 3168
rect 198 3166 1226 3200
rect 204 3162 1226 3166
rect 384 3160 1226 3162
rect 1580 3204 1782 3230
rect -188 3134 -136 3136
rect -584 3088 -136 3134
rect -1142 3064 -1096 3066
rect -1358 3054 -1312 3064
rect -1396 3052 -1312 3054
rect -1396 2988 -1352 3052
rect -4006 2892 -3742 2934
rect -4006 2818 -3968 2892
rect -6240 2814 -5886 2818
rect -6240 2776 -6210 2814
rect -6170 2810 -5886 2814
rect -6170 2776 -5932 2810
rect -5898 2776 -5886 2810
rect -6240 2772 -5886 2776
rect -5416 2772 -3968 2818
rect -6216 2770 -6164 2772
rect -5942 2766 -5886 2772
rect -4006 2716 -3968 2772
rect -3774 2716 -3742 2892
rect -1396 2930 -1382 2988
rect -1396 2876 -1352 2930
rect -1318 2876 -1312 3052
rect -1396 2866 -1312 2876
rect -1358 2864 -1312 2866
rect -1270 3054 -1096 3064
rect -1270 3052 -1136 3054
rect -1270 2876 -1264 3052
rect -1230 2878 -1136 3052
rect -1102 2878 -1096 3054
rect -1230 2876 -1096 2878
rect -1270 2866 -1096 2876
rect -1054 3064 -878 3066
rect -836 3064 -702 3066
rect -584 3064 -536 3088
rect -1054 3054 -876 3064
rect -1054 2878 -1048 3054
rect -1014 2878 -918 3054
rect -884 2878 -876 3054
rect -1054 2870 -876 2878
rect -836 3054 -656 3064
rect -836 2878 -830 3054
rect -796 3052 -656 3054
rect -796 2878 -696 3052
rect -836 2876 -696 2878
rect -662 2876 -656 3052
rect -1054 2868 -878 2870
rect -1054 2866 -1008 2868
rect -942 2866 -878 2868
rect -836 2868 -656 2876
rect -836 2866 -790 2868
rect -1270 2864 -1110 2866
rect -942 2864 -902 2866
rect -702 2864 -656 2868
rect -614 3052 -536 3064
rect -614 2876 -608 3052
rect -574 2986 -536 3052
rect -548 2928 -536 2986
rect -188 2970 -136 3088
rect 288 3108 446 3120
rect 288 3054 314 3108
rect 420 3096 446 3108
rect 1580 3116 1612 3204
rect 1746 3116 1782 3204
rect 3544 3222 3660 3236
rect 3544 3152 3562 3222
rect 3638 3210 3660 3222
rect 3784 3210 3828 3314
rect 4026 3312 4072 3324
rect 4110 3700 4182 3712
rect 4110 3538 4120 3700
rect 4154 3538 4182 3700
rect 4110 3474 4112 3538
rect 4176 3474 4182 3538
rect 4110 3324 4120 3474
rect 4154 3324 4182 3474
rect 4110 3312 4182 3324
rect 4210 3698 4300 3716
rect 4356 3710 4418 3716
rect 4466 3712 4506 3876
rect 4562 3712 4638 3714
rect 4466 3710 4518 3712
rect 4342 3708 4418 3710
rect 4210 3650 4260 3698
rect 4294 3650 4300 3698
rect 4210 3580 4218 3650
rect 4296 3580 4300 3650
rect 4210 3322 4260 3580
rect 4294 3322 4300 3580
rect 4334 3698 4418 3708
rect 4334 3546 4348 3698
rect 4342 3478 4348 3546
rect 3638 3208 3828 3210
rect 4032 3212 4060 3312
rect 4210 3310 4300 3322
rect 4334 3440 4348 3478
rect 4382 3440 4418 3698
rect 4334 3374 4342 3440
rect 4414 3374 4418 3440
rect 4334 3322 4348 3374
rect 4382 3322 4418 3374
rect 4334 3312 4418 3322
rect 4472 3700 4518 3710
rect 4472 3324 4478 3700
rect 4512 3324 4518 3700
rect 4472 3312 4518 3324
rect 4560 3700 4638 3712
rect 4560 3654 4566 3700
rect 4600 3698 4638 3700
rect 4600 3654 4994 3698
rect 4560 3588 4562 3654
rect 4634 3652 4994 3654
rect 4634 3588 4638 3652
rect 4560 3324 4566 3588
rect 4600 3324 4638 3588
rect 4560 3312 4638 3324
rect 3638 3180 3972 3208
rect 4032 3184 4188 3212
rect 3638 3176 3816 3180
rect 3638 3152 3660 3176
rect 3544 3134 3660 3152
rect 1580 3096 1782 3116
rect 420 3086 1782 3096
rect 420 3064 1698 3086
rect 3944 3076 3972 3180
rect 4152 3080 4188 3184
rect 4246 3210 4284 3310
rect 4334 3308 4410 3312
rect 4246 3182 4404 3210
rect 4152 3078 4236 3080
rect 4368 3078 4404 3182
rect 4472 3208 4506 3312
rect 4472 3180 4632 3208
rect 4034 3076 4080 3078
rect 3818 3066 3864 3076
rect 3780 3064 3864 3066
rect 420 3054 446 3064
rect 288 3040 446 3054
rect 2552 3012 2616 3028
rect 2552 2970 2564 3012
rect -190 2944 2564 2970
rect 2608 2944 2616 3012
rect -190 2934 2616 2944
rect 3780 3000 3824 3064
rect 3780 2942 3794 3000
rect -574 2876 -536 2928
rect 2552 2926 2616 2934
rect 2852 2910 3120 2942
rect 2852 2876 2878 2910
rect -614 2870 -536 2876
rect 348 2874 2878 2876
rect -614 2864 -568 2870
rect -4006 2684 -3742 2716
rect -1816 2672 -1676 2708
rect -3000 2612 -2736 2650
rect -5446 2526 -5326 2548
rect -5446 2458 -5426 2526
rect -5350 2512 -5326 2526
rect -3000 2512 -2954 2612
rect -5350 2466 -2954 2512
rect -5350 2458 -5326 2466
rect -5446 2432 -5326 2458
rect -3000 2436 -2954 2466
rect -2760 2436 -2736 2612
rect -1816 2604 -1782 2672
rect -1720 2660 -1676 2672
rect -1204 2660 -1164 2864
rect -1030 2836 -978 2838
rect -1054 2832 -700 2836
rect -1054 2794 -1024 2832
rect -984 2828 -700 2832
rect -984 2794 -746 2828
rect -712 2794 -700 2828
rect -1054 2790 -700 2794
rect -1030 2788 -978 2790
rect -756 2784 -700 2790
rect 334 2826 2878 2874
rect -1720 2640 -1160 2660
rect 334 2640 388 2826
rect 2852 2788 2878 2826
rect 3080 2788 3120 2910
rect 3780 2888 3824 2942
rect 3858 2888 3864 3064
rect 3780 2878 3864 2888
rect 3818 2876 3864 2878
rect 3906 3066 4080 3076
rect 3906 3064 4040 3066
rect 3906 2888 3912 3064
rect 3946 2890 4040 3064
rect 4074 2890 4080 3066
rect 3946 2888 4080 2890
rect 3906 2878 4080 2888
rect 4122 3076 4298 3078
rect 4340 3076 4474 3078
rect 4592 3076 4632 3180
rect 4122 3066 4300 3076
rect 4122 2890 4128 3066
rect 4162 2890 4258 3066
rect 4292 2890 4300 3066
rect 4122 2882 4300 2890
rect 4340 3066 4520 3076
rect 4340 2890 4346 3066
rect 4380 3064 4520 3066
rect 4380 2890 4480 3064
rect 4340 2888 4480 2890
rect 4514 2888 4520 3064
rect 4122 2880 4298 2882
rect 4122 2878 4168 2880
rect 4234 2878 4298 2880
rect 4340 2880 4520 2888
rect 4340 2878 4386 2880
rect 3906 2876 4066 2878
rect 4234 2876 4274 2878
rect 4474 2876 4520 2880
rect 4562 3064 4640 3076
rect 4562 2888 4568 3064
rect 4602 2998 4640 3064
rect 4628 2940 4640 2998
rect 4602 2888 4640 2940
rect 4562 2882 4640 2888
rect 4562 2876 4608 2882
rect 4146 2848 4198 2850
rect 4122 2844 4476 2848
rect 4122 2806 4152 2844
rect 4192 2840 4476 2844
rect 4192 2806 4430 2840
rect 4464 2806 4476 2840
rect 4122 2802 4476 2806
rect 4146 2800 4198 2802
rect 4420 2796 4476 2802
rect 2852 2752 3120 2788
rect -1720 2604 388 2640
rect -1816 2602 388 2604
rect 2854 2622 3112 2648
rect -1816 2580 -1676 2602
rect -1252 2598 374 2602
rect -1204 2596 -1164 2598
rect 2854 2490 2878 2622
rect 3084 2490 3112 2622
rect -3000 2400 -2736 2436
rect 851 2411 1998 2477
rect 2854 2476 3112 2490
rect 851 2310 869 2411
rect 969 2310 1998 2411
rect 851 2245 1998 2310
rect 2092 2466 3112 2476
rect 2092 2245 3012 2466
rect 3076 2414 3252 2432
rect 3076 2362 3102 2414
rect 3226 2362 3252 2414
rect 3076 2344 3252 2362
rect 1108 2236 1998 2245
rect 1108 2220 1918 2236
rect 1108 2028 1392 2220
rect 1452 2044 1918 2220
rect 1978 2044 1998 2236
rect 1452 2028 1998 2044
rect 1108 1680 1998 2028
rect 1108 1674 1920 1680
rect -2064 1566 -2008 1570
rect -3600 1522 -2008 1566
rect -5032 1250 -4700 1284
rect -3600 1274 -3554 1522
rect -2064 1520 -2008 1522
rect 1108 1482 1396 1674
rect 1456 1488 1920 1674
rect 1976 1488 1998 1680
rect 1456 1482 1998 1488
rect 1108 1390 1998 1482
rect 2122 2236 3012 2245
rect 2122 2220 2932 2236
rect 2122 2028 2406 2220
rect 2466 2044 2932 2220
rect 2992 2044 3012 2236
rect 2466 2028 3012 2044
rect 2122 1680 3012 2028
rect 2122 1674 2934 1680
rect 2122 1482 2410 1674
rect 2470 1488 2934 1674
rect 2990 1488 3012 1680
rect 2470 1482 3012 1488
rect 2122 1390 3012 1482
rect -5032 1216 -4906 1250
rect -4822 1216 -4700 1250
rect -5032 1122 -4700 1216
rect -4302 1252 -2896 1274
rect -4302 1218 -4280 1252
rect -3896 1218 -3308 1252
rect -2924 1218 -2896 1252
rect -4302 1202 -2896 1218
rect -2482 1250 -2150 1276
rect -2482 1216 -2372 1250
rect -2288 1216 -2150 1250
rect 1952 1246 2136 1274
rect -5032 1034 -5010 1122
rect -4976 1034 -4752 1122
rect -4718 1034 -4700 1122
rect -5032 944 -4700 1034
rect -4548 1136 -3514 1154
rect -4548 1124 -3502 1136
rect -4548 1036 -4534 1124
rect -4500 1036 -3562 1124
rect -3528 1036 -3502 1124
rect -4548 1014 -3502 1036
rect -4900 896 -4850 944
rect -3580 896 -3502 1014
rect -2482 1122 -2150 1216
rect 888 1214 1246 1226
rect 888 1174 902 1214
rect 944 1174 1246 1214
rect 888 1162 1246 1174
rect -2482 1034 -2476 1122
rect -2442 1034 -2218 1122
rect -2184 1034 -2150 1122
rect -2482 936 -2150 1034
rect -2368 896 -2318 936
rect -4906 860 -2318 896
rect -4906 844 -2324 860
rect -3646 538 -3604 844
rect 1200 628 1246 1162
rect 1952 1110 1980 1246
rect 2100 1224 2136 1246
rect 3078 1244 3224 1254
rect 3078 1224 3092 1244
rect 2100 1182 3092 1224
rect 3210 1182 3224 1244
rect 2100 1178 3224 1182
rect 2100 1110 2136 1178
rect 3078 1170 3224 1178
rect 3280 1190 3470 1220
rect 1952 1076 2136 1110
rect 3280 1098 3316 1190
rect 3436 1164 3470 1190
rect 4952 1164 4994 3652
rect 6144 3430 6194 3918
rect 6228 3430 6452 3918
rect 6486 3612 6532 3918
rect 7734 3930 8122 4233
rect 7734 3612 7782 3930
rect 6486 3576 7782 3612
rect 6486 3430 6532 3576
rect 6144 3108 6532 3430
rect 7734 3442 7782 3576
rect 7816 3442 8040 3930
rect 8074 3442 8122 3930
rect 7734 3136 8122 3442
rect 8826 3010 8862 4592
rect 9280 4470 9794 4566
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
rect 9002 3754 9140 3780
rect 9002 3654 9028 3754
rect 9110 3708 9140 3754
rect 9574 3708 10162 3710
rect 9110 3670 10162 3708
rect 9110 3654 9140 3670
rect 9002 3624 9140 3654
rect 9574 3508 9628 3670
rect 10112 3668 10162 3670
rect 9352 3494 9496 3508
rect 9542 3506 9628 3508
rect 9352 3348 9456 3494
rect 9352 3284 9370 3348
rect 9430 3284 9456 3348
rect 9352 3118 9456 3284
rect 9490 3118 9496 3494
rect 9352 3106 9496 3118
rect 9538 3494 9628 3506
rect 9684 3606 10052 3640
rect 9684 3504 9716 3606
rect 10002 3604 10052 3606
rect 10012 3508 10052 3604
rect 9538 3118 9544 3494
rect 9578 3118 9628 3494
rect 9538 3108 9628 3118
rect 9682 3492 9728 3504
rect 9682 3116 9688 3492
rect 9722 3116 9728 3492
rect 9538 3106 9592 3108
rect 9440 3010 9484 3106
rect 9682 3104 9728 3116
rect 9766 3492 9838 3504
rect 9766 3330 9776 3492
rect 9810 3330 9838 3492
rect 9766 3266 9768 3330
rect 9832 3266 9838 3330
rect 9766 3116 9776 3266
rect 9810 3116 9838 3266
rect 9766 3104 9838 3116
rect 9866 3490 9956 3508
rect 10012 3502 10074 3508
rect 10122 3504 10162 3668
rect 10218 3504 10294 3506
rect 10122 3502 10174 3504
rect 9998 3500 10074 3502
rect 9866 3442 9916 3490
rect 9950 3442 9956 3490
rect 9866 3372 9874 3442
rect 9952 3372 9956 3442
rect 9866 3114 9916 3372
rect 9950 3114 9956 3372
rect 9990 3490 10074 3500
rect 9990 3338 10004 3490
rect 9998 3270 10004 3338
rect 8826 3000 9484 3010
rect 9688 3004 9716 3104
rect 9866 3102 9956 3114
rect 9990 3232 10004 3270
rect 10038 3232 10074 3490
rect 9990 3166 9998 3232
rect 10070 3166 10074 3232
rect 9990 3114 10004 3166
rect 10038 3114 10074 3166
rect 9990 3104 10074 3114
rect 10128 3492 10174 3502
rect 10128 3116 10134 3492
rect 10168 3116 10174 3492
rect 10128 3104 10174 3116
rect 10216 3492 10294 3504
rect 10578 3492 10616 4714
rect 10216 3446 10222 3492
rect 10256 3454 10616 3492
rect 10256 3446 10294 3454
rect 10216 3380 10218 3446
rect 10290 3380 10294 3446
rect 10578 3442 10616 3454
rect 10216 3116 10222 3380
rect 10256 3116 10294 3380
rect 10216 3104 10294 3116
rect 8826 2974 9628 3000
rect 9688 2976 9844 3004
rect 9440 2972 9628 2974
rect 9600 2868 9628 2972
rect 9808 2872 9844 2976
rect 9902 3002 9940 3102
rect 9990 3100 10066 3104
rect 9902 2974 10060 3002
rect 9808 2870 9892 2872
rect 10024 2870 10060 2974
rect 10128 3000 10162 3104
rect 10128 2972 10288 3000
rect 9690 2868 9736 2870
rect 9474 2858 9520 2868
rect 9436 2856 9520 2858
rect 9436 2792 9480 2856
rect 9436 2734 9450 2792
rect 9436 2680 9480 2734
rect 9514 2680 9520 2856
rect 9436 2670 9520 2680
rect 9474 2668 9520 2670
rect 9562 2858 9736 2868
rect 9562 2856 9696 2858
rect 9562 2680 9568 2856
rect 9602 2682 9696 2856
rect 9730 2682 9736 2858
rect 9602 2680 9736 2682
rect 9562 2670 9736 2680
rect 9778 2868 9954 2870
rect 9996 2868 10130 2870
rect 10248 2868 10288 2972
rect 9778 2858 9956 2868
rect 9778 2682 9784 2858
rect 9818 2682 9914 2858
rect 9948 2682 9956 2858
rect 9778 2674 9956 2682
rect 9996 2858 10176 2868
rect 9996 2682 10002 2858
rect 10036 2856 10176 2858
rect 10036 2682 10136 2856
rect 9996 2680 10136 2682
rect 10170 2680 10176 2856
rect 9778 2672 9954 2674
rect 9778 2670 9824 2672
rect 9890 2670 9954 2672
rect 9996 2672 10176 2680
rect 9996 2670 10042 2672
rect 9562 2668 9722 2670
rect 9890 2668 9930 2670
rect 10130 2668 10176 2672
rect 10218 2856 10296 2868
rect 10218 2680 10224 2856
rect 10258 2790 10296 2856
rect 10284 2732 10296 2790
rect 10258 2680 10296 2732
rect 10218 2674 10296 2680
rect 10218 2668 10264 2674
rect 9802 2640 9854 2642
rect 9778 2636 10132 2640
rect 9778 2598 9808 2636
rect 9848 2632 10132 2636
rect 9848 2598 10086 2632
rect 10120 2598 10132 2632
rect 9778 2594 10132 2598
rect 9802 2592 9854 2594
rect 10076 2588 10132 2594
rect 5214 2152 5472 2162
rect 5214 2060 5240 2152
rect 5428 2122 5472 2152
rect 5428 2078 7492 2122
rect 5428 2060 5472 2078
rect 5214 2048 5472 2060
rect 5032 2022 5140 2042
rect 5032 1918 5050 2022
rect 5110 2014 5140 2022
rect 5110 2010 5686 2014
rect 5110 1968 6506 2010
rect 5110 1960 5686 1968
rect 5110 1918 5140 1960
rect 5032 1908 5140 1918
rect 5624 1832 6036 1906
rect 5624 1798 5786 1832
rect 5870 1798 6036 1832
rect 3436 1122 5006 1164
rect 3436 1098 3470 1122
rect 3280 1080 3470 1098
rect 5624 1054 6036 1798
rect 6468 1742 6506 1968
rect 4636 874 4864 916
rect 4636 742 4672 874
rect 4816 742 4864 874
rect 4636 710 4864 742
rect 1198 626 1622 628
rect 1198 606 2660 626
rect 1198 566 1612 606
rect 1810 604 2660 606
rect 1810 566 2223 604
rect 2427 566 2660 604
rect 1198 564 2660 566
rect 1470 560 2660 564
rect 1592 554 2660 560
rect -4320 344 -3008 538
rect -4320 -150 -4112 344
rect -3152 -150 -3008 344
rect -4320 -370 -3008 -150
rect 3102 160 4414 354
rect 3102 -334 3310 160
rect 4270 -334 4414 160
rect 3102 -554 4414 -334
rect 5624 -334 5682 1054
rect 5716 -334 5940 1054
rect 5974 -334 6036 1054
rect 6298 1716 6506 1742
rect 7450 1720 7492 2078
rect 7302 1716 7492 1720
rect 8214 1782 8626 1872
rect 8214 1748 8384 1782
rect 8468 1748 8626 1782
rect 6298 1698 6954 1716
rect 6298 1664 6336 1698
rect 6420 1664 6594 1698
rect 6678 1664 6852 1698
rect 6936 1664 6954 1698
rect 6298 1648 6954 1664
rect 7302 1698 7956 1716
rect 7302 1664 7336 1698
rect 7420 1664 7594 1698
rect 7678 1664 7852 1698
rect 7936 1664 7956 1698
rect 7302 1648 7956 1664
rect 6298 766 6476 1648
rect 6298 742 6956 766
rect 6298 708 6336 742
rect 6420 708 6594 742
rect 6678 708 6852 742
rect 6936 708 6956 742
rect 6298 698 6956 708
rect 7302 762 7480 1648
rect 8214 1004 8626 1748
rect 7302 742 7956 762
rect 7302 708 7336 742
rect 7420 708 7594 742
rect 7678 708 7852 742
rect 7936 708 7956 742
rect 6298 -188 6476 698
rect 7302 694 7956 708
rect 6298 -214 6958 -188
rect 6298 -248 6336 -214
rect 6420 -248 6594 -214
rect 6678 -248 6852 -214
rect 6936 -248 6958 -214
rect 6298 -256 6958 -248
rect 7302 -192 7480 694
rect 7302 -214 7956 -192
rect 7302 -248 7336 -214
rect 7420 -248 7594 -214
rect 7678 -248 7852 -214
rect 7936 -248 7956 -214
rect 6298 -282 6476 -256
rect 7302 -260 7956 -248
rect 7302 -304 7480 -260
rect 5624 -540 6036 -334
rect 8214 -384 8280 1004
rect 8314 -384 8538 1004
rect 8572 256 8626 1004
rect 9734 478 11046 672
rect 9734 256 9942 478
rect 8572 -16 9942 256
rect 10902 -16 11046 478
rect 8572 -60 11046 -16
rect 8572 -384 8626 -60
rect 9734 -236 11046 -60
rect 8214 -540 8626 -384
rect 5624 -604 8626 -540
rect 5624 -1118 6036 -604
rect 8214 -1152 8626 -604
<< via1 >>
rect 10364 10220 11324 10714
rect -2268 8770 -1836 8786
rect -2268 8732 -2250 8770
rect -2250 8732 -1853 8770
rect -1853 8732 -1836 8770
rect -2268 8716 -1836 8732
rect 2014 8770 2446 8786
rect 2014 8732 2031 8770
rect 2031 8732 2428 8770
rect 2428 8732 2446 8770
rect 2014 8716 2446 8732
rect 2928 8772 3362 8790
rect 2928 8734 2946 8772
rect 2946 8734 3343 8772
rect 3343 8734 3362 8772
rect 2928 8716 3362 8734
rect -2268 8452 -1836 8468
rect -2268 8414 -2250 8452
rect -2250 8414 -1853 8452
rect -1853 8414 -1836 8452
rect -2268 8398 -1836 8414
rect 2014 8452 2446 8468
rect 2014 8414 2031 8452
rect 2031 8414 2428 8452
rect 2428 8414 2446 8452
rect 2014 8398 2446 8414
rect -2268 8134 -1836 8150
rect -2268 8096 -2250 8134
rect -2250 8096 -1853 8134
rect -1853 8096 -1836 8134
rect -2268 8080 -1836 8096
rect 2928 8454 3362 8470
rect 2928 8416 2946 8454
rect 2946 8416 3343 8454
rect 3343 8416 3362 8454
rect 2928 8396 3362 8416
rect 7210 8772 7638 8788
rect 7210 8734 7227 8772
rect 7227 8734 7624 8772
rect 7624 8734 7638 8772
rect 7210 8718 7638 8734
rect 7212 8454 7640 8468
rect 7212 8416 7227 8454
rect 7227 8416 7624 8454
rect 7624 8416 7640 8454
rect 7212 8398 7640 8416
rect 2014 8134 2446 8150
rect 2014 8096 2031 8134
rect 2031 8096 2428 8134
rect 2428 8096 2446 8134
rect 2014 8080 2446 8096
rect 2926 8136 3360 8156
rect 2926 8098 2946 8136
rect 2946 8098 3343 8136
rect 3343 8098 3360 8136
rect 2926 8082 3360 8098
rect 7212 8136 7640 8152
rect 7212 8098 7227 8136
rect 7227 8098 7624 8136
rect 7624 8098 7640 8136
rect 7212 8082 7640 8098
rect -2268 7816 -1834 7832
rect -2268 7778 -2250 7816
rect -2250 7778 -1853 7816
rect -1853 7778 -1834 7816
rect -2268 7758 -1834 7778
rect -2270 7498 -1836 7516
rect -2270 7460 -2250 7498
rect -2250 7460 -1853 7498
rect -1853 7460 -1836 7498
rect -2270 7442 -1836 7460
rect 2014 7816 2446 7834
rect 2014 7778 2031 7816
rect 2031 7778 2428 7816
rect 2428 7778 2446 7816
rect 2014 7762 2446 7778
rect 2014 7498 2446 7516
rect 2014 7460 2031 7498
rect 2031 7460 2428 7498
rect 2428 7460 2446 7498
rect 2014 7444 2446 7460
rect -2268 7180 -1836 7196
rect -2268 7142 -2250 7180
rect -2250 7142 -1853 7180
rect -1853 7142 -1836 7180
rect -2268 7126 -1836 7142
rect 2928 7818 3360 7834
rect 2928 7780 2946 7818
rect 2946 7780 3343 7818
rect 3343 7780 3360 7818
rect 2928 7764 3360 7780
rect 7210 7818 7642 7834
rect 7210 7780 7227 7818
rect 7227 7780 7624 7818
rect 7624 7780 7642 7818
rect 7210 7764 7642 7780
rect 2928 7500 3360 7516
rect 2928 7462 2946 7500
rect 2946 7462 3343 7500
rect 3343 7462 3360 7500
rect 2928 7446 3360 7462
rect 7210 7500 7642 7516
rect 7210 7462 7227 7500
rect 7227 7462 7624 7500
rect 7624 7462 7642 7500
rect 7210 7446 7642 7462
rect 2014 7180 2446 7198
rect 2014 7142 2031 7180
rect 2031 7142 2428 7180
rect 2428 7142 2446 7180
rect 2014 7124 2446 7142
rect 2928 7182 3360 7198
rect 2928 7144 2946 7182
rect 2946 7144 3343 7182
rect 3343 7144 3360 7182
rect 2928 7128 3360 7144
rect 7210 7182 7642 7198
rect 7210 7144 7227 7182
rect 7227 7144 7624 7182
rect 7624 7144 7642 7182
rect 7210 7128 7642 7144
rect -2268 6862 -1842 6880
rect -2268 6824 -2250 6862
rect -2250 6824 -1853 6862
rect -1853 6824 -1842 6862
rect -2268 6808 -1842 6824
rect -2268 6544 -1842 6562
rect -2268 6506 -2250 6544
rect -2250 6506 -1853 6544
rect -1853 6506 -1842 6544
rect -2268 6490 -1842 6506
rect 2014 6862 2446 6878
rect 2014 6824 2031 6862
rect 2031 6824 2428 6862
rect 2428 6824 2446 6862
rect 2014 6806 2446 6824
rect 2926 6864 3364 6882
rect 2926 6826 2946 6864
rect 2946 6826 3343 6864
rect 3343 6826 3364 6864
rect 2926 6808 3364 6826
rect 7210 6864 7642 6880
rect 7210 6826 7227 6864
rect 7227 6826 7624 6864
rect 7624 6826 7642 6864
rect 7210 6810 7642 6826
rect 2014 6544 2446 6562
rect 2014 6506 2031 6544
rect 2031 6506 2428 6544
rect 2428 6506 2446 6544
rect 2014 6490 2446 6506
rect 2926 6546 3362 6564
rect 2926 6508 2946 6546
rect 2946 6508 3343 6546
rect 3343 6508 3362 6546
rect 2926 6494 3362 6508
rect -2268 6226 -1836 6244
rect -2268 6188 -2250 6226
rect -2250 6188 -1853 6226
rect -1853 6188 -1836 6226
rect -2268 6172 -1836 6188
rect 2016 6226 2444 6244
rect 2016 6188 2031 6226
rect 2031 6188 2428 6226
rect 2428 6188 2444 6226
rect 2016 6172 2444 6188
rect 2926 6228 3362 6244
rect 2926 6190 2946 6228
rect 2946 6190 3343 6228
rect 3343 6190 3362 6228
rect 2926 6174 3362 6190
rect 7210 6546 7646 6562
rect 7210 6508 7227 6546
rect 7227 6508 7624 6546
rect 7624 6508 7646 6546
rect 7210 6492 7646 6508
rect 7210 6228 7646 6244
rect 7210 6190 7227 6228
rect 7227 6190 7624 6228
rect 7624 6190 7646 6228
rect 7210 6174 7646 6190
rect -3704 5172 -3584 5250
rect -6262 4422 -5936 4662
rect -6648 3462 -6588 3526
rect -6250 3444 -6242 3508
rect -6242 3444 -6208 3508
rect -6208 3444 -6186 3508
rect -6144 3550 -6102 3620
rect -6102 3550 -6068 3620
rect -6068 3550 -6066 3620
rect -6020 3344 -6014 3410
rect -6014 3344 -5980 3410
rect -5980 3344 -5948 3410
rect -5800 3558 -5796 3624
rect -5796 3558 -5762 3624
rect -5762 3558 -5728 3624
rect -6568 2912 -6538 2970
rect -6538 2912 -6510 2970
rect -5792 2910 -5760 2968
rect -5760 2910 -5734 2968
rect -1374 4500 -1048 4740
rect -1462 3480 -1402 3544
rect -1064 3462 -1056 3526
rect -1056 3462 -1022 3526
rect -1022 3462 -1000 3526
rect -958 3568 -916 3638
rect -916 3568 -882 3638
rect -882 3568 -880 3638
rect -834 3362 -828 3428
rect -828 3362 -794 3428
rect -794 3362 -762 3428
rect -614 3576 -610 3642
rect -610 3576 -576 3642
rect -576 3576 -542 3642
rect -6 4952 46 5052
rect 174 4964 226 5048
rect 898 4972 976 5070
rect 2676 4966 2764 5098
rect 282 4712 458 4764
rect -180 4582 -72 4668
rect 5142 4752 5224 4838
rect 6582 4766 6642 4820
rect 7158 4822 7220 4882
rect 3938 4288 4264 4528
rect 3714 3492 3774 3556
rect -1382 2930 -1352 2988
rect -1352 2930 -1324 2988
rect -606 2928 -574 2986
rect -574 2928 -548 2986
rect 314 3054 420 3108
rect 4112 3474 4120 3538
rect 4120 3474 4154 3538
rect 4154 3474 4176 3538
rect 4218 3580 4260 3650
rect 4260 3580 4294 3650
rect 4294 3580 4296 3650
rect 4342 3374 4348 3440
rect 4348 3374 4382 3440
rect 4382 3374 4414 3440
rect 4562 3588 4566 3654
rect 4566 3588 4600 3654
rect 4600 3588 4634 3654
rect 3794 2942 3824 3000
rect 3824 2942 3852 3000
rect -5426 2458 -5350 2526
rect 4570 2940 4602 2998
rect 4602 2940 4628 2998
rect 3102 2362 3226 2414
rect 3092 1182 3210 1244
rect 9374 4230 9700 4470
rect 9028 3654 9110 3754
rect 9370 3284 9430 3348
rect 9768 3266 9776 3330
rect 9776 3266 9810 3330
rect 9810 3266 9832 3330
rect 9874 3372 9916 3442
rect 9916 3372 9950 3442
rect 9950 3372 9952 3442
rect 9998 3166 10004 3232
rect 10004 3166 10038 3232
rect 10038 3166 10070 3232
rect 10218 3380 10222 3446
rect 10222 3380 10256 3446
rect 10256 3380 10290 3446
rect 9450 2734 9480 2792
rect 9480 2734 9508 2792
rect 10226 2732 10258 2790
rect 10258 2732 10284 2790
rect 5240 2060 5428 2152
rect 4672 742 4816 874
rect -4112 -150 -3152 344
rect 3310 -334 4270 160
rect 9942 -16 10902 478
<< metal2 >>
rect 10156 10714 11468 10908
rect 1664 10456 1720 10466
rect 1660 10450 7194 10456
rect 10156 10450 10364 10714
rect 1660 10364 10364 10450
rect -2282 8786 -1832 8800
rect -2282 8716 -2268 8786
rect -1836 8716 -1832 8786
rect -2282 8468 -1832 8716
rect -2282 8398 -2268 8468
rect -1836 8398 -1832 8468
rect -2282 8388 -1832 8398
rect -2280 8154 -1826 8170
rect -2280 8080 -2268 8154
rect -1836 8080 -1826 8154
rect -2280 8064 -1826 8080
rect -2280 7834 -1820 7848
rect -2280 7758 -2268 7834
rect -1836 7832 -1820 7834
rect -1834 7758 -1820 7832
rect -2280 7516 -1820 7758
rect -2280 7442 -2270 7516
rect -2280 7440 -2268 7442
rect -1834 7440 -1820 7516
rect -2280 7428 -1820 7440
rect -2276 7202 -1828 7206
rect -3696 7196 -1828 7202
rect -3696 7126 -2268 7196
rect -1836 7126 -1828 7196
rect -3696 7114 -1828 7126
rect -3696 7112 -2090 7114
rect -3670 6934 -3614 7112
rect -3670 5280 -3618 6934
rect -2282 6882 -1832 6890
rect -2282 6880 -1830 6882
rect -2282 6808 -2268 6880
rect -1842 6808 -1830 6880
rect -2282 6644 -1830 6808
rect 1664 6708 1720 10364
rect 6850 10332 10364 10364
rect 2226 8868 6074 8906
rect 2226 8804 2276 8868
rect 2008 8786 2462 8804
rect 2008 8716 2014 8786
rect 2446 8716 2462 8786
rect 2008 8698 2462 8716
rect 2916 8790 3366 8800
rect 2916 8716 2928 8790
rect 3362 8716 3366 8790
rect 2006 8468 2462 8482
rect 2006 8398 2014 8468
rect 2446 8398 2462 8468
rect 2006 8150 2462 8398
rect 2916 8470 3366 8716
rect 2916 8396 2928 8470
rect 3362 8396 3366 8470
rect 2916 8384 3366 8396
rect 2006 8080 2014 8150
rect 2446 8080 2462 8150
rect 2006 8066 2462 8080
rect 2916 8156 3370 8166
rect 2916 8082 2926 8156
rect 3360 8082 3370 8156
rect 2916 8072 3370 8082
rect 3102 7978 3148 8072
rect 3102 7940 5184 7978
rect 2000 7834 2456 7852
rect 2000 7762 2014 7834
rect 2446 7762 2456 7834
rect 2000 7516 2456 7762
rect 2000 7444 2014 7516
rect 2446 7444 2456 7516
rect 2000 7198 2456 7444
rect 2918 7834 3364 7846
rect 2918 7764 2928 7834
rect 3360 7764 3364 7834
rect 2918 7516 3364 7764
rect 2918 7446 2928 7516
rect 3360 7446 3364 7516
rect 2918 7434 3364 7446
rect 2000 7124 2014 7198
rect 2446 7124 2456 7198
rect 2000 7112 2456 7124
rect 2918 7198 3366 7208
rect 2918 7128 2928 7198
rect 3360 7128 3366 7198
rect 2918 7118 3366 7128
rect 3134 7058 3200 7118
rect 4492 7058 4564 7064
rect 3134 6996 4564 7058
rect 3134 6994 3200 6996
rect 2010 6878 2456 6896
rect 2010 6806 2014 6878
rect 2446 6806 2456 6878
rect 2010 6708 2456 6806
rect 2920 6882 3374 6892
rect 2920 6808 2926 6882
rect 3364 6808 3374 6882
rect 2920 6798 3374 6808
rect 4 6644 40 6650
rect 1664 6648 2456 6708
rect 3182 6720 3220 6798
rect 3182 6672 4070 6720
rect -2282 6602 40 6644
rect -2282 6562 -1830 6602
rect -2282 6490 -2268 6562
rect -1842 6490 -1830 6562
rect -2282 6488 -1830 6490
rect -2282 6478 -1832 6488
rect -2276 6246 -1828 6256
rect -2518 6244 -1828 6246
rect -2518 6190 -2268 6244
rect -2518 5300 -2470 6190
rect -2276 6172 -2268 6190
rect -1836 6172 -1828 6244
rect -2276 6162 -1828 6172
rect -3726 5250 -3558 5280
rect -3726 5172 -3704 5250
rect -3584 5172 -3558 5250
rect -3726 5138 -3558 5172
rect -2524 4834 -2464 5300
rect 4 5072 40 6602
rect 2010 6562 2456 6648
rect 2010 6490 2014 6562
rect 2446 6490 2456 6562
rect 2010 6478 2456 6490
rect 2916 6564 3370 6580
rect 2916 6494 2926 6564
rect 3362 6494 3370 6564
rect 2916 6380 3370 6494
rect 170 6328 3370 6380
rect 170 6326 346 6328
rect 170 5072 234 6326
rect 2010 6244 2458 6254
rect 2010 6172 2016 6244
rect 2444 6172 2458 6244
rect 2010 6160 2458 6172
rect 2916 6244 3370 6328
rect 2916 6174 2926 6244
rect 3362 6174 3370 6244
rect 2158 6126 2214 6160
rect 2916 6154 3370 6174
rect 894 6090 2214 6126
rect 894 6086 2198 6090
rect 894 5090 950 6086
rect 2662 5098 2780 5124
rect -18 5052 58 5072
rect -18 4952 -6 5052
rect 46 4952 58 5052
rect -18 4932 58 4952
rect 158 5048 244 5072
rect 158 4964 174 5048
rect 226 4964 244 5048
rect 158 4940 244 4964
rect 886 5070 986 5090
rect 886 4972 898 5070
rect 976 4972 986 5070
rect 886 4940 986 4972
rect 2662 4966 2676 5098
rect 2764 5084 2780 5098
rect 4004 5084 4070 6672
rect 2764 5024 4070 5084
rect 2764 5018 4066 5024
rect 2764 4966 2780 5018
rect 2662 4946 2780 4966
rect -1468 4834 -954 4836
rect -2524 4800 -954 4834
rect -2522 4796 -954 4800
rect -6356 4662 -5842 4758
rect -6356 4422 -6262 4662
rect -5936 4422 -5842 4662
rect -6356 4324 -5842 4422
rect -1468 4740 -954 4796
rect 258 4764 490 4788
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect 58 4754 130 4756
rect 258 4754 282 4764
rect 58 4714 282 4754
rect -196 4668 -56 4686
rect -196 4582 -180 4668
rect -72 4582 -56 4668
rect -196 4562 -56 4582
rect -1468 4402 -954 4500
rect -176 4254 -72 4562
rect -6652 4202 -72 4254
rect -6652 3686 -6578 4202
rect 58 4056 130 4714
rect 258 4712 282 4714
rect 458 4712 490 4764
rect 258 4692 490 4712
rect 3844 4528 4358 4624
rect 3844 4288 3938 4528
rect 4264 4412 4358 4528
rect 4492 4412 4564 6996
rect 5142 4850 5184 7940
rect 5128 4838 5236 4850
rect 5128 4752 5142 4838
rect 5224 4752 5236 4838
rect 6034 4812 6074 8868
rect 6850 6386 6910 10332
rect 10156 10220 10364 10332
rect 11324 10220 11468 10714
rect 10156 10000 11468 10220
rect 7198 8788 7656 8800
rect 7198 8718 7210 8788
rect 7638 8718 7656 8788
rect 7198 8468 7656 8718
rect 7198 8398 7212 8468
rect 7640 8398 7656 8468
rect 7198 8298 7656 8398
rect 7198 8246 7658 8298
rect 7198 8152 7656 8246
rect 7198 8082 7212 8152
rect 7640 8082 7656 8152
rect 7198 8062 7656 8082
rect 7780 7846 7858 7848
rect 7508 7844 7858 7846
rect 7206 7834 7858 7844
rect 7206 7764 7210 7834
rect 7642 7764 7858 7834
rect 7206 7754 7858 7764
rect 7508 7750 7858 7754
rect 7206 7516 7652 7528
rect 7206 7446 7210 7516
rect 7642 7446 7652 7516
rect 7206 7198 7652 7446
rect 7206 7128 7210 7198
rect 7642 7128 7652 7198
rect 7206 7116 7652 7128
rect 7200 6880 7654 6892
rect 7200 6810 7210 6880
rect 7642 6810 7654 6880
rect 7200 6798 7654 6810
rect 7202 6562 7658 6576
rect 7202 6492 7210 6562
rect 7646 6492 7658 6562
rect 7202 6386 7658 6492
rect 6850 6308 7658 6386
rect 7202 6244 7658 6308
rect 7202 6174 7210 6244
rect 7646 6174 7658 6244
rect 7202 6158 7658 6174
rect 7780 4926 7858 7750
rect 7140 4882 7238 4900
rect 6560 4820 6658 4826
rect 6560 4812 6582 4820
rect 6034 4766 6582 4812
rect 6642 4766 6658 4820
rect 7140 4822 7158 4882
rect 7220 4860 7238 4882
rect 7778 4860 7860 4926
rect 7220 4838 7860 4860
rect 7220 4832 7858 4838
rect 7220 4822 7238 4832
rect 7140 4804 7238 4822
rect 6034 4764 6658 4766
rect 5128 4734 5236 4752
rect 6560 4750 6658 4764
rect 9280 4470 9794 4566
rect 4264 4336 4566 4412
rect 4264 4288 4358 4336
rect 4492 4330 4564 4336
rect 3844 4190 4358 4288
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
rect -5572 4000 130 4056
rect -6444 3686 -6390 3688
rect -6666 3680 -6390 3686
rect -6250 3682 -6180 3686
rect -6252 3680 -6180 3682
rect -6666 3526 -6180 3680
rect -6152 3624 -5724 3686
rect -5572 3624 -5496 4000
rect 58 3998 130 4000
rect 9002 3754 9140 3780
rect 3918 3716 3972 3718
rect 3696 3710 3972 3716
rect 4112 3712 4182 3716
rect 4110 3710 4182 3712
rect -1258 3704 -1204 3706
rect -6152 3620 -5800 3624
rect -6152 3550 -6144 3620
rect -6066 3558 -5800 3620
rect -5728 3558 -5496 3624
rect -6066 3556 -5496 3558
rect -6066 3550 -5724 3556
rect -5572 3552 -5496 3556
rect -1480 3698 -1204 3704
rect -1064 3700 -994 3704
rect -1066 3698 -994 3700
rect -6152 3532 -5724 3550
rect -6142 3530 -5724 3532
rect -1480 3544 -994 3698
rect -966 3642 -538 3704
rect -966 3638 -614 3642
rect -966 3568 -958 3638
rect -880 3576 -614 3638
rect -542 3576 -538 3642
rect -880 3568 -538 3576
rect -966 3550 -538 3568
rect -956 3548 -538 3550
rect 3696 3556 4182 3710
rect 4210 3654 4638 3716
rect 4210 3650 4562 3654
rect 4210 3580 4218 3650
rect 4296 3588 4562 3650
rect 4634 3588 4638 3654
rect 9002 3654 9028 3754
rect 9110 3654 9140 3754
rect 9002 3624 9140 3654
rect 4296 3580 4638 3588
rect 4210 3562 4638 3580
rect 4220 3560 4638 3562
rect 4254 3556 4608 3560
rect -922 3544 -568 3548
rect -6108 3526 -5754 3530
rect -6666 3462 -6648 3526
rect -6588 3508 -6180 3526
rect -6588 3462 -6250 3508
rect -6666 3444 -6250 3462
rect -6186 3444 -6180 3508
rect -6666 3286 -6180 3444
rect -1480 3480 -1462 3544
rect -1402 3526 -994 3544
rect -1402 3480 -1064 3526
rect -1480 3462 -1064 3480
rect -1000 3462 -994 3526
rect -5622 3420 -5568 3426
rect -6030 3410 -5568 3420
rect -6030 3344 -6020 3410
rect -5948 3344 -5568 3410
rect -6030 3334 -5568 3344
rect -6666 3284 -6426 3286
rect -6394 3284 -6180 3286
rect -6252 3282 -6180 3284
rect -6586 2970 -5724 3048
rect -6586 2912 -6568 2970
rect -6510 2968 -5724 2970
rect -6510 2912 -5792 2968
rect -6586 2910 -5792 2912
rect -5734 2910 -5724 2968
rect -6586 2846 -5724 2910
rect -5622 2512 -5568 3334
rect -1480 3304 -994 3462
rect 3696 3492 3714 3556
rect 3774 3538 4182 3556
rect 3774 3492 4112 3538
rect 3696 3474 4112 3492
rect 4176 3474 4182 3538
rect 9574 3508 9628 3510
rect -844 3428 -384 3438
rect -844 3362 -834 3428
rect -762 3418 -384 3428
rect 64 3418 110 3422
rect -762 3378 110 3418
rect -762 3362 -384 3378
rect -844 3352 -384 3362
rect -1480 3302 -1240 3304
rect -1208 3302 -994 3304
rect -1066 3300 -994 3302
rect 64 3100 110 3378
rect 3696 3316 4182 3474
rect 9352 3502 9628 3508
rect 9768 3504 9838 3508
rect 9766 3502 9838 3504
rect 4738 3450 4796 3452
rect 4332 3440 4796 3450
rect 4332 3374 4342 3440
rect 4414 3374 4796 3440
rect 4332 3364 4796 3374
rect 3696 3314 3936 3316
rect 3968 3314 4182 3316
rect 4110 3312 4182 3314
rect 288 3108 446 3120
rect 288 3100 314 3108
rect 64 3066 314 3100
rect -1400 2988 -538 3066
rect 66 3060 314 3066
rect 288 3054 314 3060
rect 420 3054 446 3108
rect 288 3040 446 3054
rect -1400 2930 -1382 2988
rect -1324 2986 -538 2988
rect -1324 2930 -606 2986
rect -1400 2928 -606 2930
rect -548 2928 -538 2986
rect -1400 2864 -538 2928
rect 3776 3000 4638 3078
rect 3776 2942 3794 3000
rect 3852 2998 4638 3000
rect 3852 2942 4570 2998
rect 3776 2940 4570 2942
rect 4628 2940 4638 2998
rect 3776 2876 4638 2940
rect 4738 2690 4796 3364
rect 9352 3348 9838 3502
rect 9866 3446 10294 3508
rect 9866 3442 10218 3446
rect 9866 3372 9874 3442
rect 9952 3380 10218 3442
rect 10290 3380 10294 3446
rect 9952 3372 10294 3380
rect 9866 3354 10294 3372
rect 9876 3352 10294 3354
rect 9910 3348 10264 3352
rect 9352 3284 9370 3348
rect 9430 3330 9838 3348
rect 9430 3284 9768 3330
rect 9352 3266 9768 3284
rect 9832 3266 9838 3330
rect 9352 3108 9838 3266
rect 9988 3232 10448 3242
rect 9988 3166 9998 3232
rect 10070 3166 10448 3232
rect 9988 3156 10448 3166
rect 9352 3106 9592 3108
rect 9624 3106 9838 3108
rect 9766 3104 9838 3106
rect 9432 2792 10294 2870
rect 9432 2734 9450 2792
rect 9508 2790 10294 2792
rect 9508 2734 10226 2790
rect 9432 2732 10226 2734
rect 10284 2732 10294 2790
rect -5446 2526 -5326 2548
rect -5446 2512 -5426 2526
rect -5622 2470 -5426 2512
rect -5620 2462 -5426 2470
rect -5446 2458 -5426 2462
rect -5350 2458 -5326 2526
rect -5446 2432 -5326 2458
rect 3076 2418 3252 2432
rect 3076 2362 3102 2418
rect 3226 2362 3252 2418
rect 3076 2344 3252 2362
rect 4740 2122 4792 2690
rect 9432 2668 10294 2732
rect 8592 2450 8812 2488
rect 8592 2332 8620 2450
rect 8778 2412 8812 2450
rect 10394 2412 10446 3156
rect 8778 2344 10448 2412
rect 8778 2332 8812 2344
rect 8592 2302 8812 2332
rect 5214 2152 5472 2162
rect 5214 2122 5240 2152
rect 4738 2068 5240 2122
rect 3078 1244 3224 1254
rect 3078 1182 3092 1244
rect 3210 1182 3224 1244
rect 3078 1170 3224 1182
rect 4740 916 4792 2068
rect 5214 2060 5240 2068
rect 5428 2060 5472 2152
rect 5214 2048 5472 2060
rect 4636 874 4864 916
rect 4636 742 4672 874
rect 4816 742 4864 874
rect 4636 710 4864 742
rect -4320 344 -3008 538
rect 9734 478 11046 672
rect -4320 -150 -4112 344
rect -3152 -150 -3008 344
rect -4320 -370 -3008 -150
rect 3102 160 4414 354
rect 3102 -334 3310 160
rect 4270 -334 4414 160
rect 9734 -16 9942 478
rect 10902 -16 11046 478
rect 9734 -236 11046 -16
rect 3102 -554 4414 -334
<< via2 >>
rect -2268 8150 -1836 8154
rect -2268 8080 -1836 8150
rect -2268 7832 -1836 7834
rect -2268 7760 -1836 7832
rect -2268 7442 -1836 7516
rect -1836 7442 -1834 7516
rect -2268 7440 -1834 7442
rect 2928 8718 3360 8790
rect 2928 8398 3360 8470
rect -6262 4422 -5936 4662
rect -1374 4500 -1048 4740
rect 3938 4288 4264 4528
rect 10364 10220 11324 10714
rect 7210 6810 7642 6880
rect 9374 4230 9700 4470
rect 9028 3654 9110 3754
rect 3102 2414 3226 2418
rect 3102 2362 3226 2414
rect 8620 2332 8778 2450
rect 3092 1182 3210 1244
rect -4112 -150 -3152 344
rect 3310 -334 4270 160
rect 9942 -16 10902 478
<< metal3 >>
rect 10156 10714 11468 10908
rect 2672 10434 2758 10480
rect 10156 10434 10364 10714
rect 2672 10350 10364 10434
rect 2672 8626 2758 10350
rect 10156 10220 10364 10350
rect 11324 10220 11468 10714
rect 10156 10000 11468 10220
rect 2914 8790 3368 8804
rect 2914 8718 2928 8790
rect 3360 8718 3368 8790
rect 2914 8626 3368 8718
rect 2672 8554 3368 8626
rect 2914 8470 3368 8554
rect 2914 8398 2928 8470
rect 3360 8398 3368 8470
rect 2914 8382 3368 8398
rect -2282 8154 -1824 8172
rect -2282 8080 -2268 8154
rect -1836 8080 -1824 8154
rect -2282 8062 -1824 8080
rect -2138 7992 -2072 8062
rect -2138 7924 -1248 7992
rect -2282 7834 -1822 7848
rect -2282 7760 -2268 7834
rect -1836 7760 -1822 7834
rect -2282 7640 -1822 7760
rect -1312 7640 -1248 7924
rect -2282 7576 -1240 7640
rect -2282 7516 -1822 7576
rect -2282 7440 -2268 7516
rect -1834 7440 -1822 7516
rect -2282 7422 -1822 7440
rect -1306 4836 -1240 7576
rect 7200 6884 7654 6894
rect 9448 6884 9510 6886
rect 7200 6880 9570 6884
rect 7200 6810 7210 6880
rect 7642 6810 9570 6880
rect 7200 6808 9570 6810
rect 7200 6798 7654 6808
rect -6356 4662 -5842 4758
rect -6356 4422 -6262 4662
rect -5936 4422 -5842 4662
rect -6356 4324 -5842 4422
rect -1468 4740 -954 4836
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect -1468 4402 -954 4500
rect 3844 4528 4358 4624
rect 9448 4566 9510 6808
rect 3844 4288 3938 4528
rect 4264 4288 4358 4528
rect 3844 4190 4358 4288
rect 9280 4470 9794 4566
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
rect 9002 3754 9140 3782
rect 9002 3654 9028 3754
rect 9110 3654 9140 3754
rect 9002 3624 9140 3654
rect 8592 2450 8812 2488
rect 3076 2418 3252 2432
rect 3076 2362 3102 2418
rect 3226 2408 3252 2418
rect 8592 2408 8620 2450
rect 3226 2362 8620 2408
rect 3076 2344 8620 2362
rect 8592 2332 8620 2344
rect 8778 2332 8812 2450
rect 8592 2302 8812 2332
rect 9040 1280 9106 3624
rect 8882 1278 9156 1280
rect 3118 1254 9156 1278
rect 3078 1244 9156 1254
rect 3078 1182 3092 1244
rect 3210 1192 9156 1244
rect 3210 1182 3224 1192
rect 8882 1190 9156 1192
rect 3078 1170 3224 1182
rect -4320 344 -3008 538
rect 9734 478 11046 672
rect -4320 -150 -4112 344
rect -3152 -150 -3008 344
rect -4320 -370 -3008 -150
rect 3102 160 4414 354
rect 3102 -334 3310 160
rect 4270 -334 4414 160
rect 9734 -16 9942 478
rect 10902 -16 11046 478
rect 9734 -236 11046 -16
rect 3102 -554 4414 -334
<< via3 >>
rect 10364 10220 11324 10714
rect -6262 4422 -5936 4662
rect -1374 4500 -1048 4740
rect 3938 4288 4264 4528
rect 9374 4230 9700 4470
rect -4112 -150 -3152 344
rect 3310 -334 4270 160
rect 9942 -16 10902 478
<< metal4 >>
rect 10156 10714 11468 10908
rect 10156 10474 10364 10714
rect 10150 10220 10364 10474
rect 11324 10220 11468 10714
rect 10150 10180 11468 10220
rect 10156 10000 11468 10180
rect -6356 4662 -5842 4758
rect -6356 4422 -6262 4662
rect -5936 4422 -5842 4662
rect -6356 4324 -5842 4422
rect -1468 4740 -954 4836
rect -1468 4500 -1374 4740
rect -1048 4500 -954 4740
rect -1468 4402 -954 4500
rect 3844 4528 4358 4624
rect 3844 4288 3938 4528
rect 4264 4288 4358 4528
rect 3844 4190 4358 4288
rect 9280 4470 9794 4566
rect 9280 4230 9374 4470
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
rect 10686 672 11034 10000
rect -4320 344 -3008 538
rect 9734 478 11046 672
rect -4320 -150 -4112 344
rect -3152 238 -3008 344
rect 3102 238 4414 354
rect 9734 238 9942 478
rect -3152 160 9942 238
rect -3152 -56 3310 160
rect -3152 -150 -3008 -56
rect -4320 -370 -3008 -150
rect 3102 -334 3310 -56
rect 4270 -16 9942 160
rect 10902 -16 11046 478
rect 4270 -56 11046 -16
rect 4270 -334 4414 -56
rect 9734 -236 11046 -56
rect 3102 -554 4414 -334
<< via4 >>
rect -6262 4422 -5936 4662
rect -1374 4500 -1048 4740
rect 3938 4288 4264 4528
rect 9374 4230 9700 4470
<< metal5 >>
rect -6356 4744 -5842 4758
rect -1468 4744 -954 4836
rect -6356 4740 9598 4744
rect -6356 4662 -1374 4740
rect -6356 4422 -6262 4662
rect -5936 4500 -1374 4662
rect -1048 4566 9598 4740
rect -1048 4528 9794 4566
rect -1048 4500 3938 4528
rect -5936 4422 3938 4500
rect -6356 4370 3938 4422
rect -6356 4324 -5842 4370
rect 3844 4288 3938 4370
rect 4264 4470 9794 4528
rect 4264 4370 9374 4470
rect 4264 4288 4358 4370
rect 3844 4190 4358 4288
rect 9280 4230 9374 4370
rect 9700 4230 9794 4470
rect 9280 4132 9794 4230
<< res0p35 >>
rect -7082 9376 -3228 9450
rect -1852 9376 2002 9450
rect 3378 9376 7232 9450
rect 8608 9376 12462 9450
rect -7082 9056 -3228 9130
rect -1852 9056 2002 9130
rect 3378 9056 7232 9130
rect 8608 9056 12462 9130
rect -7082 8736 -3228 8810
rect -1838 8714 2016 8788
rect 3358 8716 7212 8790
rect 8608 8736 12462 8810
rect -7082 8416 -3228 8490
rect -1838 8396 2016 8470
rect 3358 8398 7212 8472
rect 8608 8416 12462 8490
rect -7082 8096 -3228 8170
rect -1838 8078 2016 8152
rect 3358 8080 7212 8154
rect 8608 8096 12462 8170
rect -7082 7776 -3228 7850
rect -1838 7760 2016 7834
rect 3358 7762 7212 7836
rect 8608 7776 12462 7850
rect -7082 7456 -3228 7530
rect -1838 7442 2016 7516
rect 3358 7444 7212 7518
rect 8608 7456 12462 7530
rect -7082 7136 -3228 7210
rect -1838 7124 2016 7198
rect 3358 7126 7212 7200
rect 8608 7136 12462 7210
rect -7082 6816 -3228 6890
rect -1838 6806 2016 6880
rect 3358 6808 7212 6882
rect 8608 6816 12462 6890
rect -7082 6496 -3228 6570
rect -1838 6488 2016 6562
rect 3358 6490 7212 6564
rect 8608 6496 12462 6570
rect -7082 6176 -3228 6250
rect -1838 6170 2016 6244
rect 3358 6172 7212 6246
rect 8608 6176 12462 6250
rect -7082 5856 -3228 5930
rect -1818 5824 2036 5898
rect 3378 5854 7232 5928
rect 8608 5856 12462 5930
rect -7082 5536 -3228 5610
rect -1818 5504 2036 5578
rect 3378 5536 7232 5610
rect 8608 5536 12462 5610
<< labels >>
flabel metal4 -852 46 -852 46 0 FreeSans 1600 0 0 0 GND
flabel metal5 -5546 4550 -5546 4550 0 FreeSans 1600 0 0 0 VDD
flabel metal1 -86 3610 -86 3610 0 FreeSans 800 0 0 0 vinp1
flabel metal1 -170 2962 -170 2962 0 FreeSans 800 0 0 0 vinpch2
flabel metal2 -524 4224 -524 4226 0 FreeSans 800 0 0 0 outp1
flabel metal2 -538 4024 -538 4026 0 FreeSans 800 0 0 0 outp2
flabel locali 2688 2580 2688 2580 0 FreeSans 800 0 0 0 Bout
flabel locali 1512 2618 1512 2618 0 FreeSans 800 0 0 0 Bout_mirror
flabel metal3 3912 1244 3912 1244 0 FreeSans 800 0 0 0 outn1
flabel metal3 3872 2382 3872 2382 0 FreeSans 800 0 0 0 outn2
flabel locali 3568 1754 3568 1754 0 FreeSans 800 0 0 0 vinn1
flabel locali 3716 1850 3716 1850 0 FreeSans 800 0 0 0 vinnch1
flabel locali 3952 792 3952 792 0 FreeSans 800 0 0 0 vinnch2
flabel metal1 3994 1136 3994 1136 0 FreeSans 800 0 0 0 vinn2
flabel locali -3668 2058 -3668 2058 0 FreeSans 800 0 0 0 outpch1
flabel locali -2692 2038 -2692 2038 0 FreeSans 800 0 0 0 outpch2
flabel metal1 6856 4786 6856 4786 0 FreeSans 800 0 0 0 vbiasob
flabel metal1 -2036 1542 -2036 1542 0 FreeSans 800 0 0 0 vbiasot
flabel locali 3806 3846 3806 3846 0 FreeSans 400 0 0 0 Fvco_By4_QPH_bar
flabel locali -1416 3844 -1416 3844 0 FreeSans 400 0 0 0 Fvco_By4_QPH_bar
flabel locali -6684 3828 -6684 3828 0 FreeSans 400 0 0 0 Fvco_By4_QPH_bar
flabel locali -6606 3106 -6606 3106 0 FreeSans 400 0 0 0 Fvco_By4_QPH
flabel locali -1450 3118 -1450 3118 0 FreeSans 400 0 0 0 Fvco_By4_QPH
flabel locali 3812 3134 3812 3134 0 FreeSans 400 0 0 0 Fvco_By4_QPH
flabel locali 7022 2640 7022 2640 0 FreeSans 400 0 0 0 outnch1
flabel locali 7628 2648 7628 2648 0 FreeSans 400 0 0 0 outnch2
flabel metal1 -112 2610 -112 2610 0 FreeSans 400 0 0 0 vinp2
flabel metal2 -176 3408 -176 3408 0 FreeSans 400 0 0 0 vinpch1
flabel metal1 3118 4336 3118 4336 0 FreeSans 400 0 0 0 vbiaschopper
flabel locali 9446 3650 9446 3650 0 FreeSans 400 0 0 0 Fvco_By4_QPH
flabel locali 9416 2918 9416 2918 0 FreeSans 400 0 0 0 Fvco_By4_QPH_bar
<< end >>
