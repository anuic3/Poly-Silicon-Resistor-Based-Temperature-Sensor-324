magic
tech sky130A
magscale 1 2
timestamp 1634377750
<< nwell >>
rect -38 261 42358 621
<< pwell >>
rect 903 157 1089 201
rect 1633 157 2104 203
rect 3019 157 3205 201
rect 3749 157 4220 203
rect 5135 157 5321 201
rect 5865 157 6336 203
rect 7251 157 7437 201
rect 7981 157 8452 203
rect 9367 157 9553 201
rect 10097 157 10568 203
rect 11483 157 11669 201
rect 12213 157 12684 203
rect 13599 157 13785 201
rect 14329 157 14800 203
rect 15715 157 15901 201
rect 16445 157 16916 203
rect 17831 157 18017 201
rect 18561 157 19032 203
rect 19947 157 20133 201
rect 20677 157 21148 203
rect 22063 157 22249 201
rect 22793 157 23264 203
rect 24179 157 24365 201
rect 24909 157 25380 203
rect 26295 157 26481 201
rect 27025 157 27496 203
rect 28411 157 28597 201
rect 29141 157 29612 203
rect 30527 157 30713 201
rect 31257 157 31728 203
rect 32643 157 32829 201
rect 33373 157 33844 203
rect 34759 157 34945 201
rect 35489 157 35960 203
rect 36875 157 37061 201
rect 37605 157 38076 203
rect 38991 157 39177 201
rect 39721 157 40192 203
rect 41107 157 41293 201
rect 41837 157 42308 203
rect 1 48 2104 157
rect 2117 48 4220 157
rect 4233 48 6336 157
rect 6349 48 8452 157
rect 8465 48 10568 157
rect 10581 48 12684 157
rect 12697 48 14800 157
rect 14813 48 16916 157
rect 16929 48 19032 157
rect 19045 48 21148 157
rect 21161 48 23264 157
rect 23277 48 25380 157
rect 25393 48 27496 157
rect 27509 48 29612 157
rect 29625 48 31728 157
rect 31741 48 33844 157
rect 33857 48 35960 157
rect 35973 48 38076 157
rect 38089 48 40192 157
rect 40205 48 42308 157
rect 0 -77 42320 48
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 418 47 448 131
rect 513 47 543 119
rect 609 47 639 119
rect 775 47 805 131
rect 847 47 877 131
rect 979 47 1009 175
rect 1078 47 1108 119
rect 1187 47 1217 119
rect 1283 47 1313 131
rect 1432 47 1462 131
rect 1523 47 1553 131
rect 1711 47 1741 177
rect 1899 47 1929 131
rect 1996 47 2026 177
rect 2195 47 2225 131
rect 2279 47 2309 131
rect 2534 47 2564 131
rect 2629 47 2659 119
rect 2725 47 2755 119
rect 2891 47 2921 131
rect 2963 47 2993 131
rect 3095 47 3125 175
rect 3194 47 3224 119
rect 3303 47 3333 119
rect 3399 47 3429 131
rect 3548 47 3578 131
rect 3639 47 3669 131
rect 3827 47 3857 177
rect 4015 47 4045 131
rect 4112 47 4142 177
rect 4311 47 4341 131
rect 4395 47 4425 131
rect 4650 47 4680 131
rect 4745 47 4775 119
rect 4841 47 4871 119
rect 5007 47 5037 131
rect 5079 47 5109 131
rect 5211 47 5241 175
rect 5310 47 5340 119
rect 5419 47 5449 119
rect 5515 47 5545 131
rect 5664 47 5694 131
rect 5755 47 5785 131
rect 5943 47 5973 177
rect 6131 47 6161 131
rect 6228 47 6258 177
rect 6427 47 6457 131
rect 6511 47 6541 131
rect 6766 47 6796 131
rect 6861 47 6891 119
rect 6957 47 6987 119
rect 7123 47 7153 131
rect 7195 47 7225 131
rect 7327 47 7357 175
rect 7426 47 7456 119
rect 7535 47 7565 119
rect 7631 47 7661 131
rect 7780 47 7810 131
rect 7871 47 7901 131
rect 8059 47 8089 177
rect 8247 47 8277 131
rect 8344 47 8374 177
rect 8543 47 8573 131
rect 8627 47 8657 131
rect 8882 47 8912 131
rect 8977 47 9007 119
rect 9073 47 9103 119
rect 9239 47 9269 131
rect 9311 47 9341 131
rect 9443 47 9473 175
rect 9542 47 9572 119
rect 9651 47 9681 119
rect 9747 47 9777 131
rect 9896 47 9926 131
rect 9987 47 10017 131
rect 10175 47 10205 177
rect 10363 47 10393 131
rect 10460 47 10490 177
rect 10659 47 10689 131
rect 10743 47 10773 131
rect 10998 47 11028 131
rect 11093 47 11123 119
rect 11189 47 11219 119
rect 11355 47 11385 131
rect 11427 47 11457 131
rect 11559 47 11589 175
rect 11658 47 11688 119
rect 11767 47 11797 119
rect 11863 47 11893 131
rect 12012 47 12042 131
rect 12103 47 12133 131
rect 12291 47 12321 177
rect 12479 47 12509 131
rect 12576 47 12606 177
rect 12775 47 12805 131
rect 12859 47 12889 131
rect 13114 47 13144 131
rect 13209 47 13239 119
rect 13305 47 13335 119
rect 13471 47 13501 131
rect 13543 47 13573 131
rect 13675 47 13705 175
rect 13774 47 13804 119
rect 13883 47 13913 119
rect 13979 47 14009 131
rect 14128 47 14158 131
rect 14219 47 14249 131
rect 14407 47 14437 177
rect 14595 47 14625 131
rect 14692 47 14722 177
rect 14891 47 14921 131
rect 14975 47 15005 131
rect 15230 47 15260 131
rect 15325 47 15355 119
rect 15421 47 15451 119
rect 15587 47 15617 131
rect 15659 47 15689 131
rect 15791 47 15821 175
rect 15890 47 15920 119
rect 15999 47 16029 119
rect 16095 47 16125 131
rect 16244 47 16274 131
rect 16335 47 16365 131
rect 16523 47 16553 177
rect 16711 47 16741 131
rect 16808 47 16838 177
rect 17007 47 17037 131
rect 17091 47 17121 131
rect 17346 47 17376 131
rect 17441 47 17471 119
rect 17537 47 17567 119
rect 17703 47 17733 131
rect 17775 47 17805 131
rect 17907 47 17937 175
rect 18006 47 18036 119
rect 18115 47 18145 119
rect 18211 47 18241 131
rect 18360 47 18390 131
rect 18451 47 18481 131
rect 18639 47 18669 177
rect 18827 47 18857 131
rect 18924 47 18954 177
rect 19123 47 19153 131
rect 19207 47 19237 131
rect 19462 47 19492 131
rect 19557 47 19587 119
rect 19653 47 19683 119
rect 19819 47 19849 131
rect 19891 47 19921 131
rect 20023 47 20053 175
rect 20122 47 20152 119
rect 20231 47 20261 119
rect 20327 47 20357 131
rect 20476 47 20506 131
rect 20567 47 20597 131
rect 20755 47 20785 177
rect 20943 47 20973 131
rect 21040 47 21070 177
rect 21239 47 21269 131
rect 21323 47 21353 131
rect 21578 47 21608 131
rect 21673 47 21703 119
rect 21769 47 21799 119
rect 21935 47 21965 131
rect 22007 47 22037 131
rect 22139 47 22169 175
rect 22238 47 22268 119
rect 22347 47 22377 119
rect 22443 47 22473 131
rect 22592 47 22622 131
rect 22683 47 22713 131
rect 22871 47 22901 177
rect 23059 47 23089 131
rect 23156 47 23186 177
rect 23355 47 23385 131
rect 23439 47 23469 131
rect 23694 47 23724 131
rect 23789 47 23819 119
rect 23885 47 23915 119
rect 24051 47 24081 131
rect 24123 47 24153 131
rect 24255 47 24285 175
rect 24354 47 24384 119
rect 24463 47 24493 119
rect 24559 47 24589 131
rect 24708 47 24738 131
rect 24799 47 24829 131
rect 24987 47 25017 177
rect 25175 47 25205 131
rect 25272 47 25302 177
rect 25471 47 25501 131
rect 25555 47 25585 131
rect 25810 47 25840 131
rect 25905 47 25935 119
rect 26001 47 26031 119
rect 26167 47 26197 131
rect 26239 47 26269 131
rect 26371 47 26401 175
rect 26470 47 26500 119
rect 26579 47 26609 119
rect 26675 47 26705 131
rect 26824 47 26854 131
rect 26915 47 26945 131
rect 27103 47 27133 177
rect 27291 47 27321 131
rect 27388 47 27418 177
rect 27587 47 27617 131
rect 27671 47 27701 131
rect 27926 47 27956 131
rect 28021 47 28051 119
rect 28117 47 28147 119
rect 28283 47 28313 131
rect 28355 47 28385 131
rect 28487 47 28517 175
rect 28586 47 28616 119
rect 28695 47 28725 119
rect 28791 47 28821 131
rect 28940 47 28970 131
rect 29031 47 29061 131
rect 29219 47 29249 177
rect 29407 47 29437 131
rect 29504 47 29534 177
rect 29703 47 29733 131
rect 29787 47 29817 131
rect 30042 47 30072 131
rect 30137 47 30167 119
rect 30233 47 30263 119
rect 30399 47 30429 131
rect 30471 47 30501 131
rect 30603 47 30633 175
rect 30702 47 30732 119
rect 30811 47 30841 119
rect 30907 47 30937 131
rect 31056 47 31086 131
rect 31147 47 31177 131
rect 31335 47 31365 177
rect 31523 47 31553 131
rect 31620 47 31650 177
rect 31819 47 31849 131
rect 31903 47 31933 131
rect 32158 47 32188 131
rect 32253 47 32283 119
rect 32349 47 32379 119
rect 32515 47 32545 131
rect 32587 47 32617 131
rect 32719 47 32749 175
rect 32818 47 32848 119
rect 32927 47 32957 119
rect 33023 47 33053 131
rect 33172 47 33202 131
rect 33263 47 33293 131
rect 33451 47 33481 177
rect 33639 47 33669 131
rect 33736 47 33766 177
rect 33935 47 33965 131
rect 34019 47 34049 131
rect 34274 47 34304 131
rect 34369 47 34399 119
rect 34465 47 34495 119
rect 34631 47 34661 131
rect 34703 47 34733 131
rect 34835 47 34865 175
rect 34934 47 34964 119
rect 35043 47 35073 119
rect 35139 47 35169 131
rect 35288 47 35318 131
rect 35379 47 35409 131
rect 35567 47 35597 177
rect 35755 47 35785 131
rect 35852 47 35882 177
rect 36051 47 36081 131
rect 36135 47 36165 131
rect 36390 47 36420 131
rect 36485 47 36515 119
rect 36581 47 36611 119
rect 36747 47 36777 131
rect 36819 47 36849 131
rect 36951 47 36981 175
rect 37050 47 37080 119
rect 37159 47 37189 119
rect 37255 47 37285 131
rect 37404 47 37434 131
rect 37495 47 37525 131
rect 37683 47 37713 177
rect 37871 47 37901 131
rect 37968 47 37998 177
rect 38167 47 38197 131
rect 38251 47 38281 131
rect 38506 47 38536 131
rect 38601 47 38631 119
rect 38697 47 38727 119
rect 38863 47 38893 131
rect 38935 47 38965 131
rect 39067 47 39097 175
rect 39166 47 39196 119
rect 39275 47 39305 119
rect 39371 47 39401 131
rect 39520 47 39550 131
rect 39611 47 39641 131
rect 39799 47 39829 177
rect 39987 47 40017 131
rect 40084 47 40114 177
rect 40283 47 40313 131
rect 40367 47 40397 131
rect 40622 47 40652 131
rect 40717 47 40747 119
rect 40813 47 40843 119
rect 40979 47 41009 131
rect 41051 47 41081 131
rect 41183 47 41213 175
rect 41282 47 41312 119
rect 41391 47 41421 119
rect 41487 47 41517 131
rect 41636 47 41666 131
rect 41727 47 41757 131
rect 41915 47 41945 177
rect 42103 47 42133 131
rect 42200 47 42230 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 430 413 460 497
rect 522 413 552 497
rect 621 413 651 497
rect 761 413 791 497
rect 858 413 888 497
rect 1055 329 1085 497
rect 1154 413 1184 497
rect 1240 413 1270 497
rect 1324 413 1354 497
rect 1432 413 1462 497
rect 1516 413 1546 497
rect 1680 297 1710 497
rect 1899 369 1929 497
rect 1996 297 2026 497
rect 2195 363 2225 491
rect 2279 363 2309 491
rect 2546 413 2576 497
rect 2638 413 2668 497
rect 2737 413 2767 497
rect 2877 413 2907 497
rect 2974 413 3004 497
rect 3171 329 3201 497
rect 3270 413 3300 497
rect 3356 413 3386 497
rect 3440 413 3470 497
rect 3548 413 3578 497
rect 3632 413 3662 497
rect 3796 297 3826 497
rect 4015 369 4045 497
rect 4112 297 4142 497
rect 4311 363 4341 491
rect 4395 363 4425 491
rect 4662 413 4692 497
rect 4754 413 4784 497
rect 4853 413 4883 497
rect 4993 413 5023 497
rect 5090 413 5120 497
rect 5287 329 5317 497
rect 5386 413 5416 497
rect 5472 413 5502 497
rect 5556 413 5586 497
rect 5664 413 5694 497
rect 5748 413 5778 497
rect 5912 297 5942 497
rect 6131 369 6161 497
rect 6228 297 6258 497
rect 6427 363 6457 491
rect 6511 363 6541 491
rect 6778 413 6808 497
rect 6870 413 6900 497
rect 6969 413 6999 497
rect 7109 413 7139 497
rect 7206 413 7236 497
rect 7403 329 7433 497
rect 7502 413 7532 497
rect 7588 413 7618 497
rect 7672 413 7702 497
rect 7780 413 7810 497
rect 7864 413 7894 497
rect 8028 297 8058 497
rect 8247 369 8277 497
rect 8344 297 8374 497
rect 8543 363 8573 491
rect 8627 363 8657 491
rect 8894 413 8924 497
rect 8986 413 9016 497
rect 9085 413 9115 497
rect 9225 413 9255 497
rect 9322 413 9352 497
rect 9519 329 9549 497
rect 9618 413 9648 497
rect 9704 413 9734 497
rect 9788 413 9818 497
rect 9896 413 9926 497
rect 9980 413 10010 497
rect 10144 297 10174 497
rect 10363 369 10393 497
rect 10460 297 10490 497
rect 10659 363 10689 491
rect 10743 363 10773 491
rect 11010 413 11040 497
rect 11102 413 11132 497
rect 11201 413 11231 497
rect 11341 413 11371 497
rect 11438 413 11468 497
rect 11635 329 11665 497
rect 11734 413 11764 497
rect 11820 413 11850 497
rect 11904 413 11934 497
rect 12012 413 12042 497
rect 12096 413 12126 497
rect 12260 297 12290 497
rect 12479 369 12509 497
rect 12576 297 12606 497
rect 12775 363 12805 491
rect 12859 363 12889 491
rect 13126 413 13156 497
rect 13218 413 13248 497
rect 13317 413 13347 497
rect 13457 413 13487 497
rect 13554 413 13584 497
rect 13751 329 13781 497
rect 13850 413 13880 497
rect 13936 413 13966 497
rect 14020 413 14050 497
rect 14128 413 14158 497
rect 14212 413 14242 497
rect 14376 297 14406 497
rect 14595 369 14625 497
rect 14692 297 14722 497
rect 14891 363 14921 491
rect 14975 363 15005 491
rect 15242 413 15272 497
rect 15334 413 15364 497
rect 15433 413 15463 497
rect 15573 413 15603 497
rect 15670 413 15700 497
rect 15867 329 15897 497
rect 15966 413 15996 497
rect 16052 413 16082 497
rect 16136 413 16166 497
rect 16244 413 16274 497
rect 16328 413 16358 497
rect 16492 297 16522 497
rect 16711 369 16741 497
rect 16808 297 16838 497
rect 17007 363 17037 491
rect 17091 363 17121 491
rect 17358 413 17388 497
rect 17450 413 17480 497
rect 17549 413 17579 497
rect 17689 413 17719 497
rect 17786 413 17816 497
rect 17983 329 18013 497
rect 18082 413 18112 497
rect 18168 413 18198 497
rect 18252 413 18282 497
rect 18360 413 18390 497
rect 18444 413 18474 497
rect 18608 297 18638 497
rect 18827 369 18857 497
rect 18924 297 18954 497
rect 19123 363 19153 491
rect 19207 363 19237 491
rect 19474 413 19504 497
rect 19566 413 19596 497
rect 19665 413 19695 497
rect 19805 413 19835 497
rect 19902 413 19932 497
rect 20099 329 20129 497
rect 20198 413 20228 497
rect 20284 413 20314 497
rect 20368 413 20398 497
rect 20476 413 20506 497
rect 20560 413 20590 497
rect 20724 297 20754 497
rect 20943 369 20973 497
rect 21040 297 21070 497
rect 21239 363 21269 491
rect 21323 363 21353 491
rect 21590 413 21620 497
rect 21682 413 21712 497
rect 21781 413 21811 497
rect 21921 413 21951 497
rect 22018 413 22048 497
rect 22215 329 22245 497
rect 22314 413 22344 497
rect 22400 413 22430 497
rect 22484 413 22514 497
rect 22592 413 22622 497
rect 22676 413 22706 497
rect 22840 297 22870 497
rect 23059 369 23089 497
rect 23156 297 23186 497
rect 23355 363 23385 491
rect 23439 363 23469 491
rect 23706 413 23736 497
rect 23798 413 23828 497
rect 23897 413 23927 497
rect 24037 413 24067 497
rect 24134 413 24164 497
rect 24331 329 24361 497
rect 24430 413 24460 497
rect 24516 413 24546 497
rect 24600 413 24630 497
rect 24708 413 24738 497
rect 24792 413 24822 497
rect 24956 297 24986 497
rect 25175 369 25205 497
rect 25272 297 25302 497
rect 25471 363 25501 491
rect 25555 363 25585 491
rect 25822 413 25852 497
rect 25914 413 25944 497
rect 26013 413 26043 497
rect 26153 413 26183 497
rect 26250 413 26280 497
rect 26447 329 26477 497
rect 26546 413 26576 497
rect 26632 413 26662 497
rect 26716 413 26746 497
rect 26824 413 26854 497
rect 26908 413 26938 497
rect 27072 297 27102 497
rect 27291 369 27321 497
rect 27388 297 27418 497
rect 27587 363 27617 491
rect 27671 363 27701 491
rect 27938 413 27968 497
rect 28030 413 28060 497
rect 28129 413 28159 497
rect 28269 413 28299 497
rect 28366 413 28396 497
rect 28563 329 28593 497
rect 28662 413 28692 497
rect 28748 413 28778 497
rect 28832 413 28862 497
rect 28940 413 28970 497
rect 29024 413 29054 497
rect 29188 297 29218 497
rect 29407 369 29437 497
rect 29504 297 29534 497
rect 29703 363 29733 491
rect 29787 363 29817 491
rect 30054 413 30084 497
rect 30146 413 30176 497
rect 30245 413 30275 497
rect 30385 413 30415 497
rect 30482 413 30512 497
rect 30679 329 30709 497
rect 30778 413 30808 497
rect 30864 413 30894 497
rect 30948 413 30978 497
rect 31056 413 31086 497
rect 31140 413 31170 497
rect 31304 297 31334 497
rect 31523 369 31553 497
rect 31620 297 31650 497
rect 31819 363 31849 491
rect 31903 363 31933 491
rect 32170 413 32200 497
rect 32262 413 32292 497
rect 32361 413 32391 497
rect 32501 413 32531 497
rect 32598 413 32628 497
rect 32795 329 32825 497
rect 32894 413 32924 497
rect 32980 413 33010 497
rect 33064 413 33094 497
rect 33172 413 33202 497
rect 33256 413 33286 497
rect 33420 297 33450 497
rect 33639 369 33669 497
rect 33736 297 33766 497
rect 33935 363 33965 491
rect 34019 363 34049 491
rect 34286 413 34316 497
rect 34378 413 34408 497
rect 34477 413 34507 497
rect 34617 413 34647 497
rect 34714 413 34744 497
rect 34911 329 34941 497
rect 35010 413 35040 497
rect 35096 413 35126 497
rect 35180 413 35210 497
rect 35288 413 35318 497
rect 35372 413 35402 497
rect 35536 297 35566 497
rect 35755 369 35785 497
rect 35852 297 35882 497
rect 36051 363 36081 491
rect 36135 363 36165 491
rect 36402 413 36432 497
rect 36494 413 36524 497
rect 36593 413 36623 497
rect 36733 413 36763 497
rect 36830 413 36860 497
rect 37027 329 37057 497
rect 37126 413 37156 497
rect 37212 413 37242 497
rect 37296 413 37326 497
rect 37404 413 37434 497
rect 37488 413 37518 497
rect 37652 297 37682 497
rect 37871 369 37901 497
rect 37968 297 37998 497
rect 38167 363 38197 491
rect 38251 363 38281 491
rect 38518 413 38548 497
rect 38610 413 38640 497
rect 38709 413 38739 497
rect 38849 413 38879 497
rect 38946 413 38976 497
rect 39143 329 39173 497
rect 39242 413 39272 497
rect 39328 413 39358 497
rect 39412 413 39442 497
rect 39520 413 39550 497
rect 39604 413 39634 497
rect 39768 297 39798 497
rect 39987 369 40017 497
rect 40084 297 40114 497
rect 40283 363 40313 491
rect 40367 363 40397 491
rect 40634 413 40664 497
rect 40726 413 40756 497
rect 40825 413 40855 497
rect 40965 413 40995 497
rect 41062 413 41092 497
rect 41259 329 41289 497
rect 41358 413 41388 497
rect 41444 413 41474 497
rect 41528 413 41558 497
rect 41636 413 41666 497
rect 41720 413 41750 497
rect 41884 297 41914 497
rect 42103 369 42133 497
rect 42200 297 42230 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 313 89 418 131
rect 313 55 325 89
rect 359 55 418 89
rect 313 47 418 55
rect 448 119 498 131
rect 929 131 979 175
rect 657 119 775 131
rect 448 95 513 119
rect 448 61 458 95
rect 492 61 513 95
rect 448 47 513 61
rect 543 95 609 119
rect 543 61 565 95
rect 599 61 609 95
rect 543 47 609 61
rect 639 47 775 119
rect 805 47 847 131
rect 877 93 979 131
rect 877 59 911 93
rect 945 59 979 93
rect 877 47 979 59
rect 1009 119 1063 175
rect 1659 132 1711 177
rect 1233 119 1283 131
rect 1009 89 1078 119
rect 1009 55 1023 89
rect 1057 55 1078 89
rect 1009 47 1078 55
rect 1108 93 1187 119
rect 1108 59 1133 93
rect 1167 59 1187 93
rect 1108 47 1187 59
rect 1217 47 1283 119
rect 1313 89 1432 131
rect 1313 55 1345 89
rect 1379 55 1432 89
rect 1313 47 1432 55
rect 1462 47 1523 131
rect 1553 109 1605 131
rect 1553 75 1563 109
rect 1597 75 1605 109
rect 1553 47 1605 75
rect 1659 98 1667 132
rect 1701 98 1711 132
rect 1659 47 1711 98
rect 1741 165 1793 177
rect 1741 131 1751 165
rect 1785 131 1793 165
rect 1944 131 1996 177
rect 1741 97 1793 131
rect 1741 63 1751 97
rect 1785 63 1793 97
rect 1741 47 1793 63
rect 1847 119 1899 131
rect 1847 85 1855 119
rect 1889 85 1899 119
rect 1847 47 1899 85
rect 1929 113 1996 131
rect 1929 79 1952 113
rect 1986 79 1996 113
rect 1929 47 1996 79
rect 2026 143 2078 177
rect 2026 109 2036 143
rect 2070 109 2078 143
rect 2026 47 2078 109
rect 2143 119 2195 131
rect 2143 85 2151 119
rect 2185 85 2195 119
rect 2143 47 2195 85
rect 2225 93 2279 131
rect 2225 59 2235 93
rect 2269 59 2279 93
rect 2225 47 2279 59
rect 2309 119 2361 131
rect 2309 85 2319 119
rect 2353 85 2361 119
rect 2309 47 2361 85
rect 2429 89 2534 131
rect 2429 55 2441 89
rect 2475 55 2534 89
rect 2429 47 2534 55
rect 2564 119 2614 131
rect 3045 131 3095 175
rect 2773 119 2891 131
rect 2564 95 2629 119
rect 2564 61 2574 95
rect 2608 61 2629 95
rect 2564 47 2629 61
rect 2659 95 2725 119
rect 2659 61 2681 95
rect 2715 61 2725 95
rect 2659 47 2725 61
rect 2755 47 2891 119
rect 2921 47 2963 131
rect 2993 93 3095 131
rect 2993 59 3027 93
rect 3061 59 3095 93
rect 2993 47 3095 59
rect 3125 119 3179 175
rect 3775 132 3827 177
rect 3349 119 3399 131
rect 3125 89 3194 119
rect 3125 55 3139 89
rect 3173 55 3194 89
rect 3125 47 3194 55
rect 3224 93 3303 119
rect 3224 59 3249 93
rect 3283 59 3303 93
rect 3224 47 3303 59
rect 3333 47 3399 119
rect 3429 89 3548 131
rect 3429 55 3461 89
rect 3495 55 3548 89
rect 3429 47 3548 55
rect 3578 47 3639 131
rect 3669 109 3721 131
rect 3669 75 3679 109
rect 3713 75 3721 109
rect 3669 47 3721 75
rect 3775 98 3783 132
rect 3817 98 3827 132
rect 3775 47 3827 98
rect 3857 165 3909 177
rect 3857 131 3867 165
rect 3901 131 3909 165
rect 4060 131 4112 177
rect 3857 97 3909 131
rect 3857 63 3867 97
rect 3901 63 3909 97
rect 3857 47 3909 63
rect 3963 119 4015 131
rect 3963 85 3971 119
rect 4005 85 4015 119
rect 3963 47 4015 85
rect 4045 113 4112 131
rect 4045 79 4068 113
rect 4102 79 4112 113
rect 4045 47 4112 79
rect 4142 143 4194 177
rect 4142 109 4152 143
rect 4186 109 4194 143
rect 4142 47 4194 109
rect 4259 119 4311 131
rect 4259 85 4267 119
rect 4301 85 4311 119
rect 4259 47 4311 85
rect 4341 93 4395 131
rect 4341 59 4351 93
rect 4385 59 4395 93
rect 4341 47 4395 59
rect 4425 119 4477 131
rect 4425 85 4435 119
rect 4469 85 4477 119
rect 4425 47 4477 85
rect 4545 89 4650 131
rect 4545 55 4557 89
rect 4591 55 4650 89
rect 4545 47 4650 55
rect 4680 119 4730 131
rect 5161 131 5211 175
rect 4889 119 5007 131
rect 4680 95 4745 119
rect 4680 61 4690 95
rect 4724 61 4745 95
rect 4680 47 4745 61
rect 4775 95 4841 119
rect 4775 61 4797 95
rect 4831 61 4841 95
rect 4775 47 4841 61
rect 4871 47 5007 119
rect 5037 47 5079 131
rect 5109 93 5211 131
rect 5109 59 5143 93
rect 5177 59 5211 93
rect 5109 47 5211 59
rect 5241 119 5295 175
rect 5891 132 5943 177
rect 5465 119 5515 131
rect 5241 89 5310 119
rect 5241 55 5255 89
rect 5289 55 5310 89
rect 5241 47 5310 55
rect 5340 93 5419 119
rect 5340 59 5365 93
rect 5399 59 5419 93
rect 5340 47 5419 59
rect 5449 47 5515 119
rect 5545 89 5664 131
rect 5545 55 5577 89
rect 5611 55 5664 89
rect 5545 47 5664 55
rect 5694 47 5755 131
rect 5785 109 5837 131
rect 5785 75 5795 109
rect 5829 75 5837 109
rect 5785 47 5837 75
rect 5891 98 5899 132
rect 5933 98 5943 132
rect 5891 47 5943 98
rect 5973 165 6025 177
rect 5973 131 5983 165
rect 6017 131 6025 165
rect 6176 131 6228 177
rect 5973 97 6025 131
rect 5973 63 5983 97
rect 6017 63 6025 97
rect 5973 47 6025 63
rect 6079 119 6131 131
rect 6079 85 6087 119
rect 6121 85 6131 119
rect 6079 47 6131 85
rect 6161 113 6228 131
rect 6161 79 6184 113
rect 6218 79 6228 113
rect 6161 47 6228 79
rect 6258 143 6310 177
rect 6258 109 6268 143
rect 6302 109 6310 143
rect 6258 47 6310 109
rect 6375 119 6427 131
rect 6375 85 6383 119
rect 6417 85 6427 119
rect 6375 47 6427 85
rect 6457 93 6511 131
rect 6457 59 6467 93
rect 6501 59 6511 93
rect 6457 47 6511 59
rect 6541 119 6593 131
rect 6541 85 6551 119
rect 6585 85 6593 119
rect 6541 47 6593 85
rect 6661 89 6766 131
rect 6661 55 6673 89
rect 6707 55 6766 89
rect 6661 47 6766 55
rect 6796 119 6846 131
rect 7277 131 7327 175
rect 7005 119 7123 131
rect 6796 95 6861 119
rect 6796 61 6806 95
rect 6840 61 6861 95
rect 6796 47 6861 61
rect 6891 95 6957 119
rect 6891 61 6913 95
rect 6947 61 6957 95
rect 6891 47 6957 61
rect 6987 47 7123 119
rect 7153 47 7195 131
rect 7225 93 7327 131
rect 7225 59 7259 93
rect 7293 59 7327 93
rect 7225 47 7327 59
rect 7357 119 7411 175
rect 8007 132 8059 177
rect 7581 119 7631 131
rect 7357 89 7426 119
rect 7357 55 7371 89
rect 7405 55 7426 89
rect 7357 47 7426 55
rect 7456 93 7535 119
rect 7456 59 7481 93
rect 7515 59 7535 93
rect 7456 47 7535 59
rect 7565 47 7631 119
rect 7661 89 7780 131
rect 7661 55 7693 89
rect 7727 55 7780 89
rect 7661 47 7780 55
rect 7810 47 7871 131
rect 7901 109 7953 131
rect 7901 75 7911 109
rect 7945 75 7953 109
rect 7901 47 7953 75
rect 8007 98 8015 132
rect 8049 98 8059 132
rect 8007 47 8059 98
rect 8089 165 8141 177
rect 8089 131 8099 165
rect 8133 131 8141 165
rect 8292 131 8344 177
rect 8089 97 8141 131
rect 8089 63 8099 97
rect 8133 63 8141 97
rect 8089 47 8141 63
rect 8195 119 8247 131
rect 8195 85 8203 119
rect 8237 85 8247 119
rect 8195 47 8247 85
rect 8277 113 8344 131
rect 8277 79 8300 113
rect 8334 79 8344 113
rect 8277 47 8344 79
rect 8374 143 8426 177
rect 8374 109 8384 143
rect 8418 109 8426 143
rect 8374 47 8426 109
rect 8491 119 8543 131
rect 8491 85 8499 119
rect 8533 85 8543 119
rect 8491 47 8543 85
rect 8573 93 8627 131
rect 8573 59 8583 93
rect 8617 59 8627 93
rect 8573 47 8627 59
rect 8657 119 8709 131
rect 8657 85 8667 119
rect 8701 85 8709 119
rect 8657 47 8709 85
rect 8777 89 8882 131
rect 8777 55 8789 89
rect 8823 55 8882 89
rect 8777 47 8882 55
rect 8912 119 8962 131
rect 9393 131 9443 175
rect 9121 119 9239 131
rect 8912 95 8977 119
rect 8912 61 8922 95
rect 8956 61 8977 95
rect 8912 47 8977 61
rect 9007 95 9073 119
rect 9007 61 9029 95
rect 9063 61 9073 95
rect 9007 47 9073 61
rect 9103 47 9239 119
rect 9269 47 9311 131
rect 9341 93 9443 131
rect 9341 59 9375 93
rect 9409 59 9443 93
rect 9341 47 9443 59
rect 9473 119 9527 175
rect 10123 132 10175 177
rect 9697 119 9747 131
rect 9473 89 9542 119
rect 9473 55 9487 89
rect 9521 55 9542 89
rect 9473 47 9542 55
rect 9572 93 9651 119
rect 9572 59 9597 93
rect 9631 59 9651 93
rect 9572 47 9651 59
rect 9681 47 9747 119
rect 9777 89 9896 131
rect 9777 55 9809 89
rect 9843 55 9896 89
rect 9777 47 9896 55
rect 9926 47 9987 131
rect 10017 109 10069 131
rect 10017 75 10027 109
rect 10061 75 10069 109
rect 10017 47 10069 75
rect 10123 98 10131 132
rect 10165 98 10175 132
rect 10123 47 10175 98
rect 10205 165 10257 177
rect 10205 131 10215 165
rect 10249 131 10257 165
rect 10408 131 10460 177
rect 10205 97 10257 131
rect 10205 63 10215 97
rect 10249 63 10257 97
rect 10205 47 10257 63
rect 10311 119 10363 131
rect 10311 85 10319 119
rect 10353 85 10363 119
rect 10311 47 10363 85
rect 10393 113 10460 131
rect 10393 79 10416 113
rect 10450 79 10460 113
rect 10393 47 10460 79
rect 10490 143 10542 177
rect 10490 109 10500 143
rect 10534 109 10542 143
rect 10490 47 10542 109
rect 10607 119 10659 131
rect 10607 85 10615 119
rect 10649 85 10659 119
rect 10607 47 10659 85
rect 10689 93 10743 131
rect 10689 59 10699 93
rect 10733 59 10743 93
rect 10689 47 10743 59
rect 10773 119 10825 131
rect 10773 85 10783 119
rect 10817 85 10825 119
rect 10773 47 10825 85
rect 10893 89 10998 131
rect 10893 55 10905 89
rect 10939 55 10998 89
rect 10893 47 10998 55
rect 11028 119 11078 131
rect 11509 131 11559 175
rect 11237 119 11355 131
rect 11028 95 11093 119
rect 11028 61 11038 95
rect 11072 61 11093 95
rect 11028 47 11093 61
rect 11123 95 11189 119
rect 11123 61 11145 95
rect 11179 61 11189 95
rect 11123 47 11189 61
rect 11219 47 11355 119
rect 11385 47 11427 131
rect 11457 93 11559 131
rect 11457 59 11491 93
rect 11525 59 11559 93
rect 11457 47 11559 59
rect 11589 119 11643 175
rect 12239 132 12291 177
rect 11813 119 11863 131
rect 11589 89 11658 119
rect 11589 55 11603 89
rect 11637 55 11658 89
rect 11589 47 11658 55
rect 11688 93 11767 119
rect 11688 59 11713 93
rect 11747 59 11767 93
rect 11688 47 11767 59
rect 11797 47 11863 119
rect 11893 89 12012 131
rect 11893 55 11925 89
rect 11959 55 12012 89
rect 11893 47 12012 55
rect 12042 47 12103 131
rect 12133 109 12185 131
rect 12133 75 12143 109
rect 12177 75 12185 109
rect 12133 47 12185 75
rect 12239 98 12247 132
rect 12281 98 12291 132
rect 12239 47 12291 98
rect 12321 165 12373 177
rect 12321 131 12331 165
rect 12365 131 12373 165
rect 12524 131 12576 177
rect 12321 97 12373 131
rect 12321 63 12331 97
rect 12365 63 12373 97
rect 12321 47 12373 63
rect 12427 119 12479 131
rect 12427 85 12435 119
rect 12469 85 12479 119
rect 12427 47 12479 85
rect 12509 113 12576 131
rect 12509 79 12532 113
rect 12566 79 12576 113
rect 12509 47 12576 79
rect 12606 143 12658 177
rect 12606 109 12616 143
rect 12650 109 12658 143
rect 12606 47 12658 109
rect 12723 119 12775 131
rect 12723 85 12731 119
rect 12765 85 12775 119
rect 12723 47 12775 85
rect 12805 93 12859 131
rect 12805 59 12815 93
rect 12849 59 12859 93
rect 12805 47 12859 59
rect 12889 119 12941 131
rect 12889 85 12899 119
rect 12933 85 12941 119
rect 12889 47 12941 85
rect 13009 89 13114 131
rect 13009 55 13021 89
rect 13055 55 13114 89
rect 13009 47 13114 55
rect 13144 119 13194 131
rect 13625 131 13675 175
rect 13353 119 13471 131
rect 13144 95 13209 119
rect 13144 61 13154 95
rect 13188 61 13209 95
rect 13144 47 13209 61
rect 13239 95 13305 119
rect 13239 61 13261 95
rect 13295 61 13305 95
rect 13239 47 13305 61
rect 13335 47 13471 119
rect 13501 47 13543 131
rect 13573 93 13675 131
rect 13573 59 13607 93
rect 13641 59 13675 93
rect 13573 47 13675 59
rect 13705 119 13759 175
rect 14355 132 14407 177
rect 13929 119 13979 131
rect 13705 89 13774 119
rect 13705 55 13719 89
rect 13753 55 13774 89
rect 13705 47 13774 55
rect 13804 93 13883 119
rect 13804 59 13829 93
rect 13863 59 13883 93
rect 13804 47 13883 59
rect 13913 47 13979 119
rect 14009 89 14128 131
rect 14009 55 14041 89
rect 14075 55 14128 89
rect 14009 47 14128 55
rect 14158 47 14219 131
rect 14249 109 14301 131
rect 14249 75 14259 109
rect 14293 75 14301 109
rect 14249 47 14301 75
rect 14355 98 14363 132
rect 14397 98 14407 132
rect 14355 47 14407 98
rect 14437 165 14489 177
rect 14437 131 14447 165
rect 14481 131 14489 165
rect 14640 131 14692 177
rect 14437 97 14489 131
rect 14437 63 14447 97
rect 14481 63 14489 97
rect 14437 47 14489 63
rect 14543 119 14595 131
rect 14543 85 14551 119
rect 14585 85 14595 119
rect 14543 47 14595 85
rect 14625 113 14692 131
rect 14625 79 14648 113
rect 14682 79 14692 113
rect 14625 47 14692 79
rect 14722 143 14774 177
rect 14722 109 14732 143
rect 14766 109 14774 143
rect 14722 47 14774 109
rect 14839 119 14891 131
rect 14839 85 14847 119
rect 14881 85 14891 119
rect 14839 47 14891 85
rect 14921 93 14975 131
rect 14921 59 14931 93
rect 14965 59 14975 93
rect 14921 47 14975 59
rect 15005 119 15057 131
rect 15005 85 15015 119
rect 15049 85 15057 119
rect 15005 47 15057 85
rect 15125 89 15230 131
rect 15125 55 15137 89
rect 15171 55 15230 89
rect 15125 47 15230 55
rect 15260 119 15310 131
rect 15741 131 15791 175
rect 15469 119 15587 131
rect 15260 95 15325 119
rect 15260 61 15270 95
rect 15304 61 15325 95
rect 15260 47 15325 61
rect 15355 95 15421 119
rect 15355 61 15377 95
rect 15411 61 15421 95
rect 15355 47 15421 61
rect 15451 47 15587 119
rect 15617 47 15659 131
rect 15689 93 15791 131
rect 15689 59 15723 93
rect 15757 59 15791 93
rect 15689 47 15791 59
rect 15821 119 15875 175
rect 16471 132 16523 177
rect 16045 119 16095 131
rect 15821 89 15890 119
rect 15821 55 15835 89
rect 15869 55 15890 89
rect 15821 47 15890 55
rect 15920 93 15999 119
rect 15920 59 15945 93
rect 15979 59 15999 93
rect 15920 47 15999 59
rect 16029 47 16095 119
rect 16125 89 16244 131
rect 16125 55 16157 89
rect 16191 55 16244 89
rect 16125 47 16244 55
rect 16274 47 16335 131
rect 16365 109 16417 131
rect 16365 75 16375 109
rect 16409 75 16417 109
rect 16365 47 16417 75
rect 16471 98 16479 132
rect 16513 98 16523 132
rect 16471 47 16523 98
rect 16553 165 16605 177
rect 16553 131 16563 165
rect 16597 131 16605 165
rect 16756 131 16808 177
rect 16553 97 16605 131
rect 16553 63 16563 97
rect 16597 63 16605 97
rect 16553 47 16605 63
rect 16659 119 16711 131
rect 16659 85 16667 119
rect 16701 85 16711 119
rect 16659 47 16711 85
rect 16741 113 16808 131
rect 16741 79 16764 113
rect 16798 79 16808 113
rect 16741 47 16808 79
rect 16838 143 16890 177
rect 16838 109 16848 143
rect 16882 109 16890 143
rect 16838 47 16890 109
rect 16955 119 17007 131
rect 16955 85 16963 119
rect 16997 85 17007 119
rect 16955 47 17007 85
rect 17037 93 17091 131
rect 17037 59 17047 93
rect 17081 59 17091 93
rect 17037 47 17091 59
rect 17121 119 17173 131
rect 17121 85 17131 119
rect 17165 85 17173 119
rect 17121 47 17173 85
rect 17241 89 17346 131
rect 17241 55 17253 89
rect 17287 55 17346 89
rect 17241 47 17346 55
rect 17376 119 17426 131
rect 17857 131 17907 175
rect 17585 119 17703 131
rect 17376 95 17441 119
rect 17376 61 17386 95
rect 17420 61 17441 95
rect 17376 47 17441 61
rect 17471 95 17537 119
rect 17471 61 17493 95
rect 17527 61 17537 95
rect 17471 47 17537 61
rect 17567 47 17703 119
rect 17733 47 17775 131
rect 17805 93 17907 131
rect 17805 59 17839 93
rect 17873 59 17907 93
rect 17805 47 17907 59
rect 17937 119 17991 175
rect 18587 132 18639 177
rect 18161 119 18211 131
rect 17937 89 18006 119
rect 17937 55 17951 89
rect 17985 55 18006 89
rect 17937 47 18006 55
rect 18036 93 18115 119
rect 18036 59 18061 93
rect 18095 59 18115 93
rect 18036 47 18115 59
rect 18145 47 18211 119
rect 18241 89 18360 131
rect 18241 55 18273 89
rect 18307 55 18360 89
rect 18241 47 18360 55
rect 18390 47 18451 131
rect 18481 109 18533 131
rect 18481 75 18491 109
rect 18525 75 18533 109
rect 18481 47 18533 75
rect 18587 98 18595 132
rect 18629 98 18639 132
rect 18587 47 18639 98
rect 18669 165 18721 177
rect 18669 131 18679 165
rect 18713 131 18721 165
rect 18872 131 18924 177
rect 18669 97 18721 131
rect 18669 63 18679 97
rect 18713 63 18721 97
rect 18669 47 18721 63
rect 18775 119 18827 131
rect 18775 85 18783 119
rect 18817 85 18827 119
rect 18775 47 18827 85
rect 18857 113 18924 131
rect 18857 79 18880 113
rect 18914 79 18924 113
rect 18857 47 18924 79
rect 18954 143 19006 177
rect 18954 109 18964 143
rect 18998 109 19006 143
rect 18954 47 19006 109
rect 19071 119 19123 131
rect 19071 85 19079 119
rect 19113 85 19123 119
rect 19071 47 19123 85
rect 19153 93 19207 131
rect 19153 59 19163 93
rect 19197 59 19207 93
rect 19153 47 19207 59
rect 19237 119 19289 131
rect 19237 85 19247 119
rect 19281 85 19289 119
rect 19237 47 19289 85
rect 19357 89 19462 131
rect 19357 55 19369 89
rect 19403 55 19462 89
rect 19357 47 19462 55
rect 19492 119 19542 131
rect 19973 131 20023 175
rect 19701 119 19819 131
rect 19492 95 19557 119
rect 19492 61 19502 95
rect 19536 61 19557 95
rect 19492 47 19557 61
rect 19587 95 19653 119
rect 19587 61 19609 95
rect 19643 61 19653 95
rect 19587 47 19653 61
rect 19683 47 19819 119
rect 19849 47 19891 131
rect 19921 93 20023 131
rect 19921 59 19955 93
rect 19989 59 20023 93
rect 19921 47 20023 59
rect 20053 119 20107 175
rect 20703 132 20755 177
rect 20277 119 20327 131
rect 20053 89 20122 119
rect 20053 55 20067 89
rect 20101 55 20122 89
rect 20053 47 20122 55
rect 20152 93 20231 119
rect 20152 59 20177 93
rect 20211 59 20231 93
rect 20152 47 20231 59
rect 20261 47 20327 119
rect 20357 89 20476 131
rect 20357 55 20389 89
rect 20423 55 20476 89
rect 20357 47 20476 55
rect 20506 47 20567 131
rect 20597 109 20649 131
rect 20597 75 20607 109
rect 20641 75 20649 109
rect 20597 47 20649 75
rect 20703 98 20711 132
rect 20745 98 20755 132
rect 20703 47 20755 98
rect 20785 165 20837 177
rect 20785 131 20795 165
rect 20829 131 20837 165
rect 20988 131 21040 177
rect 20785 97 20837 131
rect 20785 63 20795 97
rect 20829 63 20837 97
rect 20785 47 20837 63
rect 20891 119 20943 131
rect 20891 85 20899 119
rect 20933 85 20943 119
rect 20891 47 20943 85
rect 20973 113 21040 131
rect 20973 79 20996 113
rect 21030 79 21040 113
rect 20973 47 21040 79
rect 21070 143 21122 177
rect 21070 109 21080 143
rect 21114 109 21122 143
rect 21070 47 21122 109
rect 21187 119 21239 131
rect 21187 85 21195 119
rect 21229 85 21239 119
rect 21187 47 21239 85
rect 21269 93 21323 131
rect 21269 59 21279 93
rect 21313 59 21323 93
rect 21269 47 21323 59
rect 21353 119 21405 131
rect 21353 85 21363 119
rect 21397 85 21405 119
rect 21353 47 21405 85
rect 21473 89 21578 131
rect 21473 55 21485 89
rect 21519 55 21578 89
rect 21473 47 21578 55
rect 21608 119 21658 131
rect 22089 131 22139 175
rect 21817 119 21935 131
rect 21608 95 21673 119
rect 21608 61 21618 95
rect 21652 61 21673 95
rect 21608 47 21673 61
rect 21703 95 21769 119
rect 21703 61 21725 95
rect 21759 61 21769 95
rect 21703 47 21769 61
rect 21799 47 21935 119
rect 21965 47 22007 131
rect 22037 93 22139 131
rect 22037 59 22071 93
rect 22105 59 22139 93
rect 22037 47 22139 59
rect 22169 119 22223 175
rect 22819 132 22871 177
rect 22393 119 22443 131
rect 22169 89 22238 119
rect 22169 55 22183 89
rect 22217 55 22238 89
rect 22169 47 22238 55
rect 22268 93 22347 119
rect 22268 59 22293 93
rect 22327 59 22347 93
rect 22268 47 22347 59
rect 22377 47 22443 119
rect 22473 89 22592 131
rect 22473 55 22505 89
rect 22539 55 22592 89
rect 22473 47 22592 55
rect 22622 47 22683 131
rect 22713 109 22765 131
rect 22713 75 22723 109
rect 22757 75 22765 109
rect 22713 47 22765 75
rect 22819 98 22827 132
rect 22861 98 22871 132
rect 22819 47 22871 98
rect 22901 165 22953 177
rect 22901 131 22911 165
rect 22945 131 22953 165
rect 23104 131 23156 177
rect 22901 97 22953 131
rect 22901 63 22911 97
rect 22945 63 22953 97
rect 22901 47 22953 63
rect 23007 119 23059 131
rect 23007 85 23015 119
rect 23049 85 23059 119
rect 23007 47 23059 85
rect 23089 113 23156 131
rect 23089 79 23112 113
rect 23146 79 23156 113
rect 23089 47 23156 79
rect 23186 143 23238 177
rect 23186 109 23196 143
rect 23230 109 23238 143
rect 23186 47 23238 109
rect 23303 119 23355 131
rect 23303 85 23311 119
rect 23345 85 23355 119
rect 23303 47 23355 85
rect 23385 93 23439 131
rect 23385 59 23395 93
rect 23429 59 23439 93
rect 23385 47 23439 59
rect 23469 119 23521 131
rect 23469 85 23479 119
rect 23513 85 23521 119
rect 23469 47 23521 85
rect 23589 89 23694 131
rect 23589 55 23601 89
rect 23635 55 23694 89
rect 23589 47 23694 55
rect 23724 119 23774 131
rect 24205 131 24255 175
rect 23933 119 24051 131
rect 23724 95 23789 119
rect 23724 61 23734 95
rect 23768 61 23789 95
rect 23724 47 23789 61
rect 23819 95 23885 119
rect 23819 61 23841 95
rect 23875 61 23885 95
rect 23819 47 23885 61
rect 23915 47 24051 119
rect 24081 47 24123 131
rect 24153 93 24255 131
rect 24153 59 24187 93
rect 24221 59 24255 93
rect 24153 47 24255 59
rect 24285 119 24339 175
rect 24935 132 24987 177
rect 24509 119 24559 131
rect 24285 89 24354 119
rect 24285 55 24299 89
rect 24333 55 24354 89
rect 24285 47 24354 55
rect 24384 93 24463 119
rect 24384 59 24409 93
rect 24443 59 24463 93
rect 24384 47 24463 59
rect 24493 47 24559 119
rect 24589 89 24708 131
rect 24589 55 24621 89
rect 24655 55 24708 89
rect 24589 47 24708 55
rect 24738 47 24799 131
rect 24829 109 24881 131
rect 24829 75 24839 109
rect 24873 75 24881 109
rect 24829 47 24881 75
rect 24935 98 24943 132
rect 24977 98 24987 132
rect 24935 47 24987 98
rect 25017 165 25069 177
rect 25017 131 25027 165
rect 25061 131 25069 165
rect 25220 131 25272 177
rect 25017 97 25069 131
rect 25017 63 25027 97
rect 25061 63 25069 97
rect 25017 47 25069 63
rect 25123 119 25175 131
rect 25123 85 25131 119
rect 25165 85 25175 119
rect 25123 47 25175 85
rect 25205 113 25272 131
rect 25205 79 25228 113
rect 25262 79 25272 113
rect 25205 47 25272 79
rect 25302 143 25354 177
rect 25302 109 25312 143
rect 25346 109 25354 143
rect 25302 47 25354 109
rect 25419 119 25471 131
rect 25419 85 25427 119
rect 25461 85 25471 119
rect 25419 47 25471 85
rect 25501 93 25555 131
rect 25501 59 25511 93
rect 25545 59 25555 93
rect 25501 47 25555 59
rect 25585 119 25637 131
rect 25585 85 25595 119
rect 25629 85 25637 119
rect 25585 47 25637 85
rect 25705 89 25810 131
rect 25705 55 25717 89
rect 25751 55 25810 89
rect 25705 47 25810 55
rect 25840 119 25890 131
rect 26321 131 26371 175
rect 26049 119 26167 131
rect 25840 95 25905 119
rect 25840 61 25850 95
rect 25884 61 25905 95
rect 25840 47 25905 61
rect 25935 95 26001 119
rect 25935 61 25957 95
rect 25991 61 26001 95
rect 25935 47 26001 61
rect 26031 47 26167 119
rect 26197 47 26239 131
rect 26269 93 26371 131
rect 26269 59 26303 93
rect 26337 59 26371 93
rect 26269 47 26371 59
rect 26401 119 26455 175
rect 27051 132 27103 177
rect 26625 119 26675 131
rect 26401 89 26470 119
rect 26401 55 26415 89
rect 26449 55 26470 89
rect 26401 47 26470 55
rect 26500 93 26579 119
rect 26500 59 26525 93
rect 26559 59 26579 93
rect 26500 47 26579 59
rect 26609 47 26675 119
rect 26705 89 26824 131
rect 26705 55 26737 89
rect 26771 55 26824 89
rect 26705 47 26824 55
rect 26854 47 26915 131
rect 26945 109 26997 131
rect 26945 75 26955 109
rect 26989 75 26997 109
rect 26945 47 26997 75
rect 27051 98 27059 132
rect 27093 98 27103 132
rect 27051 47 27103 98
rect 27133 165 27185 177
rect 27133 131 27143 165
rect 27177 131 27185 165
rect 27336 131 27388 177
rect 27133 97 27185 131
rect 27133 63 27143 97
rect 27177 63 27185 97
rect 27133 47 27185 63
rect 27239 119 27291 131
rect 27239 85 27247 119
rect 27281 85 27291 119
rect 27239 47 27291 85
rect 27321 113 27388 131
rect 27321 79 27344 113
rect 27378 79 27388 113
rect 27321 47 27388 79
rect 27418 143 27470 177
rect 27418 109 27428 143
rect 27462 109 27470 143
rect 27418 47 27470 109
rect 27535 119 27587 131
rect 27535 85 27543 119
rect 27577 85 27587 119
rect 27535 47 27587 85
rect 27617 93 27671 131
rect 27617 59 27627 93
rect 27661 59 27671 93
rect 27617 47 27671 59
rect 27701 119 27753 131
rect 27701 85 27711 119
rect 27745 85 27753 119
rect 27701 47 27753 85
rect 27821 89 27926 131
rect 27821 55 27833 89
rect 27867 55 27926 89
rect 27821 47 27926 55
rect 27956 119 28006 131
rect 28437 131 28487 175
rect 28165 119 28283 131
rect 27956 95 28021 119
rect 27956 61 27966 95
rect 28000 61 28021 95
rect 27956 47 28021 61
rect 28051 95 28117 119
rect 28051 61 28073 95
rect 28107 61 28117 95
rect 28051 47 28117 61
rect 28147 47 28283 119
rect 28313 47 28355 131
rect 28385 93 28487 131
rect 28385 59 28419 93
rect 28453 59 28487 93
rect 28385 47 28487 59
rect 28517 119 28571 175
rect 29167 132 29219 177
rect 28741 119 28791 131
rect 28517 89 28586 119
rect 28517 55 28531 89
rect 28565 55 28586 89
rect 28517 47 28586 55
rect 28616 93 28695 119
rect 28616 59 28641 93
rect 28675 59 28695 93
rect 28616 47 28695 59
rect 28725 47 28791 119
rect 28821 89 28940 131
rect 28821 55 28853 89
rect 28887 55 28940 89
rect 28821 47 28940 55
rect 28970 47 29031 131
rect 29061 109 29113 131
rect 29061 75 29071 109
rect 29105 75 29113 109
rect 29061 47 29113 75
rect 29167 98 29175 132
rect 29209 98 29219 132
rect 29167 47 29219 98
rect 29249 165 29301 177
rect 29249 131 29259 165
rect 29293 131 29301 165
rect 29452 131 29504 177
rect 29249 97 29301 131
rect 29249 63 29259 97
rect 29293 63 29301 97
rect 29249 47 29301 63
rect 29355 119 29407 131
rect 29355 85 29363 119
rect 29397 85 29407 119
rect 29355 47 29407 85
rect 29437 113 29504 131
rect 29437 79 29460 113
rect 29494 79 29504 113
rect 29437 47 29504 79
rect 29534 143 29586 177
rect 29534 109 29544 143
rect 29578 109 29586 143
rect 29534 47 29586 109
rect 29651 119 29703 131
rect 29651 85 29659 119
rect 29693 85 29703 119
rect 29651 47 29703 85
rect 29733 93 29787 131
rect 29733 59 29743 93
rect 29777 59 29787 93
rect 29733 47 29787 59
rect 29817 119 29869 131
rect 29817 85 29827 119
rect 29861 85 29869 119
rect 29817 47 29869 85
rect 29937 89 30042 131
rect 29937 55 29949 89
rect 29983 55 30042 89
rect 29937 47 30042 55
rect 30072 119 30122 131
rect 30553 131 30603 175
rect 30281 119 30399 131
rect 30072 95 30137 119
rect 30072 61 30082 95
rect 30116 61 30137 95
rect 30072 47 30137 61
rect 30167 95 30233 119
rect 30167 61 30189 95
rect 30223 61 30233 95
rect 30167 47 30233 61
rect 30263 47 30399 119
rect 30429 47 30471 131
rect 30501 93 30603 131
rect 30501 59 30535 93
rect 30569 59 30603 93
rect 30501 47 30603 59
rect 30633 119 30687 175
rect 31283 132 31335 177
rect 30857 119 30907 131
rect 30633 89 30702 119
rect 30633 55 30647 89
rect 30681 55 30702 89
rect 30633 47 30702 55
rect 30732 93 30811 119
rect 30732 59 30757 93
rect 30791 59 30811 93
rect 30732 47 30811 59
rect 30841 47 30907 119
rect 30937 89 31056 131
rect 30937 55 30969 89
rect 31003 55 31056 89
rect 30937 47 31056 55
rect 31086 47 31147 131
rect 31177 109 31229 131
rect 31177 75 31187 109
rect 31221 75 31229 109
rect 31177 47 31229 75
rect 31283 98 31291 132
rect 31325 98 31335 132
rect 31283 47 31335 98
rect 31365 165 31417 177
rect 31365 131 31375 165
rect 31409 131 31417 165
rect 31568 131 31620 177
rect 31365 97 31417 131
rect 31365 63 31375 97
rect 31409 63 31417 97
rect 31365 47 31417 63
rect 31471 119 31523 131
rect 31471 85 31479 119
rect 31513 85 31523 119
rect 31471 47 31523 85
rect 31553 113 31620 131
rect 31553 79 31576 113
rect 31610 79 31620 113
rect 31553 47 31620 79
rect 31650 143 31702 177
rect 31650 109 31660 143
rect 31694 109 31702 143
rect 31650 47 31702 109
rect 31767 119 31819 131
rect 31767 85 31775 119
rect 31809 85 31819 119
rect 31767 47 31819 85
rect 31849 93 31903 131
rect 31849 59 31859 93
rect 31893 59 31903 93
rect 31849 47 31903 59
rect 31933 119 31985 131
rect 31933 85 31943 119
rect 31977 85 31985 119
rect 31933 47 31985 85
rect 32053 89 32158 131
rect 32053 55 32065 89
rect 32099 55 32158 89
rect 32053 47 32158 55
rect 32188 119 32238 131
rect 32669 131 32719 175
rect 32397 119 32515 131
rect 32188 95 32253 119
rect 32188 61 32198 95
rect 32232 61 32253 95
rect 32188 47 32253 61
rect 32283 95 32349 119
rect 32283 61 32305 95
rect 32339 61 32349 95
rect 32283 47 32349 61
rect 32379 47 32515 119
rect 32545 47 32587 131
rect 32617 93 32719 131
rect 32617 59 32651 93
rect 32685 59 32719 93
rect 32617 47 32719 59
rect 32749 119 32803 175
rect 33399 132 33451 177
rect 32973 119 33023 131
rect 32749 89 32818 119
rect 32749 55 32763 89
rect 32797 55 32818 89
rect 32749 47 32818 55
rect 32848 93 32927 119
rect 32848 59 32873 93
rect 32907 59 32927 93
rect 32848 47 32927 59
rect 32957 47 33023 119
rect 33053 89 33172 131
rect 33053 55 33085 89
rect 33119 55 33172 89
rect 33053 47 33172 55
rect 33202 47 33263 131
rect 33293 109 33345 131
rect 33293 75 33303 109
rect 33337 75 33345 109
rect 33293 47 33345 75
rect 33399 98 33407 132
rect 33441 98 33451 132
rect 33399 47 33451 98
rect 33481 165 33533 177
rect 33481 131 33491 165
rect 33525 131 33533 165
rect 33684 131 33736 177
rect 33481 97 33533 131
rect 33481 63 33491 97
rect 33525 63 33533 97
rect 33481 47 33533 63
rect 33587 119 33639 131
rect 33587 85 33595 119
rect 33629 85 33639 119
rect 33587 47 33639 85
rect 33669 113 33736 131
rect 33669 79 33692 113
rect 33726 79 33736 113
rect 33669 47 33736 79
rect 33766 143 33818 177
rect 33766 109 33776 143
rect 33810 109 33818 143
rect 33766 47 33818 109
rect 33883 119 33935 131
rect 33883 85 33891 119
rect 33925 85 33935 119
rect 33883 47 33935 85
rect 33965 93 34019 131
rect 33965 59 33975 93
rect 34009 59 34019 93
rect 33965 47 34019 59
rect 34049 119 34101 131
rect 34049 85 34059 119
rect 34093 85 34101 119
rect 34049 47 34101 85
rect 34169 89 34274 131
rect 34169 55 34181 89
rect 34215 55 34274 89
rect 34169 47 34274 55
rect 34304 119 34354 131
rect 34785 131 34835 175
rect 34513 119 34631 131
rect 34304 95 34369 119
rect 34304 61 34314 95
rect 34348 61 34369 95
rect 34304 47 34369 61
rect 34399 95 34465 119
rect 34399 61 34421 95
rect 34455 61 34465 95
rect 34399 47 34465 61
rect 34495 47 34631 119
rect 34661 47 34703 131
rect 34733 93 34835 131
rect 34733 59 34767 93
rect 34801 59 34835 93
rect 34733 47 34835 59
rect 34865 119 34919 175
rect 35515 132 35567 177
rect 35089 119 35139 131
rect 34865 89 34934 119
rect 34865 55 34879 89
rect 34913 55 34934 89
rect 34865 47 34934 55
rect 34964 93 35043 119
rect 34964 59 34989 93
rect 35023 59 35043 93
rect 34964 47 35043 59
rect 35073 47 35139 119
rect 35169 89 35288 131
rect 35169 55 35201 89
rect 35235 55 35288 89
rect 35169 47 35288 55
rect 35318 47 35379 131
rect 35409 109 35461 131
rect 35409 75 35419 109
rect 35453 75 35461 109
rect 35409 47 35461 75
rect 35515 98 35523 132
rect 35557 98 35567 132
rect 35515 47 35567 98
rect 35597 165 35649 177
rect 35597 131 35607 165
rect 35641 131 35649 165
rect 35800 131 35852 177
rect 35597 97 35649 131
rect 35597 63 35607 97
rect 35641 63 35649 97
rect 35597 47 35649 63
rect 35703 119 35755 131
rect 35703 85 35711 119
rect 35745 85 35755 119
rect 35703 47 35755 85
rect 35785 113 35852 131
rect 35785 79 35808 113
rect 35842 79 35852 113
rect 35785 47 35852 79
rect 35882 143 35934 177
rect 35882 109 35892 143
rect 35926 109 35934 143
rect 35882 47 35934 109
rect 35999 119 36051 131
rect 35999 85 36007 119
rect 36041 85 36051 119
rect 35999 47 36051 85
rect 36081 93 36135 131
rect 36081 59 36091 93
rect 36125 59 36135 93
rect 36081 47 36135 59
rect 36165 119 36217 131
rect 36165 85 36175 119
rect 36209 85 36217 119
rect 36165 47 36217 85
rect 36285 89 36390 131
rect 36285 55 36297 89
rect 36331 55 36390 89
rect 36285 47 36390 55
rect 36420 119 36470 131
rect 36901 131 36951 175
rect 36629 119 36747 131
rect 36420 95 36485 119
rect 36420 61 36430 95
rect 36464 61 36485 95
rect 36420 47 36485 61
rect 36515 95 36581 119
rect 36515 61 36537 95
rect 36571 61 36581 95
rect 36515 47 36581 61
rect 36611 47 36747 119
rect 36777 47 36819 131
rect 36849 93 36951 131
rect 36849 59 36883 93
rect 36917 59 36951 93
rect 36849 47 36951 59
rect 36981 119 37035 175
rect 37631 132 37683 177
rect 37205 119 37255 131
rect 36981 89 37050 119
rect 36981 55 36995 89
rect 37029 55 37050 89
rect 36981 47 37050 55
rect 37080 93 37159 119
rect 37080 59 37105 93
rect 37139 59 37159 93
rect 37080 47 37159 59
rect 37189 47 37255 119
rect 37285 89 37404 131
rect 37285 55 37317 89
rect 37351 55 37404 89
rect 37285 47 37404 55
rect 37434 47 37495 131
rect 37525 109 37577 131
rect 37525 75 37535 109
rect 37569 75 37577 109
rect 37525 47 37577 75
rect 37631 98 37639 132
rect 37673 98 37683 132
rect 37631 47 37683 98
rect 37713 165 37765 177
rect 37713 131 37723 165
rect 37757 131 37765 165
rect 37916 131 37968 177
rect 37713 97 37765 131
rect 37713 63 37723 97
rect 37757 63 37765 97
rect 37713 47 37765 63
rect 37819 119 37871 131
rect 37819 85 37827 119
rect 37861 85 37871 119
rect 37819 47 37871 85
rect 37901 113 37968 131
rect 37901 79 37924 113
rect 37958 79 37968 113
rect 37901 47 37968 79
rect 37998 143 38050 177
rect 37998 109 38008 143
rect 38042 109 38050 143
rect 37998 47 38050 109
rect 38115 119 38167 131
rect 38115 85 38123 119
rect 38157 85 38167 119
rect 38115 47 38167 85
rect 38197 93 38251 131
rect 38197 59 38207 93
rect 38241 59 38251 93
rect 38197 47 38251 59
rect 38281 119 38333 131
rect 38281 85 38291 119
rect 38325 85 38333 119
rect 38281 47 38333 85
rect 38401 89 38506 131
rect 38401 55 38413 89
rect 38447 55 38506 89
rect 38401 47 38506 55
rect 38536 119 38586 131
rect 39017 131 39067 175
rect 38745 119 38863 131
rect 38536 95 38601 119
rect 38536 61 38546 95
rect 38580 61 38601 95
rect 38536 47 38601 61
rect 38631 95 38697 119
rect 38631 61 38653 95
rect 38687 61 38697 95
rect 38631 47 38697 61
rect 38727 47 38863 119
rect 38893 47 38935 131
rect 38965 93 39067 131
rect 38965 59 38999 93
rect 39033 59 39067 93
rect 38965 47 39067 59
rect 39097 119 39151 175
rect 39747 132 39799 177
rect 39321 119 39371 131
rect 39097 89 39166 119
rect 39097 55 39111 89
rect 39145 55 39166 89
rect 39097 47 39166 55
rect 39196 93 39275 119
rect 39196 59 39221 93
rect 39255 59 39275 93
rect 39196 47 39275 59
rect 39305 47 39371 119
rect 39401 89 39520 131
rect 39401 55 39433 89
rect 39467 55 39520 89
rect 39401 47 39520 55
rect 39550 47 39611 131
rect 39641 109 39693 131
rect 39641 75 39651 109
rect 39685 75 39693 109
rect 39641 47 39693 75
rect 39747 98 39755 132
rect 39789 98 39799 132
rect 39747 47 39799 98
rect 39829 165 39881 177
rect 39829 131 39839 165
rect 39873 131 39881 165
rect 40032 131 40084 177
rect 39829 97 39881 131
rect 39829 63 39839 97
rect 39873 63 39881 97
rect 39829 47 39881 63
rect 39935 119 39987 131
rect 39935 85 39943 119
rect 39977 85 39987 119
rect 39935 47 39987 85
rect 40017 113 40084 131
rect 40017 79 40040 113
rect 40074 79 40084 113
rect 40017 47 40084 79
rect 40114 143 40166 177
rect 40114 109 40124 143
rect 40158 109 40166 143
rect 40114 47 40166 109
rect 40231 119 40283 131
rect 40231 85 40239 119
rect 40273 85 40283 119
rect 40231 47 40283 85
rect 40313 93 40367 131
rect 40313 59 40323 93
rect 40357 59 40367 93
rect 40313 47 40367 59
rect 40397 119 40449 131
rect 40397 85 40407 119
rect 40441 85 40449 119
rect 40397 47 40449 85
rect 40517 89 40622 131
rect 40517 55 40529 89
rect 40563 55 40622 89
rect 40517 47 40622 55
rect 40652 119 40702 131
rect 41133 131 41183 175
rect 40861 119 40979 131
rect 40652 95 40717 119
rect 40652 61 40662 95
rect 40696 61 40717 95
rect 40652 47 40717 61
rect 40747 95 40813 119
rect 40747 61 40769 95
rect 40803 61 40813 95
rect 40747 47 40813 61
rect 40843 47 40979 119
rect 41009 47 41051 131
rect 41081 93 41183 131
rect 41081 59 41115 93
rect 41149 59 41183 93
rect 41081 47 41183 59
rect 41213 119 41267 175
rect 41863 132 41915 177
rect 41437 119 41487 131
rect 41213 89 41282 119
rect 41213 55 41227 89
rect 41261 55 41282 89
rect 41213 47 41282 55
rect 41312 93 41391 119
rect 41312 59 41337 93
rect 41371 59 41391 93
rect 41312 47 41391 59
rect 41421 47 41487 119
rect 41517 89 41636 131
rect 41517 55 41549 89
rect 41583 55 41636 89
rect 41517 47 41636 55
rect 41666 47 41727 131
rect 41757 109 41809 131
rect 41757 75 41767 109
rect 41801 75 41809 109
rect 41757 47 41809 75
rect 41863 98 41871 132
rect 41905 98 41915 132
rect 41863 47 41915 98
rect 41945 165 41997 177
rect 41945 131 41955 165
rect 41989 131 41997 165
rect 42148 131 42200 177
rect 41945 97 41997 131
rect 41945 63 41955 97
rect 41989 63 41997 97
rect 41945 47 41997 63
rect 42051 119 42103 131
rect 42051 85 42059 119
rect 42093 85 42103 119
rect 42051 47 42103 85
rect 42133 113 42200 131
rect 42133 79 42156 113
rect 42190 79 42200 113
rect 42133 47 42200 79
rect 42230 143 42282 177
rect 42230 109 42240 143
rect 42274 109 42282 143
rect 42230 47 42282 109
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 378 485 430 497
rect 378 451 386 485
rect 420 451 430 485
rect 378 413 430 451
rect 460 477 522 497
rect 460 443 470 477
rect 504 443 522 477
rect 460 413 522 443
rect 552 483 621 497
rect 552 449 563 483
rect 597 449 621 483
rect 552 413 621 449
rect 651 459 761 497
rect 651 425 717 459
rect 751 425 761 459
rect 651 413 761 425
rect 791 475 858 497
rect 791 441 814 475
rect 848 441 858 475
rect 791 413 858 441
rect 888 459 940 497
rect 888 425 898 459
rect 932 425 940 459
rect 888 413 940 425
rect 1003 485 1055 497
rect 1003 451 1011 485
rect 1045 451 1055 485
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 1003 329 1055 451
rect 1085 477 1154 497
rect 1085 443 1099 477
rect 1133 443 1154 477
rect 1085 413 1154 443
rect 1184 484 1240 497
rect 1184 450 1196 484
rect 1230 450 1240 484
rect 1184 413 1240 450
rect 1270 413 1324 497
rect 1354 485 1432 497
rect 1354 451 1388 485
rect 1422 451 1432 485
rect 1354 413 1432 451
rect 1462 459 1516 497
rect 1462 425 1472 459
rect 1506 425 1516 459
rect 1462 413 1516 425
rect 1546 485 1680 497
rect 1546 451 1558 485
rect 1592 451 1636 485
rect 1670 451 1680 485
rect 1546 413 1680 451
rect 1085 329 1139 413
rect 1630 297 1680 413
rect 1710 477 1766 497
rect 1710 443 1720 477
rect 1754 443 1766 477
rect 1710 409 1766 443
rect 1710 375 1720 409
rect 1754 375 1766 409
rect 1710 341 1766 375
rect 1847 485 1899 497
rect 1847 451 1855 485
rect 1889 451 1899 485
rect 1847 417 1899 451
rect 1847 383 1855 417
rect 1889 383 1899 417
rect 1847 369 1899 383
rect 1929 485 1996 497
rect 1929 451 1952 485
rect 1986 451 1996 485
rect 1929 417 1996 451
rect 1929 383 1952 417
rect 1986 383 1996 417
rect 1929 369 1996 383
rect 1710 307 1720 341
rect 1754 307 1766 341
rect 1710 297 1766 307
rect 1944 349 1996 369
rect 1944 315 1952 349
rect 1986 315 1996 349
rect 1944 297 1996 315
rect 2026 449 2078 497
rect 2026 415 2036 449
rect 2070 415 2078 449
rect 2026 381 2078 415
rect 2026 347 2036 381
rect 2070 347 2078 381
rect 2143 477 2195 491
rect 2143 443 2151 477
rect 2185 443 2195 477
rect 2143 409 2195 443
rect 2143 375 2151 409
rect 2185 375 2195 409
rect 2143 363 2195 375
rect 2225 461 2279 491
rect 2225 427 2235 461
rect 2269 427 2279 461
rect 2225 363 2279 427
rect 2309 477 2361 491
rect 2309 443 2319 477
rect 2353 443 2361 477
rect 2309 409 2361 443
rect 2494 485 2546 497
rect 2494 451 2502 485
rect 2536 451 2546 485
rect 2494 413 2546 451
rect 2576 477 2638 497
rect 2576 443 2586 477
rect 2620 443 2638 477
rect 2576 413 2638 443
rect 2668 483 2737 497
rect 2668 449 2679 483
rect 2713 449 2737 483
rect 2668 413 2737 449
rect 2767 459 2877 497
rect 2767 425 2833 459
rect 2867 425 2877 459
rect 2767 413 2877 425
rect 2907 475 2974 497
rect 2907 441 2930 475
rect 2964 441 2974 475
rect 2907 413 2974 441
rect 3004 459 3056 497
rect 3004 425 3014 459
rect 3048 425 3056 459
rect 3004 413 3056 425
rect 3119 485 3171 497
rect 3119 451 3127 485
rect 3161 451 3171 485
rect 2309 375 2319 409
rect 2353 375 2361 409
rect 2309 363 2361 375
rect 2026 297 2078 347
rect 3119 329 3171 451
rect 3201 477 3270 497
rect 3201 443 3215 477
rect 3249 443 3270 477
rect 3201 413 3270 443
rect 3300 484 3356 497
rect 3300 450 3312 484
rect 3346 450 3356 484
rect 3300 413 3356 450
rect 3386 413 3440 497
rect 3470 485 3548 497
rect 3470 451 3504 485
rect 3538 451 3548 485
rect 3470 413 3548 451
rect 3578 459 3632 497
rect 3578 425 3588 459
rect 3622 425 3632 459
rect 3578 413 3632 425
rect 3662 485 3796 497
rect 3662 451 3674 485
rect 3708 451 3752 485
rect 3786 451 3796 485
rect 3662 413 3796 451
rect 3201 329 3255 413
rect 3746 297 3796 413
rect 3826 477 3882 497
rect 3826 443 3836 477
rect 3870 443 3882 477
rect 3826 409 3882 443
rect 3826 375 3836 409
rect 3870 375 3882 409
rect 3826 341 3882 375
rect 3963 485 4015 497
rect 3963 451 3971 485
rect 4005 451 4015 485
rect 3963 417 4015 451
rect 3963 383 3971 417
rect 4005 383 4015 417
rect 3963 369 4015 383
rect 4045 485 4112 497
rect 4045 451 4068 485
rect 4102 451 4112 485
rect 4045 417 4112 451
rect 4045 383 4068 417
rect 4102 383 4112 417
rect 4045 369 4112 383
rect 3826 307 3836 341
rect 3870 307 3882 341
rect 3826 297 3882 307
rect 4060 349 4112 369
rect 4060 315 4068 349
rect 4102 315 4112 349
rect 4060 297 4112 315
rect 4142 449 4194 497
rect 4142 415 4152 449
rect 4186 415 4194 449
rect 4142 381 4194 415
rect 4142 347 4152 381
rect 4186 347 4194 381
rect 4259 477 4311 491
rect 4259 443 4267 477
rect 4301 443 4311 477
rect 4259 409 4311 443
rect 4259 375 4267 409
rect 4301 375 4311 409
rect 4259 363 4311 375
rect 4341 461 4395 491
rect 4341 427 4351 461
rect 4385 427 4395 461
rect 4341 363 4395 427
rect 4425 477 4477 491
rect 4425 443 4435 477
rect 4469 443 4477 477
rect 4425 409 4477 443
rect 4610 485 4662 497
rect 4610 451 4618 485
rect 4652 451 4662 485
rect 4610 413 4662 451
rect 4692 477 4754 497
rect 4692 443 4702 477
rect 4736 443 4754 477
rect 4692 413 4754 443
rect 4784 483 4853 497
rect 4784 449 4795 483
rect 4829 449 4853 483
rect 4784 413 4853 449
rect 4883 459 4993 497
rect 4883 425 4949 459
rect 4983 425 4993 459
rect 4883 413 4993 425
rect 5023 475 5090 497
rect 5023 441 5046 475
rect 5080 441 5090 475
rect 5023 413 5090 441
rect 5120 459 5172 497
rect 5120 425 5130 459
rect 5164 425 5172 459
rect 5120 413 5172 425
rect 5235 485 5287 497
rect 5235 451 5243 485
rect 5277 451 5287 485
rect 4425 375 4435 409
rect 4469 375 4477 409
rect 4425 363 4477 375
rect 4142 297 4194 347
rect 5235 329 5287 451
rect 5317 477 5386 497
rect 5317 443 5331 477
rect 5365 443 5386 477
rect 5317 413 5386 443
rect 5416 484 5472 497
rect 5416 450 5428 484
rect 5462 450 5472 484
rect 5416 413 5472 450
rect 5502 413 5556 497
rect 5586 485 5664 497
rect 5586 451 5620 485
rect 5654 451 5664 485
rect 5586 413 5664 451
rect 5694 459 5748 497
rect 5694 425 5704 459
rect 5738 425 5748 459
rect 5694 413 5748 425
rect 5778 485 5912 497
rect 5778 451 5790 485
rect 5824 451 5868 485
rect 5902 451 5912 485
rect 5778 413 5912 451
rect 5317 329 5371 413
rect 5862 297 5912 413
rect 5942 477 5998 497
rect 5942 443 5952 477
rect 5986 443 5998 477
rect 5942 409 5998 443
rect 5942 375 5952 409
rect 5986 375 5998 409
rect 5942 341 5998 375
rect 6079 485 6131 497
rect 6079 451 6087 485
rect 6121 451 6131 485
rect 6079 417 6131 451
rect 6079 383 6087 417
rect 6121 383 6131 417
rect 6079 369 6131 383
rect 6161 485 6228 497
rect 6161 451 6184 485
rect 6218 451 6228 485
rect 6161 417 6228 451
rect 6161 383 6184 417
rect 6218 383 6228 417
rect 6161 369 6228 383
rect 5942 307 5952 341
rect 5986 307 5998 341
rect 5942 297 5998 307
rect 6176 349 6228 369
rect 6176 315 6184 349
rect 6218 315 6228 349
rect 6176 297 6228 315
rect 6258 449 6310 497
rect 6258 415 6268 449
rect 6302 415 6310 449
rect 6258 381 6310 415
rect 6258 347 6268 381
rect 6302 347 6310 381
rect 6375 477 6427 491
rect 6375 443 6383 477
rect 6417 443 6427 477
rect 6375 409 6427 443
rect 6375 375 6383 409
rect 6417 375 6427 409
rect 6375 363 6427 375
rect 6457 461 6511 491
rect 6457 427 6467 461
rect 6501 427 6511 461
rect 6457 363 6511 427
rect 6541 477 6593 491
rect 6541 443 6551 477
rect 6585 443 6593 477
rect 6541 409 6593 443
rect 6726 485 6778 497
rect 6726 451 6734 485
rect 6768 451 6778 485
rect 6726 413 6778 451
rect 6808 477 6870 497
rect 6808 443 6818 477
rect 6852 443 6870 477
rect 6808 413 6870 443
rect 6900 483 6969 497
rect 6900 449 6911 483
rect 6945 449 6969 483
rect 6900 413 6969 449
rect 6999 459 7109 497
rect 6999 425 7065 459
rect 7099 425 7109 459
rect 6999 413 7109 425
rect 7139 475 7206 497
rect 7139 441 7162 475
rect 7196 441 7206 475
rect 7139 413 7206 441
rect 7236 459 7288 497
rect 7236 425 7246 459
rect 7280 425 7288 459
rect 7236 413 7288 425
rect 7351 485 7403 497
rect 7351 451 7359 485
rect 7393 451 7403 485
rect 6541 375 6551 409
rect 6585 375 6593 409
rect 6541 363 6593 375
rect 6258 297 6310 347
rect 7351 329 7403 451
rect 7433 477 7502 497
rect 7433 443 7447 477
rect 7481 443 7502 477
rect 7433 413 7502 443
rect 7532 484 7588 497
rect 7532 450 7544 484
rect 7578 450 7588 484
rect 7532 413 7588 450
rect 7618 413 7672 497
rect 7702 485 7780 497
rect 7702 451 7736 485
rect 7770 451 7780 485
rect 7702 413 7780 451
rect 7810 459 7864 497
rect 7810 425 7820 459
rect 7854 425 7864 459
rect 7810 413 7864 425
rect 7894 485 8028 497
rect 7894 451 7906 485
rect 7940 451 7984 485
rect 8018 451 8028 485
rect 7894 413 8028 451
rect 7433 329 7487 413
rect 7978 297 8028 413
rect 8058 477 8114 497
rect 8058 443 8068 477
rect 8102 443 8114 477
rect 8058 409 8114 443
rect 8058 375 8068 409
rect 8102 375 8114 409
rect 8058 341 8114 375
rect 8195 485 8247 497
rect 8195 451 8203 485
rect 8237 451 8247 485
rect 8195 417 8247 451
rect 8195 383 8203 417
rect 8237 383 8247 417
rect 8195 369 8247 383
rect 8277 485 8344 497
rect 8277 451 8300 485
rect 8334 451 8344 485
rect 8277 417 8344 451
rect 8277 383 8300 417
rect 8334 383 8344 417
rect 8277 369 8344 383
rect 8058 307 8068 341
rect 8102 307 8114 341
rect 8058 297 8114 307
rect 8292 349 8344 369
rect 8292 315 8300 349
rect 8334 315 8344 349
rect 8292 297 8344 315
rect 8374 449 8426 497
rect 8374 415 8384 449
rect 8418 415 8426 449
rect 8374 381 8426 415
rect 8374 347 8384 381
rect 8418 347 8426 381
rect 8491 477 8543 491
rect 8491 443 8499 477
rect 8533 443 8543 477
rect 8491 409 8543 443
rect 8491 375 8499 409
rect 8533 375 8543 409
rect 8491 363 8543 375
rect 8573 461 8627 491
rect 8573 427 8583 461
rect 8617 427 8627 461
rect 8573 363 8627 427
rect 8657 477 8709 491
rect 8657 443 8667 477
rect 8701 443 8709 477
rect 8657 409 8709 443
rect 8842 485 8894 497
rect 8842 451 8850 485
rect 8884 451 8894 485
rect 8842 413 8894 451
rect 8924 477 8986 497
rect 8924 443 8934 477
rect 8968 443 8986 477
rect 8924 413 8986 443
rect 9016 483 9085 497
rect 9016 449 9027 483
rect 9061 449 9085 483
rect 9016 413 9085 449
rect 9115 459 9225 497
rect 9115 425 9181 459
rect 9215 425 9225 459
rect 9115 413 9225 425
rect 9255 475 9322 497
rect 9255 441 9278 475
rect 9312 441 9322 475
rect 9255 413 9322 441
rect 9352 459 9404 497
rect 9352 425 9362 459
rect 9396 425 9404 459
rect 9352 413 9404 425
rect 9467 485 9519 497
rect 9467 451 9475 485
rect 9509 451 9519 485
rect 8657 375 8667 409
rect 8701 375 8709 409
rect 8657 363 8709 375
rect 8374 297 8426 347
rect 9467 329 9519 451
rect 9549 477 9618 497
rect 9549 443 9563 477
rect 9597 443 9618 477
rect 9549 413 9618 443
rect 9648 484 9704 497
rect 9648 450 9660 484
rect 9694 450 9704 484
rect 9648 413 9704 450
rect 9734 413 9788 497
rect 9818 485 9896 497
rect 9818 451 9852 485
rect 9886 451 9896 485
rect 9818 413 9896 451
rect 9926 459 9980 497
rect 9926 425 9936 459
rect 9970 425 9980 459
rect 9926 413 9980 425
rect 10010 485 10144 497
rect 10010 451 10022 485
rect 10056 451 10100 485
rect 10134 451 10144 485
rect 10010 413 10144 451
rect 9549 329 9603 413
rect 10094 297 10144 413
rect 10174 477 10230 497
rect 10174 443 10184 477
rect 10218 443 10230 477
rect 10174 409 10230 443
rect 10174 375 10184 409
rect 10218 375 10230 409
rect 10174 341 10230 375
rect 10311 485 10363 497
rect 10311 451 10319 485
rect 10353 451 10363 485
rect 10311 417 10363 451
rect 10311 383 10319 417
rect 10353 383 10363 417
rect 10311 369 10363 383
rect 10393 485 10460 497
rect 10393 451 10416 485
rect 10450 451 10460 485
rect 10393 417 10460 451
rect 10393 383 10416 417
rect 10450 383 10460 417
rect 10393 369 10460 383
rect 10174 307 10184 341
rect 10218 307 10230 341
rect 10174 297 10230 307
rect 10408 349 10460 369
rect 10408 315 10416 349
rect 10450 315 10460 349
rect 10408 297 10460 315
rect 10490 449 10542 497
rect 10490 415 10500 449
rect 10534 415 10542 449
rect 10490 381 10542 415
rect 10490 347 10500 381
rect 10534 347 10542 381
rect 10607 477 10659 491
rect 10607 443 10615 477
rect 10649 443 10659 477
rect 10607 409 10659 443
rect 10607 375 10615 409
rect 10649 375 10659 409
rect 10607 363 10659 375
rect 10689 461 10743 491
rect 10689 427 10699 461
rect 10733 427 10743 461
rect 10689 363 10743 427
rect 10773 477 10825 491
rect 10773 443 10783 477
rect 10817 443 10825 477
rect 10773 409 10825 443
rect 10958 485 11010 497
rect 10958 451 10966 485
rect 11000 451 11010 485
rect 10958 413 11010 451
rect 11040 477 11102 497
rect 11040 443 11050 477
rect 11084 443 11102 477
rect 11040 413 11102 443
rect 11132 483 11201 497
rect 11132 449 11143 483
rect 11177 449 11201 483
rect 11132 413 11201 449
rect 11231 459 11341 497
rect 11231 425 11297 459
rect 11331 425 11341 459
rect 11231 413 11341 425
rect 11371 475 11438 497
rect 11371 441 11394 475
rect 11428 441 11438 475
rect 11371 413 11438 441
rect 11468 459 11520 497
rect 11468 425 11478 459
rect 11512 425 11520 459
rect 11468 413 11520 425
rect 11583 485 11635 497
rect 11583 451 11591 485
rect 11625 451 11635 485
rect 10773 375 10783 409
rect 10817 375 10825 409
rect 10773 363 10825 375
rect 10490 297 10542 347
rect 11583 329 11635 451
rect 11665 477 11734 497
rect 11665 443 11679 477
rect 11713 443 11734 477
rect 11665 413 11734 443
rect 11764 484 11820 497
rect 11764 450 11776 484
rect 11810 450 11820 484
rect 11764 413 11820 450
rect 11850 413 11904 497
rect 11934 485 12012 497
rect 11934 451 11968 485
rect 12002 451 12012 485
rect 11934 413 12012 451
rect 12042 459 12096 497
rect 12042 425 12052 459
rect 12086 425 12096 459
rect 12042 413 12096 425
rect 12126 485 12260 497
rect 12126 451 12138 485
rect 12172 451 12216 485
rect 12250 451 12260 485
rect 12126 413 12260 451
rect 11665 329 11719 413
rect 12210 297 12260 413
rect 12290 477 12346 497
rect 12290 443 12300 477
rect 12334 443 12346 477
rect 12290 409 12346 443
rect 12290 375 12300 409
rect 12334 375 12346 409
rect 12290 341 12346 375
rect 12427 485 12479 497
rect 12427 451 12435 485
rect 12469 451 12479 485
rect 12427 417 12479 451
rect 12427 383 12435 417
rect 12469 383 12479 417
rect 12427 369 12479 383
rect 12509 485 12576 497
rect 12509 451 12532 485
rect 12566 451 12576 485
rect 12509 417 12576 451
rect 12509 383 12532 417
rect 12566 383 12576 417
rect 12509 369 12576 383
rect 12290 307 12300 341
rect 12334 307 12346 341
rect 12290 297 12346 307
rect 12524 349 12576 369
rect 12524 315 12532 349
rect 12566 315 12576 349
rect 12524 297 12576 315
rect 12606 449 12658 497
rect 12606 415 12616 449
rect 12650 415 12658 449
rect 12606 381 12658 415
rect 12606 347 12616 381
rect 12650 347 12658 381
rect 12723 477 12775 491
rect 12723 443 12731 477
rect 12765 443 12775 477
rect 12723 409 12775 443
rect 12723 375 12731 409
rect 12765 375 12775 409
rect 12723 363 12775 375
rect 12805 461 12859 491
rect 12805 427 12815 461
rect 12849 427 12859 461
rect 12805 363 12859 427
rect 12889 477 12941 491
rect 12889 443 12899 477
rect 12933 443 12941 477
rect 12889 409 12941 443
rect 13074 485 13126 497
rect 13074 451 13082 485
rect 13116 451 13126 485
rect 13074 413 13126 451
rect 13156 477 13218 497
rect 13156 443 13166 477
rect 13200 443 13218 477
rect 13156 413 13218 443
rect 13248 483 13317 497
rect 13248 449 13259 483
rect 13293 449 13317 483
rect 13248 413 13317 449
rect 13347 459 13457 497
rect 13347 425 13413 459
rect 13447 425 13457 459
rect 13347 413 13457 425
rect 13487 475 13554 497
rect 13487 441 13510 475
rect 13544 441 13554 475
rect 13487 413 13554 441
rect 13584 459 13636 497
rect 13584 425 13594 459
rect 13628 425 13636 459
rect 13584 413 13636 425
rect 13699 485 13751 497
rect 13699 451 13707 485
rect 13741 451 13751 485
rect 12889 375 12899 409
rect 12933 375 12941 409
rect 12889 363 12941 375
rect 12606 297 12658 347
rect 13699 329 13751 451
rect 13781 477 13850 497
rect 13781 443 13795 477
rect 13829 443 13850 477
rect 13781 413 13850 443
rect 13880 484 13936 497
rect 13880 450 13892 484
rect 13926 450 13936 484
rect 13880 413 13936 450
rect 13966 413 14020 497
rect 14050 485 14128 497
rect 14050 451 14084 485
rect 14118 451 14128 485
rect 14050 413 14128 451
rect 14158 459 14212 497
rect 14158 425 14168 459
rect 14202 425 14212 459
rect 14158 413 14212 425
rect 14242 485 14376 497
rect 14242 451 14254 485
rect 14288 451 14332 485
rect 14366 451 14376 485
rect 14242 413 14376 451
rect 13781 329 13835 413
rect 14326 297 14376 413
rect 14406 477 14462 497
rect 14406 443 14416 477
rect 14450 443 14462 477
rect 14406 409 14462 443
rect 14406 375 14416 409
rect 14450 375 14462 409
rect 14406 341 14462 375
rect 14543 485 14595 497
rect 14543 451 14551 485
rect 14585 451 14595 485
rect 14543 417 14595 451
rect 14543 383 14551 417
rect 14585 383 14595 417
rect 14543 369 14595 383
rect 14625 485 14692 497
rect 14625 451 14648 485
rect 14682 451 14692 485
rect 14625 417 14692 451
rect 14625 383 14648 417
rect 14682 383 14692 417
rect 14625 369 14692 383
rect 14406 307 14416 341
rect 14450 307 14462 341
rect 14406 297 14462 307
rect 14640 349 14692 369
rect 14640 315 14648 349
rect 14682 315 14692 349
rect 14640 297 14692 315
rect 14722 449 14774 497
rect 14722 415 14732 449
rect 14766 415 14774 449
rect 14722 381 14774 415
rect 14722 347 14732 381
rect 14766 347 14774 381
rect 14839 477 14891 491
rect 14839 443 14847 477
rect 14881 443 14891 477
rect 14839 409 14891 443
rect 14839 375 14847 409
rect 14881 375 14891 409
rect 14839 363 14891 375
rect 14921 461 14975 491
rect 14921 427 14931 461
rect 14965 427 14975 461
rect 14921 363 14975 427
rect 15005 477 15057 491
rect 15005 443 15015 477
rect 15049 443 15057 477
rect 15005 409 15057 443
rect 15190 485 15242 497
rect 15190 451 15198 485
rect 15232 451 15242 485
rect 15190 413 15242 451
rect 15272 477 15334 497
rect 15272 443 15282 477
rect 15316 443 15334 477
rect 15272 413 15334 443
rect 15364 483 15433 497
rect 15364 449 15375 483
rect 15409 449 15433 483
rect 15364 413 15433 449
rect 15463 459 15573 497
rect 15463 425 15529 459
rect 15563 425 15573 459
rect 15463 413 15573 425
rect 15603 475 15670 497
rect 15603 441 15626 475
rect 15660 441 15670 475
rect 15603 413 15670 441
rect 15700 459 15752 497
rect 15700 425 15710 459
rect 15744 425 15752 459
rect 15700 413 15752 425
rect 15815 485 15867 497
rect 15815 451 15823 485
rect 15857 451 15867 485
rect 15005 375 15015 409
rect 15049 375 15057 409
rect 15005 363 15057 375
rect 14722 297 14774 347
rect 15815 329 15867 451
rect 15897 477 15966 497
rect 15897 443 15911 477
rect 15945 443 15966 477
rect 15897 413 15966 443
rect 15996 484 16052 497
rect 15996 450 16008 484
rect 16042 450 16052 484
rect 15996 413 16052 450
rect 16082 413 16136 497
rect 16166 485 16244 497
rect 16166 451 16200 485
rect 16234 451 16244 485
rect 16166 413 16244 451
rect 16274 459 16328 497
rect 16274 425 16284 459
rect 16318 425 16328 459
rect 16274 413 16328 425
rect 16358 485 16492 497
rect 16358 451 16370 485
rect 16404 451 16448 485
rect 16482 451 16492 485
rect 16358 413 16492 451
rect 15897 329 15951 413
rect 16442 297 16492 413
rect 16522 477 16578 497
rect 16522 443 16532 477
rect 16566 443 16578 477
rect 16522 409 16578 443
rect 16522 375 16532 409
rect 16566 375 16578 409
rect 16522 341 16578 375
rect 16659 485 16711 497
rect 16659 451 16667 485
rect 16701 451 16711 485
rect 16659 417 16711 451
rect 16659 383 16667 417
rect 16701 383 16711 417
rect 16659 369 16711 383
rect 16741 485 16808 497
rect 16741 451 16764 485
rect 16798 451 16808 485
rect 16741 417 16808 451
rect 16741 383 16764 417
rect 16798 383 16808 417
rect 16741 369 16808 383
rect 16522 307 16532 341
rect 16566 307 16578 341
rect 16522 297 16578 307
rect 16756 349 16808 369
rect 16756 315 16764 349
rect 16798 315 16808 349
rect 16756 297 16808 315
rect 16838 449 16890 497
rect 16838 415 16848 449
rect 16882 415 16890 449
rect 16838 381 16890 415
rect 16838 347 16848 381
rect 16882 347 16890 381
rect 16955 477 17007 491
rect 16955 443 16963 477
rect 16997 443 17007 477
rect 16955 409 17007 443
rect 16955 375 16963 409
rect 16997 375 17007 409
rect 16955 363 17007 375
rect 17037 461 17091 491
rect 17037 427 17047 461
rect 17081 427 17091 461
rect 17037 363 17091 427
rect 17121 477 17173 491
rect 17121 443 17131 477
rect 17165 443 17173 477
rect 17121 409 17173 443
rect 17306 485 17358 497
rect 17306 451 17314 485
rect 17348 451 17358 485
rect 17306 413 17358 451
rect 17388 477 17450 497
rect 17388 443 17398 477
rect 17432 443 17450 477
rect 17388 413 17450 443
rect 17480 483 17549 497
rect 17480 449 17491 483
rect 17525 449 17549 483
rect 17480 413 17549 449
rect 17579 459 17689 497
rect 17579 425 17645 459
rect 17679 425 17689 459
rect 17579 413 17689 425
rect 17719 475 17786 497
rect 17719 441 17742 475
rect 17776 441 17786 475
rect 17719 413 17786 441
rect 17816 459 17868 497
rect 17816 425 17826 459
rect 17860 425 17868 459
rect 17816 413 17868 425
rect 17931 485 17983 497
rect 17931 451 17939 485
rect 17973 451 17983 485
rect 17121 375 17131 409
rect 17165 375 17173 409
rect 17121 363 17173 375
rect 16838 297 16890 347
rect 17931 329 17983 451
rect 18013 477 18082 497
rect 18013 443 18027 477
rect 18061 443 18082 477
rect 18013 413 18082 443
rect 18112 484 18168 497
rect 18112 450 18124 484
rect 18158 450 18168 484
rect 18112 413 18168 450
rect 18198 413 18252 497
rect 18282 485 18360 497
rect 18282 451 18316 485
rect 18350 451 18360 485
rect 18282 413 18360 451
rect 18390 459 18444 497
rect 18390 425 18400 459
rect 18434 425 18444 459
rect 18390 413 18444 425
rect 18474 485 18608 497
rect 18474 451 18486 485
rect 18520 451 18564 485
rect 18598 451 18608 485
rect 18474 413 18608 451
rect 18013 329 18067 413
rect 18558 297 18608 413
rect 18638 477 18694 497
rect 18638 443 18648 477
rect 18682 443 18694 477
rect 18638 409 18694 443
rect 18638 375 18648 409
rect 18682 375 18694 409
rect 18638 341 18694 375
rect 18775 485 18827 497
rect 18775 451 18783 485
rect 18817 451 18827 485
rect 18775 417 18827 451
rect 18775 383 18783 417
rect 18817 383 18827 417
rect 18775 369 18827 383
rect 18857 485 18924 497
rect 18857 451 18880 485
rect 18914 451 18924 485
rect 18857 417 18924 451
rect 18857 383 18880 417
rect 18914 383 18924 417
rect 18857 369 18924 383
rect 18638 307 18648 341
rect 18682 307 18694 341
rect 18638 297 18694 307
rect 18872 349 18924 369
rect 18872 315 18880 349
rect 18914 315 18924 349
rect 18872 297 18924 315
rect 18954 449 19006 497
rect 18954 415 18964 449
rect 18998 415 19006 449
rect 18954 381 19006 415
rect 18954 347 18964 381
rect 18998 347 19006 381
rect 19071 477 19123 491
rect 19071 443 19079 477
rect 19113 443 19123 477
rect 19071 409 19123 443
rect 19071 375 19079 409
rect 19113 375 19123 409
rect 19071 363 19123 375
rect 19153 461 19207 491
rect 19153 427 19163 461
rect 19197 427 19207 461
rect 19153 363 19207 427
rect 19237 477 19289 491
rect 19237 443 19247 477
rect 19281 443 19289 477
rect 19237 409 19289 443
rect 19422 485 19474 497
rect 19422 451 19430 485
rect 19464 451 19474 485
rect 19422 413 19474 451
rect 19504 477 19566 497
rect 19504 443 19514 477
rect 19548 443 19566 477
rect 19504 413 19566 443
rect 19596 483 19665 497
rect 19596 449 19607 483
rect 19641 449 19665 483
rect 19596 413 19665 449
rect 19695 459 19805 497
rect 19695 425 19761 459
rect 19795 425 19805 459
rect 19695 413 19805 425
rect 19835 475 19902 497
rect 19835 441 19858 475
rect 19892 441 19902 475
rect 19835 413 19902 441
rect 19932 459 19984 497
rect 19932 425 19942 459
rect 19976 425 19984 459
rect 19932 413 19984 425
rect 20047 485 20099 497
rect 20047 451 20055 485
rect 20089 451 20099 485
rect 19237 375 19247 409
rect 19281 375 19289 409
rect 19237 363 19289 375
rect 18954 297 19006 347
rect 20047 329 20099 451
rect 20129 477 20198 497
rect 20129 443 20143 477
rect 20177 443 20198 477
rect 20129 413 20198 443
rect 20228 484 20284 497
rect 20228 450 20240 484
rect 20274 450 20284 484
rect 20228 413 20284 450
rect 20314 413 20368 497
rect 20398 485 20476 497
rect 20398 451 20432 485
rect 20466 451 20476 485
rect 20398 413 20476 451
rect 20506 459 20560 497
rect 20506 425 20516 459
rect 20550 425 20560 459
rect 20506 413 20560 425
rect 20590 485 20724 497
rect 20590 451 20602 485
rect 20636 451 20680 485
rect 20714 451 20724 485
rect 20590 413 20724 451
rect 20129 329 20183 413
rect 20674 297 20724 413
rect 20754 477 20810 497
rect 20754 443 20764 477
rect 20798 443 20810 477
rect 20754 409 20810 443
rect 20754 375 20764 409
rect 20798 375 20810 409
rect 20754 341 20810 375
rect 20891 485 20943 497
rect 20891 451 20899 485
rect 20933 451 20943 485
rect 20891 417 20943 451
rect 20891 383 20899 417
rect 20933 383 20943 417
rect 20891 369 20943 383
rect 20973 485 21040 497
rect 20973 451 20996 485
rect 21030 451 21040 485
rect 20973 417 21040 451
rect 20973 383 20996 417
rect 21030 383 21040 417
rect 20973 369 21040 383
rect 20754 307 20764 341
rect 20798 307 20810 341
rect 20754 297 20810 307
rect 20988 349 21040 369
rect 20988 315 20996 349
rect 21030 315 21040 349
rect 20988 297 21040 315
rect 21070 449 21122 497
rect 21070 415 21080 449
rect 21114 415 21122 449
rect 21070 381 21122 415
rect 21070 347 21080 381
rect 21114 347 21122 381
rect 21187 477 21239 491
rect 21187 443 21195 477
rect 21229 443 21239 477
rect 21187 409 21239 443
rect 21187 375 21195 409
rect 21229 375 21239 409
rect 21187 363 21239 375
rect 21269 461 21323 491
rect 21269 427 21279 461
rect 21313 427 21323 461
rect 21269 363 21323 427
rect 21353 477 21405 491
rect 21353 443 21363 477
rect 21397 443 21405 477
rect 21353 409 21405 443
rect 21538 485 21590 497
rect 21538 451 21546 485
rect 21580 451 21590 485
rect 21538 413 21590 451
rect 21620 477 21682 497
rect 21620 443 21630 477
rect 21664 443 21682 477
rect 21620 413 21682 443
rect 21712 483 21781 497
rect 21712 449 21723 483
rect 21757 449 21781 483
rect 21712 413 21781 449
rect 21811 459 21921 497
rect 21811 425 21877 459
rect 21911 425 21921 459
rect 21811 413 21921 425
rect 21951 475 22018 497
rect 21951 441 21974 475
rect 22008 441 22018 475
rect 21951 413 22018 441
rect 22048 459 22100 497
rect 22048 425 22058 459
rect 22092 425 22100 459
rect 22048 413 22100 425
rect 22163 485 22215 497
rect 22163 451 22171 485
rect 22205 451 22215 485
rect 21353 375 21363 409
rect 21397 375 21405 409
rect 21353 363 21405 375
rect 21070 297 21122 347
rect 22163 329 22215 451
rect 22245 477 22314 497
rect 22245 443 22259 477
rect 22293 443 22314 477
rect 22245 413 22314 443
rect 22344 484 22400 497
rect 22344 450 22356 484
rect 22390 450 22400 484
rect 22344 413 22400 450
rect 22430 413 22484 497
rect 22514 485 22592 497
rect 22514 451 22548 485
rect 22582 451 22592 485
rect 22514 413 22592 451
rect 22622 459 22676 497
rect 22622 425 22632 459
rect 22666 425 22676 459
rect 22622 413 22676 425
rect 22706 485 22840 497
rect 22706 451 22718 485
rect 22752 451 22796 485
rect 22830 451 22840 485
rect 22706 413 22840 451
rect 22245 329 22299 413
rect 22790 297 22840 413
rect 22870 477 22926 497
rect 22870 443 22880 477
rect 22914 443 22926 477
rect 22870 409 22926 443
rect 22870 375 22880 409
rect 22914 375 22926 409
rect 22870 341 22926 375
rect 23007 485 23059 497
rect 23007 451 23015 485
rect 23049 451 23059 485
rect 23007 417 23059 451
rect 23007 383 23015 417
rect 23049 383 23059 417
rect 23007 369 23059 383
rect 23089 485 23156 497
rect 23089 451 23112 485
rect 23146 451 23156 485
rect 23089 417 23156 451
rect 23089 383 23112 417
rect 23146 383 23156 417
rect 23089 369 23156 383
rect 22870 307 22880 341
rect 22914 307 22926 341
rect 22870 297 22926 307
rect 23104 349 23156 369
rect 23104 315 23112 349
rect 23146 315 23156 349
rect 23104 297 23156 315
rect 23186 449 23238 497
rect 23186 415 23196 449
rect 23230 415 23238 449
rect 23186 381 23238 415
rect 23186 347 23196 381
rect 23230 347 23238 381
rect 23303 477 23355 491
rect 23303 443 23311 477
rect 23345 443 23355 477
rect 23303 409 23355 443
rect 23303 375 23311 409
rect 23345 375 23355 409
rect 23303 363 23355 375
rect 23385 461 23439 491
rect 23385 427 23395 461
rect 23429 427 23439 461
rect 23385 363 23439 427
rect 23469 477 23521 491
rect 23469 443 23479 477
rect 23513 443 23521 477
rect 23469 409 23521 443
rect 23654 485 23706 497
rect 23654 451 23662 485
rect 23696 451 23706 485
rect 23654 413 23706 451
rect 23736 477 23798 497
rect 23736 443 23746 477
rect 23780 443 23798 477
rect 23736 413 23798 443
rect 23828 483 23897 497
rect 23828 449 23839 483
rect 23873 449 23897 483
rect 23828 413 23897 449
rect 23927 459 24037 497
rect 23927 425 23993 459
rect 24027 425 24037 459
rect 23927 413 24037 425
rect 24067 475 24134 497
rect 24067 441 24090 475
rect 24124 441 24134 475
rect 24067 413 24134 441
rect 24164 459 24216 497
rect 24164 425 24174 459
rect 24208 425 24216 459
rect 24164 413 24216 425
rect 24279 485 24331 497
rect 24279 451 24287 485
rect 24321 451 24331 485
rect 23469 375 23479 409
rect 23513 375 23521 409
rect 23469 363 23521 375
rect 23186 297 23238 347
rect 24279 329 24331 451
rect 24361 477 24430 497
rect 24361 443 24375 477
rect 24409 443 24430 477
rect 24361 413 24430 443
rect 24460 484 24516 497
rect 24460 450 24472 484
rect 24506 450 24516 484
rect 24460 413 24516 450
rect 24546 413 24600 497
rect 24630 485 24708 497
rect 24630 451 24664 485
rect 24698 451 24708 485
rect 24630 413 24708 451
rect 24738 459 24792 497
rect 24738 425 24748 459
rect 24782 425 24792 459
rect 24738 413 24792 425
rect 24822 485 24956 497
rect 24822 451 24834 485
rect 24868 451 24912 485
rect 24946 451 24956 485
rect 24822 413 24956 451
rect 24361 329 24415 413
rect 24906 297 24956 413
rect 24986 477 25042 497
rect 24986 443 24996 477
rect 25030 443 25042 477
rect 24986 409 25042 443
rect 24986 375 24996 409
rect 25030 375 25042 409
rect 24986 341 25042 375
rect 25123 485 25175 497
rect 25123 451 25131 485
rect 25165 451 25175 485
rect 25123 417 25175 451
rect 25123 383 25131 417
rect 25165 383 25175 417
rect 25123 369 25175 383
rect 25205 485 25272 497
rect 25205 451 25228 485
rect 25262 451 25272 485
rect 25205 417 25272 451
rect 25205 383 25228 417
rect 25262 383 25272 417
rect 25205 369 25272 383
rect 24986 307 24996 341
rect 25030 307 25042 341
rect 24986 297 25042 307
rect 25220 349 25272 369
rect 25220 315 25228 349
rect 25262 315 25272 349
rect 25220 297 25272 315
rect 25302 449 25354 497
rect 25302 415 25312 449
rect 25346 415 25354 449
rect 25302 381 25354 415
rect 25302 347 25312 381
rect 25346 347 25354 381
rect 25419 477 25471 491
rect 25419 443 25427 477
rect 25461 443 25471 477
rect 25419 409 25471 443
rect 25419 375 25427 409
rect 25461 375 25471 409
rect 25419 363 25471 375
rect 25501 461 25555 491
rect 25501 427 25511 461
rect 25545 427 25555 461
rect 25501 363 25555 427
rect 25585 477 25637 491
rect 25585 443 25595 477
rect 25629 443 25637 477
rect 25585 409 25637 443
rect 25770 485 25822 497
rect 25770 451 25778 485
rect 25812 451 25822 485
rect 25770 413 25822 451
rect 25852 477 25914 497
rect 25852 443 25862 477
rect 25896 443 25914 477
rect 25852 413 25914 443
rect 25944 483 26013 497
rect 25944 449 25955 483
rect 25989 449 26013 483
rect 25944 413 26013 449
rect 26043 459 26153 497
rect 26043 425 26109 459
rect 26143 425 26153 459
rect 26043 413 26153 425
rect 26183 475 26250 497
rect 26183 441 26206 475
rect 26240 441 26250 475
rect 26183 413 26250 441
rect 26280 459 26332 497
rect 26280 425 26290 459
rect 26324 425 26332 459
rect 26280 413 26332 425
rect 26395 485 26447 497
rect 26395 451 26403 485
rect 26437 451 26447 485
rect 25585 375 25595 409
rect 25629 375 25637 409
rect 25585 363 25637 375
rect 25302 297 25354 347
rect 26395 329 26447 451
rect 26477 477 26546 497
rect 26477 443 26491 477
rect 26525 443 26546 477
rect 26477 413 26546 443
rect 26576 484 26632 497
rect 26576 450 26588 484
rect 26622 450 26632 484
rect 26576 413 26632 450
rect 26662 413 26716 497
rect 26746 485 26824 497
rect 26746 451 26780 485
rect 26814 451 26824 485
rect 26746 413 26824 451
rect 26854 459 26908 497
rect 26854 425 26864 459
rect 26898 425 26908 459
rect 26854 413 26908 425
rect 26938 485 27072 497
rect 26938 451 26950 485
rect 26984 451 27028 485
rect 27062 451 27072 485
rect 26938 413 27072 451
rect 26477 329 26531 413
rect 27022 297 27072 413
rect 27102 477 27158 497
rect 27102 443 27112 477
rect 27146 443 27158 477
rect 27102 409 27158 443
rect 27102 375 27112 409
rect 27146 375 27158 409
rect 27102 341 27158 375
rect 27239 485 27291 497
rect 27239 451 27247 485
rect 27281 451 27291 485
rect 27239 417 27291 451
rect 27239 383 27247 417
rect 27281 383 27291 417
rect 27239 369 27291 383
rect 27321 485 27388 497
rect 27321 451 27344 485
rect 27378 451 27388 485
rect 27321 417 27388 451
rect 27321 383 27344 417
rect 27378 383 27388 417
rect 27321 369 27388 383
rect 27102 307 27112 341
rect 27146 307 27158 341
rect 27102 297 27158 307
rect 27336 349 27388 369
rect 27336 315 27344 349
rect 27378 315 27388 349
rect 27336 297 27388 315
rect 27418 449 27470 497
rect 27418 415 27428 449
rect 27462 415 27470 449
rect 27418 381 27470 415
rect 27418 347 27428 381
rect 27462 347 27470 381
rect 27535 477 27587 491
rect 27535 443 27543 477
rect 27577 443 27587 477
rect 27535 409 27587 443
rect 27535 375 27543 409
rect 27577 375 27587 409
rect 27535 363 27587 375
rect 27617 461 27671 491
rect 27617 427 27627 461
rect 27661 427 27671 461
rect 27617 363 27671 427
rect 27701 477 27753 491
rect 27701 443 27711 477
rect 27745 443 27753 477
rect 27701 409 27753 443
rect 27886 485 27938 497
rect 27886 451 27894 485
rect 27928 451 27938 485
rect 27886 413 27938 451
rect 27968 477 28030 497
rect 27968 443 27978 477
rect 28012 443 28030 477
rect 27968 413 28030 443
rect 28060 483 28129 497
rect 28060 449 28071 483
rect 28105 449 28129 483
rect 28060 413 28129 449
rect 28159 459 28269 497
rect 28159 425 28225 459
rect 28259 425 28269 459
rect 28159 413 28269 425
rect 28299 475 28366 497
rect 28299 441 28322 475
rect 28356 441 28366 475
rect 28299 413 28366 441
rect 28396 459 28448 497
rect 28396 425 28406 459
rect 28440 425 28448 459
rect 28396 413 28448 425
rect 28511 485 28563 497
rect 28511 451 28519 485
rect 28553 451 28563 485
rect 27701 375 27711 409
rect 27745 375 27753 409
rect 27701 363 27753 375
rect 27418 297 27470 347
rect 28511 329 28563 451
rect 28593 477 28662 497
rect 28593 443 28607 477
rect 28641 443 28662 477
rect 28593 413 28662 443
rect 28692 484 28748 497
rect 28692 450 28704 484
rect 28738 450 28748 484
rect 28692 413 28748 450
rect 28778 413 28832 497
rect 28862 485 28940 497
rect 28862 451 28896 485
rect 28930 451 28940 485
rect 28862 413 28940 451
rect 28970 459 29024 497
rect 28970 425 28980 459
rect 29014 425 29024 459
rect 28970 413 29024 425
rect 29054 485 29188 497
rect 29054 451 29066 485
rect 29100 451 29144 485
rect 29178 451 29188 485
rect 29054 413 29188 451
rect 28593 329 28647 413
rect 29138 297 29188 413
rect 29218 477 29274 497
rect 29218 443 29228 477
rect 29262 443 29274 477
rect 29218 409 29274 443
rect 29218 375 29228 409
rect 29262 375 29274 409
rect 29218 341 29274 375
rect 29355 485 29407 497
rect 29355 451 29363 485
rect 29397 451 29407 485
rect 29355 417 29407 451
rect 29355 383 29363 417
rect 29397 383 29407 417
rect 29355 369 29407 383
rect 29437 485 29504 497
rect 29437 451 29460 485
rect 29494 451 29504 485
rect 29437 417 29504 451
rect 29437 383 29460 417
rect 29494 383 29504 417
rect 29437 369 29504 383
rect 29218 307 29228 341
rect 29262 307 29274 341
rect 29218 297 29274 307
rect 29452 349 29504 369
rect 29452 315 29460 349
rect 29494 315 29504 349
rect 29452 297 29504 315
rect 29534 449 29586 497
rect 29534 415 29544 449
rect 29578 415 29586 449
rect 29534 381 29586 415
rect 29534 347 29544 381
rect 29578 347 29586 381
rect 29651 477 29703 491
rect 29651 443 29659 477
rect 29693 443 29703 477
rect 29651 409 29703 443
rect 29651 375 29659 409
rect 29693 375 29703 409
rect 29651 363 29703 375
rect 29733 461 29787 491
rect 29733 427 29743 461
rect 29777 427 29787 461
rect 29733 363 29787 427
rect 29817 477 29869 491
rect 29817 443 29827 477
rect 29861 443 29869 477
rect 29817 409 29869 443
rect 30002 485 30054 497
rect 30002 451 30010 485
rect 30044 451 30054 485
rect 30002 413 30054 451
rect 30084 477 30146 497
rect 30084 443 30094 477
rect 30128 443 30146 477
rect 30084 413 30146 443
rect 30176 483 30245 497
rect 30176 449 30187 483
rect 30221 449 30245 483
rect 30176 413 30245 449
rect 30275 459 30385 497
rect 30275 425 30341 459
rect 30375 425 30385 459
rect 30275 413 30385 425
rect 30415 475 30482 497
rect 30415 441 30438 475
rect 30472 441 30482 475
rect 30415 413 30482 441
rect 30512 459 30564 497
rect 30512 425 30522 459
rect 30556 425 30564 459
rect 30512 413 30564 425
rect 30627 485 30679 497
rect 30627 451 30635 485
rect 30669 451 30679 485
rect 29817 375 29827 409
rect 29861 375 29869 409
rect 29817 363 29869 375
rect 29534 297 29586 347
rect 30627 329 30679 451
rect 30709 477 30778 497
rect 30709 443 30723 477
rect 30757 443 30778 477
rect 30709 413 30778 443
rect 30808 484 30864 497
rect 30808 450 30820 484
rect 30854 450 30864 484
rect 30808 413 30864 450
rect 30894 413 30948 497
rect 30978 485 31056 497
rect 30978 451 31012 485
rect 31046 451 31056 485
rect 30978 413 31056 451
rect 31086 459 31140 497
rect 31086 425 31096 459
rect 31130 425 31140 459
rect 31086 413 31140 425
rect 31170 485 31304 497
rect 31170 451 31182 485
rect 31216 451 31260 485
rect 31294 451 31304 485
rect 31170 413 31304 451
rect 30709 329 30763 413
rect 31254 297 31304 413
rect 31334 477 31390 497
rect 31334 443 31344 477
rect 31378 443 31390 477
rect 31334 409 31390 443
rect 31334 375 31344 409
rect 31378 375 31390 409
rect 31334 341 31390 375
rect 31471 485 31523 497
rect 31471 451 31479 485
rect 31513 451 31523 485
rect 31471 417 31523 451
rect 31471 383 31479 417
rect 31513 383 31523 417
rect 31471 369 31523 383
rect 31553 485 31620 497
rect 31553 451 31576 485
rect 31610 451 31620 485
rect 31553 417 31620 451
rect 31553 383 31576 417
rect 31610 383 31620 417
rect 31553 369 31620 383
rect 31334 307 31344 341
rect 31378 307 31390 341
rect 31334 297 31390 307
rect 31568 349 31620 369
rect 31568 315 31576 349
rect 31610 315 31620 349
rect 31568 297 31620 315
rect 31650 449 31702 497
rect 31650 415 31660 449
rect 31694 415 31702 449
rect 31650 381 31702 415
rect 31650 347 31660 381
rect 31694 347 31702 381
rect 31767 477 31819 491
rect 31767 443 31775 477
rect 31809 443 31819 477
rect 31767 409 31819 443
rect 31767 375 31775 409
rect 31809 375 31819 409
rect 31767 363 31819 375
rect 31849 461 31903 491
rect 31849 427 31859 461
rect 31893 427 31903 461
rect 31849 363 31903 427
rect 31933 477 31985 491
rect 31933 443 31943 477
rect 31977 443 31985 477
rect 31933 409 31985 443
rect 32118 485 32170 497
rect 32118 451 32126 485
rect 32160 451 32170 485
rect 32118 413 32170 451
rect 32200 477 32262 497
rect 32200 443 32210 477
rect 32244 443 32262 477
rect 32200 413 32262 443
rect 32292 483 32361 497
rect 32292 449 32303 483
rect 32337 449 32361 483
rect 32292 413 32361 449
rect 32391 459 32501 497
rect 32391 425 32457 459
rect 32491 425 32501 459
rect 32391 413 32501 425
rect 32531 475 32598 497
rect 32531 441 32554 475
rect 32588 441 32598 475
rect 32531 413 32598 441
rect 32628 459 32680 497
rect 32628 425 32638 459
rect 32672 425 32680 459
rect 32628 413 32680 425
rect 32743 485 32795 497
rect 32743 451 32751 485
rect 32785 451 32795 485
rect 31933 375 31943 409
rect 31977 375 31985 409
rect 31933 363 31985 375
rect 31650 297 31702 347
rect 32743 329 32795 451
rect 32825 477 32894 497
rect 32825 443 32839 477
rect 32873 443 32894 477
rect 32825 413 32894 443
rect 32924 484 32980 497
rect 32924 450 32936 484
rect 32970 450 32980 484
rect 32924 413 32980 450
rect 33010 413 33064 497
rect 33094 485 33172 497
rect 33094 451 33128 485
rect 33162 451 33172 485
rect 33094 413 33172 451
rect 33202 459 33256 497
rect 33202 425 33212 459
rect 33246 425 33256 459
rect 33202 413 33256 425
rect 33286 485 33420 497
rect 33286 451 33298 485
rect 33332 451 33376 485
rect 33410 451 33420 485
rect 33286 413 33420 451
rect 32825 329 32879 413
rect 33370 297 33420 413
rect 33450 477 33506 497
rect 33450 443 33460 477
rect 33494 443 33506 477
rect 33450 409 33506 443
rect 33450 375 33460 409
rect 33494 375 33506 409
rect 33450 341 33506 375
rect 33587 485 33639 497
rect 33587 451 33595 485
rect 33629 451 33639 485
rect 33587 417 33639 451
rect 33587 383 33595 417
rect 33629 383 33639 417
rect 33587 369 33639 383
rect 33669 485 33736 497
rect 33669 451 33692 485
rect 33726 451 33736 485
rect 33669 417 33736 451
rect 33669 383 33692 417
rect 33726 383 33736 417
rect 33669 369 33736 383
rect 33450 307 33460 341
rect 33494 307 33506 341
rect 33450 297 33506 307
rect 33684 349 33736 369
rect 33684 315 33692 349
rect 33726 315 33736 349
rect 33684 297 33736 315
rect 33766 449 33818 497
rect 33766 415 33776 449
rect 33810 415 33818 449
rect 33766 381 33818 415
rect 33766 347 33776 381
rect 33810 347 33818 381
rect 33883 477 33935 491
rect 33883 443 33891 477
rect 33925 443 33935 477
rect 33883 409 33935 443
rect 33883 375 33891 409
rect 33925 375 33935 409
rect 33883 363 33935 375
rect 33965 461 34019 491
rect 33965 427 33975 461
rect 34009 427 34019 461
rect 33965 363 34019 427
rect 34049 477 34101 491
rect 34049 443 34059 477
rect 34093 443 34101 477
rect 34049 409 34101 443
rect 34234 485 34286 497
rect 34234 451 34242 485
rect 34276 451 34286 485
rect 34234 413 34286 451
rect 34316 477 34378 497
rect 34316 443 34326 477
rect 34360 443 34378 477
rect 34316 413 34378 443
rect 34408 483 34477 497
rect 34408 449 34419 483
rect 34453 449 34477 483
rect 34408 413 34477 449
rect 34507 459 34617 497
rect 34507 425 34573 459
rect 34607 425 34617 459
rect 34507 413 34617 425
rect 34647 475 34714 497
rect 34647 441 34670 475
rect 34704 441 34714 475
rect 34647 413 34714 441
rect 34744 459 34796 497
rect 34744 425 34754 459
rect 34788 425 34796 459
rect 34744 413 34796 425
rect 34859 485 34911 497
rect 34859 451 34867 485
rect 34901 451 34911 485
rect 34049 375 34059 409
rect 34093 375 34101 409
rect 34049 363 34101 375
rect 33766 297 33818 347
rect 34859 329 34911 451
rect 34941 477 35010 497
rect 34941 443 34955 477
rect 34989 443 35010 477
rect 34941 413 35010 443
rect 35040 484 35096 497
rect 35040 450 35052 484
rect 35086 450 35096 484
rect 35040 413 35096 450
rect 35126 413 35180 497
rect 35210 485 35288 497
rect 35210 451 35244 485
rect 35278 451 35288 485
rect 35210 413 35288 451
rect 35318 459 35372 497
rect 35318 425 35328 459
rect 35362 425 35372 459
rect 35318 413 35372 425
rect 35402 485 35536 497
rect 35402 451 35414 485
rect 35448 451 35492 485
rect 35526 451 35536 485
rect 35402 413 35536 451
rect 34941 329 34995 413
rect 35486 297 35536 413
rect 35566 477 35622 497
rect 35566 443 35576 477
rect 35610 443 35622 477
rect 35566 409 35622 443
rect 35566 375 35576 409
rect 35610 375 35622 409
rect 35566 341 35622 375
rect 35703 485 35755 497
rect 35703 451 35711 485
rect 35745 451 35755 485
rect 35703 417 35755 451
rect 35703 383 35711 417
rect 35745 383 35755 417
rect 35703 369 35755 383
rect 35785 485 35852 497
rect 35785 451 35808 485
rect 35842 451 35852 485
rect 35785 417 35852 451
rect 35785 383 35808 417
rect 35842 383 35852 417
rect 35785 369 35852 383
rect 35566 307 35576 341
rect 35610 307 35622 341
rect 35566 297 35622 307
rect 35800 349 35852 369
rect 35800 315 35808 349
rect 35842 315 35852 349
rect 35800 297 35852 315
rect 35882 449 35934 497
rect 35882 415 35892 449
rect 35926 415 35934 449
rect 35882 381 35934 415
rect 35882 347 35892 381
rect 35926 347 35934 381
rect 35999 477 36051 491
rect 35999 443 36007 477
rect 36041 443 36051 477
rect 35999 409 36051 443
rect 35999 375 36007 409
rect 36041 375 36051 409
rect 35999 363 36051 375
rect 36081 461 36135 491
rect 36081 427 36091 461
rect 36125 427 36135 461
rect 36081 363 36135 427
rect 36165 477 36217 491
rect 36165 443 36175 477
rect 36209 443 36217 477
rect 36165 409 36217 443
rect 36350 485 36402 497
rect 36350 451 36358 485
rect 36392 451 36402 485
rect 36350 413 36402 451
rect 36432 477 36494 497
rect 36432 443 36442 477
rect 36476 443 36494 477
rect 36432 413 36494 443
rect 36524 483 36593 497
rect 36524 449 36535 483
rect 36569 449 36593 483
rect 36524 413 36593 449
rect 36623 459 36733 497
rect 36623 425 36689 459
rect 36723 425 36733 459
rect 36623 413 36733 425
rect 36763 475 36830 497
rect 36763 441 36786 475
rect 36820 441 36830 475
rect 36763 413 36830 441
rect 36860 459 36912 497
rect 36860 425 36870 459
rect 36904 425 36912 459
rect 36860 413 36912 425
rect 36975 485 37027 497
rect 36975 451 36983 485
rect 37017 451 37027 485
rect 36165 375 36175 409
rect 36209 375 36217 409
rect 36165 363 36217 375
rect 35882 297 35934 347
rect 36975 329 37027 451
rect 37057 477 37126 497
rect 37057 443 37071 477
rect 37105 443 37126 477
rect 37057 413 37126 443
rect 37156 484 37212 497
rect 37156 450 37168 484
rect 37202 450 37212 484
rect 37156 413 37212 450
rect 37242 413 37296 497
rect 37326 485 37404 497
rect 37326 451 37360 485
rect 37394 451 37404 485
rect 37326 413 37404 451
rect 37434 459 37488 497
rect 37434 425 37444 459
rect 37478 425 37488 459
rect 37434 413 37488 425
rect 37518 485 37652 497
rect 37518 451 37530 485
rect 37564 451 37608 485
rect 37642 451 37652 485
rect 37518 413 37652 451
rect 37057 329 37111 413
rect 37602 297 37652 413
rect 37682 477 37738 497
rect 37682 443 37692 477
rect 37726 443 37738 477
rect 37682 409 37738 443
rect 37682 375 37692 409
rect 37726 375 37738 409
rect 37682 341 37738 375
rect 37819 485 37871 497
rect 37819 451 37827 485
rect 37861 451 37871 485
rect 37819 417 37871 451
rect 37819 383 37827 417
rect 37861 383 37871 417
rect 37819 369 37871 383
rect 37901 485 37968 497
rect 37901 451 37924 485
rect 37958 451 37968 485
rect 37901 417 37968 451
rect 37901 383 37924 417
rect 37958 383 37968 417
rect 37901 369 37968 383
rect 37682 307 37692 341
rect 37726 307 37738 341
rect 37682 297 37738 307
rect 37916 349 37968 369
rect 37916 315 37924 349
rect 37958 315 37968 349
rect 37916 297 37968 315
rect 37998 449 38050 497
rect 37998 415 38008 449
rect 38042 415 38050 449
rect 37998 381 38050 415
rect 37998 347 38008 381
rect 38042 347 38050 381
rect 38115 477 38167 491
rect 38115 443 38123 477
rect 38157 443 38167 477
rect 38115 409 38167 443
rect 38115 375 38123 409
rect 38157 375 38167 409
rect 38115 363 38167 375
rect 38197 461 38251 491
rect 38197 427 38207 461
rect 38241 427 38251 461
rect 38197 363 38251 427
rect 38281 477 38333 491
rect 38281 443 38291 477
rect 38325 443 38333 477
rect 38281 409 38333 443
rect 38466 485 38518 497
rect 38466 451 38474 485
rect 38508 451 38518 485
rect 38466 413 38518 451
rect 38548 477 38610 497
rect 38548 443 38558 477
rect 38592 443 38610 477
rect 38548 413 38610 443
rect 38640 483 38709 497
rect 38640 449 38651 483
rect 38685 449 38709 483
rect 38640 413 38709 449
rect 38739 459 38849 497
rect 38739 425 38805 459
rect 38839 425 38849 459
rect 38739 413 38849 425
rect 38879 475 38946 497
rect 38879 441 38902 475
rect 38936 441 38946 475
rect 38879 413 38946 441
rect 38976 459 39028 497
rect 38976 425 38986 459
rect 39020 425 39028 459
rect 38976 413 39028 425
rect 39091 485 39143 497
rect 39091 451 39099 485
rect 39133 451 39143 485
rect 38281 375 38291 409
rect 38325 375 38333 409
rect 38281 363 38333 375
rect 37998 297 38050 347
rect 39091 329 39143 451
rect 39173 477 39242 497
rect 39173 443 39187 477
rect 39221 443 39242 477
rect 39173 413 39242 443
rect 39272 484 39328 497
rect 39272 450 39284 484
rect 39318 450 39328 484
rect 39272 413 39328 450
rect 39358 413 39412 497
rect 39442 485 39520 497
rect 39442 451 39476 485
rect 39510 451 39520 485
rect 39442 413 39520 451
rect 39550 459 39604 497
rect 39550 425 39560 459
rect 39594 425 39604 459
rect 39550 413 39604 425
rect 39634 485 39768 497
rect 39634 451 39646 485
rect 39680 451 39724 485
rect 39758 451 39768 485
rect 39634 413 39768 451
rect 39173 329 39227 413
rect 39718 297 39768 413
rect 39798 477 39854 497
rect 39798 443 39808 477
rect 39842 443 39854 477
rect 39798 409 39854 443
rect 39798 375 39808 409
rect 39842 375 39854 409
rect 39798 341 39854 375
rect 39935 485 39987 497
rect 39935 451 39943 485
rect 39977 451 39987 485
rect 39935 417 39987 451
rect 39935 383 39943 417
rect 39977 383 39987 417
rect 39935 369 39987 383
rect 40017 485 40084 497
rect 40017 451 40040 485
rect 40074 451 40084 485
rect 40017 417 40084 451
rect 40017 383 40040 417
rect 40074 383 40084 417
rect 40017 369 40084 383
rect 39798 307 39808 341
rect 39842 307 39854 341
rect 39798 297 39854 307
rect 40032 349 40084 369
rect 40032 315 40040 349
rect 40074 315 40084 349
rect 40032 297 40084 315
rect 40114 449 40166 497
rect 40114 415 40124 449
rect 40158 415 40166 449
rect 40114 381 40166 415
rect 40114 347 40124 381
rect 40158 347 40166 381
rect 40231 477 40283 491
rect 40231 443 40239 477
rect 40273 443 40283 477
rect 40231 409 40283 443
rect 40231 375 40239 409
rect 40273 375 40283 409
rect 40231 363 40283 375
rect 40313 461 40367 491
rect 40313 427 40323 461
rect 40357 427 40367 461
rect 40313 363 40367 427
rect 40397 477 40449 491
rect 40397 443 40407 477
rect 40441 443 40449 477
rect 40397 409 40449 443
rect 40582 485 40634 497
rect 40582 451 40590 485
rect 40624 451 40634 485
rect 40582 413 40634 451
rect 40664 477 40726 497
rect 40664 443 40674 477
rect 40708 443 40726 477
rect 40664 413 40726 443
rect 40756 483 40825 497
rect 40756 449 40767 483
rect 40801 449 40825 483
rect 40756 413 40825 449
rect 40855 459 40965 497
rect 40855 425 40921 459
rect 40955 425 40965 459
rect 40855 413 40965 425
rect 40995 475 41062 497
rect 40995 441 41018 475
rect 41052 441 41062 475
rect 40995 413 41062 441
rect 41092 459 41144 497
rect 41092 425 41102 459
rect 41136 425 41144 459
rect 41092 413 41144 425
rect 41207 485 41259 497
rect 41207 451 41215 485
rect 41249 451 41259 485
rect 40397 375 40407 409
rect 40441 375 40449 409
rect 40397 363 40449 375
rect 40114 297 40166 347
rect 41207 329 41259 451
rect 41289 477 41358 497
rect 41289 443 41303 477
rect 41337 443 41358 477
rect 41289 413 41358 443
rect 41388 484 41444 497
rect 41388 450 41400 484
rect 41434 450 41444 484
rect 41388 413 41444 450
rect 41474 413 41528 497
rect 41558 485 41636 497
rect 41558 451 41592 485
rect 41626 451 41636 485
rect 41558 413 41636 451
rect 41666 459 41720 497
rect 41666 425 41676 459
rect 41710 425 41720 459
rect 41666 413 41720 425
rect 41750 485 41884 497
rect 41750 451 41762 485
rect 41796 451 41840 485
rect 41874 451 41884 485
rect 41750 413 41884 451
rect 41289 329 41343 413
rect 41834 297 41884 413
rect 41914 477 41970 497
rect 41914 443 41924 477
rect 41958 443 41970 477
rect 41914 409 41970 443
rect 41914 375 41924 409
rect 41958 375 41970 409
rect 41914 341 41970 375
rect 42051 485 42103 497
rect 42051 451 42059 485
rect 42093 451 42103 485
rect 42051 417 42103 451
rect 42051 383 42059 417
rect 42093 383 42103 417
rect 42051 369 42103 383
rect 42133 485 42200 497
rect 42133 451 42156 485
rect 42190 451 42200 485
rect 42133 417 42200 451
rect 42133 383 42156 417
rect 42190 383 42200 417
rect 42133 369 42200 383
rect 41914 307 41924 341
rect 41958 307 41970 341
rect 41914 297 41970 307
rect 42148 349 42200 369
rect 42148 315 42156 349
rect 42190 315 42200 349
rect 42148 297 42200 315
rect 42230 449 42282 497
rect 42230 415 42240 449
rect 42274 415 42282 449
rect 42230 381 42282 415
rect 42230 347 42240 381
rect 42274 347 42282 381
rect 42230 297 42282 347
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 325 55 359 89
rect 458 61 492 95
rect 565 61 599 95
rect 911 59 945 93
rect 1023 55 1057 89
rect 1133 59 1167 93
rect 1345 55 1379 89
rect 1563 75 1597 109
rect 1667 98 1701 132
rect 1751 131 1785 165
rect 1751 63 1785 97
rect 1855 85 1889 119
rect 1952 79 1986 113
rect 2036 109 2070 143
rect 2151 85 2185 119
rect 2235 59 2269 93
rect 2319 85 2353 119
rect 2441 55 2475 89
rect 2574 61 2608 95
rect 2681 61 2715 95
rect 3027 59 3061 93
rect 3139 55 3173 89
rect 3249 59 3283 93
rect 3461 55 3495 89
rect 3679 75 3713 109
rect 3783 98 3817 132
rect 3867 131 3901 165
rect 3867 63 3901 97
rect 3971 85 4005 119
rect 4068 79 4102 113
rect 4152 109 4186 143
rect 4267 85 4301 119
rect 4351 59 4385 93
rect 4435 85 4469 119
rect 4557 55 4591 89
rect 4690 61 4724 95
rect 4797 61 4831 95
rect 5143 59 5177 93
rect 5255 55 5289 89
rect 5365 59 5399 93
rect 5577 55 5611 89
rect 5795 75 5829 109
rect 5899 98 5933 132
rect 5983 131 6017 165
rect 5983 63 6017 97
rect 6087 85 6121 119
rect 6184 79 6218 113
rect 6268 109 6302 143
rect 6383 85 6417 119
rect 6467 59 6501 93
rect 6551 85 6585 119
rect 6673 55 6707 89
rect 6806 61 6840 95
rect 6913 61 6947 95
rect 7259 59 7293 93
rect 7371 55 7405 89
rect 7481 59 7515 93
rect 7693 55 7727 89
rect 7911 75 7945 109
rect 8015 98 8049 132
rect 8099 131 8133 165
rect 8099 63 8133 97
rect 8203 85 8237 119
rect 8300 79 8334 113
rect 8384 109 8418 143
rect 8499 85 8533 119
rect 8583 59 8617 93
rect 8667 85 8701 119
rect 8789 55 8823 89
rect 8922 61 8956 95
rect 9029 61 9063 95
rect 9375 59 9409 93
rect 9487 55 9521 89
rect 9597 59 9631 93
rect 9809 55 9843 89
rect 10027 75 10061 109
rect 10131 98 10165 132
rect 10215 131 10249 165
rect 10215 63 10249 97
rect 10319 85 10353 119
rect 10416 79 10450 113
rect 10500 109 10534 143
rect 10615 85 10649 119
rect 10699 59 10733 93
rect 10783 85 10817 119
rect 10905 55 10939 89
rect 11038 61 11072 95
rect 11145 61 11179 95
rect 11491 59 11525 93
rect 11603 55 11637 89
rect 11713 59 11747 93
rect 11925 55 11959 89
rect 12143 75 12177 109
rect 12247 98 12281 132
rect 12331 131 12365 165
rect 12331 63 12365 97
rect 12435 85 12469 119
rect 12532 79 12566 113
rect 12616 109 12650 143
rect 12731 85 12765 119
rect 12815 59 12849 93
rect 12899 85 12933 119
rect 13021 55 13055 89
rect 13154 61 13188 95
rect 13261 61 13295 95
rect 13607 59 13641 93
rect 13719 55 13753 89
rect 13829 59 13863 93
rect 14041 55 14075 89
rect 14259 75 14293 109
rect 14363 98 14397 132
rect 14447 131 14481 165
rect 14447 63 14481 97
rect 14551 85 14585 119
rect 14648 79 14682 113
rect 14732 109 14766 143
rect 14847 85 14881 119
rect 14931 59 14965 93
rect 15015 85 15049 119
rect 15137 55 15171 89
rect 15270 61 15304 95
rect 15377 61 15411 95
rect 15723 59 15757 93
rect 15835 55 15869 89
rect 15945 59 15979 93
rect 16157 55 16191 89
rect 16375 75 16409 109
rect 16479 98 16513 132
rect 16563 131 16597 165
rect 16563 63 16597 97
rect 16667 85 16701 119
rect 16764 79 16798 113
rect 16848 109 16882 143
rect 16963 85 16997 119
rect 17047 59 17081 93
rect 17131 85 17165 119
rect 17253 55 17287 89
rect 17386 61 17420 95
rect 17493 61 17527 95
rect 17839 59 17873 93
rect 17951 55 17985 89
rect 18061 59 18095 93
rect 18273 55 18307 89
rect 18491 75 18525 109
rect 18595 98 18629 132
rect 18679 131 18713 165
rect 18679 63 18713 97
rect 18783 85 18817 119
rect 18880 79 18914 113
rect 18964 109 18998 143
rect 19079 85 19113 119
rect 19163 59 19197 93
rect 19247 85 19281 119
rect 19369 55 19403 89
rect 19502 61 19536 95
rect 19609 61 19643 95
rect 19955 59 19989 93
rect 20067 55 20101 89
rect 20177 59 20211 93
rect 20389 55 20423 89
rect 20607 75 20641 109
rect 20711 98 20745 132
rect 20795 131 20829 165
rect 20795 63 20829 97
rect 20899 85 20933 119
rect 20996 79 21030 113
rect 21080 109 21114 143
rect 21195 85 21229 119
rect 21279 59 21313 93
rect 21363 85 21397 119
rect 21485 55 21519 89
rect 21618 61 21652 95
rect 21725 61 21759 95
rect 22071 59 22105 93
rect 22183 55 22217 89
rect 22293 59 22327 93
rect 22505 55 22539 89
rect 22723 75 22757 109
rect 22827 98 22861 132
rect 22911 131 22945 165
rect 22911 63 22945 97
rect 23015 85 23049 119
rect 23112 79 23146 113
rect 23196 109 23230 143
rect 23311 85 23345 119
rect 23395 59 23429 93
rect 23479 85 23513 119
rect 23601 55 23635 89
rect 23734 61 23768 95
rect 23841 61 23875 95
rect 24187 59 24221 93
rect 24299 55 24333 89
rect 24409 59 24443 93
rect 24621 55 24655 89
rect 24839 75 24873 109
rect 24943 98 24977 132
rect 25027 131 25061 165
rect 25027 63 25061 97
rect 25131 85 25165 119
rect 25228 79 25262 113
rect 25312 109 25346 143
rect 25427 85 25461 119
rect 25511 59 25545 93
rect 25595 85 25629 119
rect 25717 55 25751 89
rect 25850 61 25884 95
rect 25957 61 25991 95
rect 26303 59 26337 93
rect 26415 55 26449 89
rect 26525 59 26559 93
rect 26737 55 26771 89
rect 26955 75 26989 109
rect 27059 98 27093 132
rect 27143 131 27177 165
rect 27143 63 27177 97
rect 27247 85 27281 119
rect 27344 79 27378 113
rect 27428 109 27462 143
rect 27543 85 27577 119
rect 27627 59 27661 93
rect 27711 85 27745 119
rect 27833 55 27867 89
rect 27966 61 28000 95
rect 28073 61 28107 95
rect 28419 59 28453 93
rect 28531 55 28565 89
rect 28641 59 28675 93
rect 28853 55 28887 89
rect 29071 75 29105 109
rect 29175 98 29209 132
rect 29259 131 29293 165
rect 29259 63 29293 97
rect 29363 85 29397 119
rect 29460 79 29494 113
rect 29544 109 29578 143
rect 29659 85 29693 119
rect 29743 59 29777 93
rect 29827 85 29861 119
rect 29949 55 29983 89
rect 30082 61 30116 95
rect 30189 61 30223 95
rect 30535 59 30569 93
rect 30647 55 30681 89
rect 30757 59 30791 93
rect 30969 55 31003 89
rect 31187 75 31221 109
rect 31291 98 31325 132
rect 31375 131 31409 165
rect 31375 63 31409 97
rect 31479 85 31513 119
rect 31576 79 31610 113
rect 31660 109 31694 143
rect 31775 85 31809 119
rect 31859 59 31893 93
rect 31943 85 31977 119
rect 32065 55 32099 89
rect 32198 61 32232 95
rect 32305 61 32339 95
rect 32651 59 32685 93
rect 32763 55 32797 89
rect 32873 59 32907 93
rect 33085 55 33119 89
rect 33303 75 33337 109
rect 33407 98 33441 132
rect 33491 131 33525 165
rect 33491 63 33525 97
rect 33595 85 33629 119
rect 33692 79 33726 113
rect 33776 109 33810 143
rect 33891 85 33925 119
rect 33975 59 34009 93
rect 34059 85 34093 119
rect 34181 55 34215 89
rect 34314 61 34348 95
rect 34421 61 34455 95
rect 34767 59 34801 93
rect 34879 55 34913 89
rect 34989 59 35023 93
rect 35201 55 35235 89
rect 35419 75 35453 109
rect 35523 98 35557 132
rect 35607 131 35641 165
rect 35607 63 35641 97
rect 35711 85 35745 119
rect 35808 79 35842 113
rect 35892 109 35926 143
rect 36007 85 36041 119
rect 36091 59 36125 93
rect 36175 85 36209 119
rect 36297 55 36331 89
rect 36430 61 36464 95
rect 36537 61 36571 95
rect 36883 59 36917 93
rect 36995 55 37029 89
rect 37105 59 37139 93
rect 37317 55 37351 89
rect 37535 75 37569 109
rect 37639 98 37673 132
rect 37723 131 37757 165
rect 37723 63 37757 97
rect 37827 85 37861 119
rect 37924 79 37958 113
rect 38008 109 38042 143
rect 38123 85 38157 119
rect 38207 59 38241 93
rect 38291 85 38325 119
rect 38413 55 38447 89
rect 38546 61 38580 95
rect 38653 61 38687 95
rect 38999 59 39033 93
rect 39111 55 39145 89
rect 39221 59 39255 93
rect 39433 55 39467 89
rect 39651 75 39685 109
rect 39755 98 39789 132
rect 39839 131 39873 165
rect 39839 63 39873 97
rect 39943 85 39977 119
rect 40040 79 40074 113
rect 40124 109 40158 143
rect 40239 85 40273 119
rect 40323 59 40357 93
rect 40407 85 40441 119
rect 40529 55 40563 89
rect 40662 61 40696 95
rect 40769 61 40803 95
rect 41115 59 41149 93
rect 41227 55 41261 89
rect 41337 59 41371 93
rect 41549 55 41583 89
rect 41767 75 41801 109
rect 41871 98 41905 132
rect 41955 131 41989 165
rect 41955 63 41989 97
rect 42059 85 42093 119
rect 42156 79 42190 113
rect 42240 109 42274 143
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 386 451 420 485
rect 470 443 504 477
rect 563 449 597 483
rect 717 425 751 459
rect 814 441 848 475
rect 898 425 932 459
rect 1011 451 1045 485
rect 203 375 237 409
rect 1099 443 1133 477
rect 1196 450 1230 484
rect 1388 451 1422 485
rect 1472 425 1506 459
rect 1558 451 1592 485
rect 1636 451 1670 485
rect 1720 443 1754 477
rect 1720 375 1754 409
rect 1855 451 1889 485
rect 1855 383 1889 417
rect 1952 451 1986 485
rect 1952 383 1986 417
rect 1720 307 1754 341
rect 1952 315 1986 349
rect 2036 415 2070 449
rect 2036 347 2070 381
rect 2151 443 2185 477
rect 2151 375 2185 409
rect 2235 427 2269 461
rect 2319 443 2353 477
rect 2502 451 2536 485
rect 2586 443 2620 477
rect 2679 449 2713 483
rect 2833 425 2867 459
rect 2930 441 2964 475
rect 3014 425 3048 459
rect 3127 451 3161 485
rect 2319 375 2353 409
rect 3215 443 3249 477
rect 3312 450 3346 484
rect 3504 451 3538 485
rect 3588 425 3622 459
rect 3674 451 3708 485
rect 3752 451 3786 485
rect 3836 443 3870 477
rect 3836 375 3870 409
rect 3971 451 4005 485
rect 3971 383 4005 417
rect 4068 451 4102 485
rect 4068 383 4102 417
rect 3836 307 3870 341
rect 4068 315 4102 349
rect 4152 415 4186 449
rect 4152 347 4186 381
rect 4267 443 4301 477
rect 4267 375 4301 409
rect 4351 427 4385 461
rect 4435 443 4469 477
rect 4618 451 4652 485
rect 4702 443 4736 477
rect 4795 449 4829 483
rect 4949 425 4983 459
rect 5046 441 5080 475
rect 5130 425 5164 459
rect 5243 451 5277 485
rect 4435 375 4469 409
rect 5331 443 5365 477
rect 5428 450 5462 484
rect 5620 451 5654 485
rect 5704 425 5738 459
rect 5790 451 5824 485
rect 5868 451 5902 485
rect 5952 443 5986 477
rect 5952 375 5986 409
rect 6087 451 6121 485
rect 6087 383 6121 417
rect 6184 451 6218 485
rect 6184 383 6218 417
rect 5952 307 5986 341
rect 6184 315 6218 349
rect 6268 415 6302 449
rect 6268 347 6302 381
rect 6383 443 6417 477
rect 6383 375 6417 409
rect 6467 427 6501 461
rect 6551 443 6585 477
rect 6734 451 6768 485
rect 6818 443 6852 477
rect 6911 449 6945 483
rect 7065 425 7099 459
rect 7162 441 7196 475
rect 7246 425 7280 459
rect 7359 451 7393 485
rect 6551 375 6585 409
rect 7447 443 7481 477
rect 7544 450 7578 484
rect 7736 451 7770 485
rect 7820 425 7854 459
rect 7906 451 7940 485
rect 7984 451 8018 485
rect 8068 443 8102 477
rect 8068 375 8102 409
rect 8203 451 8237 485
rect 8203 383 8237 417
rect 8300 451 8334 485
rect 8300 383 8334 417
rect 8068 307 8102 341
rect 8300 315 8334 349
rect 8384 415 8418 449
rect 8384 347 8418 381
rect 8499 443 8533 477
rect 8499 375 8533 409
rect 8583 427 8617 461
rect 8667 443 8701 477
rect 8850 451 8884 485
rect 8934 443 8968 477
rect 9027 449 9061 483
rect 9181 425 9215 459
rect 9278 441 9312 475
rect 9362 425 9396 459
rect 9475 451 9509 485
rect 8667 375 8701 409
rect 9563 443 9597 477
rect 9660 450 9694 484
rect 9852 451 9886 485
rect 9936 425 9970 459
rect 10022 451 10056 485
rect 10100 451 10134 485
rect 10184 443 10218 477
rect 10184 375 10218 409
rect 10319 451 10353 485
rect 10319 383 10353 417
rect 10416 451 10450 485
rect 10416 383 10450 417
rect 10184 307 10218 341
rect 10416 315 10450 349
rect 10500 415 10534 449
rect 10500 347 10534 381
rect 10615 443 10649 477
rect 10615 375 10649 409
rect 10699 427 10733 461
rect 10783 443 10817 477
rect 10966 451 11000 485
rect 11050 443 11084 477
rect 11143 449 11177 483
rect 11297 425 11331 459
rect 11394 441 11428 475
rect 11478 425 11512 459
rect 11591 451 11625 485
rect 10783 375 10817 409
rect 11679 443 11713 477
rect 11776 450 11810 484
rect 11968 451 12002 485
rect 12052 425 12086 459
rect 12138 451 12172 485
rect 12216 451 12250 485
rect 12300 443 12334 477
rect 12300 375 12334 409
rect 12435 451 12469 485
rect 12435 383 12469 417
rect 12532 451 12566 485
rect 12532 383 12566 417
rect 12300 307 12334 341
rect 12532 315 12566 349
rect 12616 415 12650 449
rect 12616 347 12650 381
rect 12731 443 12765 477
rect 12731 375 12765 409
rect 12815 427 12849 461
rect 12899 443 12933 477
rect 13082 451 13116 485
rect 13166 443 13200 477
rect 13259 449 13293 483
rect 13413 425 13447 459
rect 13510 441 13544 475
rect 13594 425 13628 459
rect 13707 451 13741 485
rect 12899 375 12933 409
rect 13795 443 13829 477
rect 13892 450 13926 484
rect 14084 451 14118 485
rect 14168 425 14202 459
rect 14254 451 14288 485
rect 14332 451 14366 485
rect 14416 443 14450 477
rect 14416 375 14450 409
rect 14551 451 14585 485
rect 14551 383 14585 417
rect 14648 451 14682 485
rect 14648 383 14682 417
rect 14416 307 14450 341
rect 14648 315 14682 349
rect 14732 415 14766 449
rect 14732 347 14766 381
rect 14847 443 14881 477
rect 14847 375 14881 409
rect 14931 427 14965 461
rect 15015 443 15049 477
rect 15198 451 15232 485
rect 15282 443 15316 477
rect 15375 449 15409 483
rect 15529 425 15563 459
rect 15626 441 15660 475
rect 15710 425 15744 459
rect 15823 451 15857 485
rect 15015 375 15049 409
rect 15911 443 15945 477
rect 16008 450 16042 484
rect 16200 451 16234 485
rect 16284 425 16318 459
rect 16370 451 16404 485
rect 16448 451 16482 485
rect 16532 443 16566 477
rect 16532 375 16566 409
rect 16667 451 16701 485
rect 16667 383 16701 417
rect 16764 451 16798 485
rect 16764 383 16798 417
rect 16532 307 16566 341
rect 16764 315 16798 349
rect 16848 415 16882 449
rect 16848 347 16882 381
rect 16963 443 16997 477
rect 16963 375 16997 409
rect 17047 427 17081 461
rect 17131 443 17165 477
rect 17314 451 17348 485
rect 17398 443 17432 477
rect 17491 449 17525 483
rect 17645 425 17679 459
rect 17742 441 17776 475
rect 17826 425 17860 459
rect 17939 451 17973 485
rect 17131 375 17165 409
rect 18027 443 18061 477
rect 18124 450 18158 484
rect 18316 451 18350 485
rect 18400 425 18434 459
rect 18486 451 18520 485
rect 18564 451 18598 485
rect 18648 443 18682 477
rect 18648 375 18682 409
rect 18783 451 18817 485
rect 18783 383 18817 417
rect 18880 451 18914 485
rect 18880 383 18914 417
rect 18648 307 18682 341
rect 18880 315 18914 349
rect 18964 415 18998 449
rect 18964 347 18998 381
rect 19079 443 19113 477
rect 19079 375 19113 409
rect 19163 427 19197 461
rect 19247 443 19281 477
rect 19430 451 19464 485
rect 19514 443 19548 477
rect 19607 449 19641 483
rect 19761 425 19795 459
rect 19858 441 19892 475
rect 19942 425 19976 459
rect 20055 451 20089 485
rect 19247 375 19281 409
rect 20143 443 20177 477
rect 20240 450 20274 484
rect 20432 451 20466 485
rect 20516 425 20550 459
rect 20602 451 20636 485
rect 20680 451 20714 485
rect 20764 443 20798 477
rect 20764 375 20798 409
rect 20899 451 20933 485
rect 20899 383 20933 417
rect 20996 451 21030 485
rect 20996 383 21030 417
rect 20764 307 20798 341
rect 20996 315 21030 349
rect 21080 415 21114 449
rect 21080 347 21114 381
rect 21195 443 21229 477
rect 21195 375 21229 409
rect 21279 427 21313 461
rect 21363 443 21397 477
rect 21546 451 21580 485
rect 21630 443 21664 477
rect 21723 449 21757 483
rect 21877 425 21911 459
rect 21974 441 22008 475
rect 22058 425 22092 459
rect 22171 451 22205 485
rect 21363 375 21397 409
rect 22259 443 22293 477
rect 22356 450 22390 484
rect 22548 451 22582 485
rect 22632 425 22666 459
rect 22718 451 22752 485
rect 22796 451 22830 485
rect 22880 443 22914 477
rect 22880 375 22914 409
rect 23015 451 23049 485
rect 23015 383 23049 417
rect 23112 451 23146 485
rect 23112 383 23146 417
rect 22880 307 22914 341
rect 23112 315 23146 349
rect 23196 415 23230 449
rect 23196 347 23230 381
rect 23311 443 23345 477
rect 23311 375 23345 409
rect 23395 427 23429 461
rect 23479 443 23513 477
rect 23662 451 23696 485
rect 23746 443 23780 477
rect 23839 449 23873 483
rect 23993 425 24027 459
rect 24090 441 24124 475
rect 24174 425 24208 459
rect 24287 451 24321 485
rect 23479 375 23513 409
rect 24375 443 24409 477
rect 24472 450 24506 484
rect 24664 451 24698 485
rect 24748 425 24782 459
rect 24834 451 24868 485
rect 24912 451 24946 485
rect 24996 443 25030 477
rect 24996 375 25030 409
rect 25131 451 25165 485
rect 25131 383 25165 417
rect 25228 451 25262 485
rect 25228 383 25262 417
rect 24996 307 25030 341
rect 25228 315 25262 349
rect 25312 415 25346 449
rect 25312 347 25346 381
rect 25427 443 25461 477
rect 25427 375 25461 409
rect 25511 427 25545 461
rect 25595 443 25629 477
rect 25778 451 25812 485
rect 25862 443 25896 477
rect 25955 449 25989 483
rect 26109 425 26143 459
rect 26206 441 26240 475
rect 26290 425 26324 459
rect 26403 451 26437 485
rect 25595 375 25629 409
rect 26491 443 26525 477
rect 26588 450 26622 484
rect 26780 451 26814 485
rect 26864 425 26898 459
rect 26950 451 26984 485
rect 27028 451 27062 485
rect 27112 443 27146 477
rect 27112 375 27146 409
rect 27247 451 27281 485
rect 27247 383 27281 417
rect 27344 451 27378 485
rect 27344 383 27378 417
rect 27112 307 27146 341
rect 27344 315 27378 349
rect 27428 415 27462 449
rect 27428 347 27462 381
rect 27543 443 27577 477
rect 27543 375 27577 409
rect 27627 427 27661 461
rect 27711 443 27745 477
rect 27894 451 27928 485
rect 27978 443 28012 477
rect 28071 449 28105 483
rect 28225 425 28259 459
rect 28322 441 28356 475
rect 28406 425 28440 459
rect 28519 451 28553 485
rect 27711 375 27745 409
rect 28607 443 28641 477
rect 28704 450 28738 484
rect 28896 451 28930 485
rect 28980 425 29014 459
rect 29066 451 29100 485
rect 29144 451 29178 485
rect 29228 443 29262 477
rect 29228 375 29262 409
rect 29363 451 29397 485
rect 29363 383 29397 417
rect 29460 451 29494 485
rect 29460 383 29494 417
rect 29228 307 29262 341
rect 29460 315 29494 349
rect 29544 415 29578 449
rect 29544 347 29578 381
rect 29659 443 29693 477
rect 29659 375 29693 409
rect 29743 427 29777 461
rect 29827 443 29861 477
rect 30010 451 30044 485
rect 30094 443 30128 477
rect 30187 449 30221 483
rect 30341 425 30375 459
rect 30438 441 30472 475
rect 30522 425 30556 459
rect 30635 451 30669 485
rect 29827 375 29861 409
rect 30723 443 30757 477
rect 30820 450 30854 484
rect 31012 451 31046 485
rect 31096 425 31130 459
rect 31182 451 31216 485
rect 31260 451 31294 485
rect 31344 443 31378 477
rect 31344 375 31378 409
rect 31479 451 31513 485
rect 31479 383 31513 417
rect 31576 451 31610 485
rect 31576 383 31610 417
rect 31344 307 31378 341
rect 31576 315 31610 349
rect 31660 415 31694 449
rect 31660 347 31694 381
rect 31775 443 31809 477
rect 31775 375 31809 409
rect 31859 427 31893 461
rect 31943 443 31977 477
rect 32126 451 32160 485
rect 32210 443 32244 477
rect 32303 449 32337 483
rect 32457 425 32491 459
rect 32554 441 32588 475
rect 32638 425 32672 459
rect 32751 451 32785 485
rect 31943 375 31977 409
rect 32839 443 32873 477
rect 32936 450 32970 484
rect 33128 451 33162 485
rect 33212 425 33246 459
rect 33298 451 33332 485
rect 33376 451 33410 485
rect 33460 443 33494 477
rect 33460 375 33494 409
rect 33595 451 33629 485
rect 33595 383 33629 417
rect 33692 451 33726 485
rect 33692 383 33726 417
rect 33460 307 33494 341
rect 33692 315 33726 349
rect 33776 415 33810 449
rect 33776 347 33810 381
rect 33891 443 33925 477
rect 33891 375 33925 409
rect 33975 427 34009 461
rect 34059 443 34093 477
rect 34242 451 34276 485
rect 34326 443 34360 477
rect 34419 449 34453 483
rect 34573 425 34607 459
rect 34670 441 34704 475
rect 34754 425 34788 459
rect 34867 451 34901 485
rect 34059 375 34093 409
rect 34955 443 34989 477
rect 35052 450 35086 484
rect 35244 451 35278 485
rect 35328 425 35362 459
rect 35414 451 35448 485
rect 35492 451 35526 485
rect 35576 443 35610 477
rect 35576 375 35610 409
rect 35711 451 35745 485
rect 35711 383 35745 417
rect 35808 451 35842 485
rect 35808 383 35842 417
rect 35576 307 35610 341
rect 35808 315 35842 349
rect 35892 415 35926 449
rect 35892 347 35926 381
rect 36007 443 36041 477
rect 36007 375 36041 409
rect 36091 427 36125 461
rect 36175 443 36209 477
rect 36358 451 36392 485
rect 36442 443 36476 477
rect 36535 449 36569 483
rect 36689 425 36723 459
rect 36786 441 36820 475
rect 36870 425 36904 459
rect 36983 451 37017 485
rect 36175 375 36209 409
rect 37071 443 37105 477
rect 37168 450 37202 484
rect 37360 451 37394 485
rect 37444 425 37478 459
rect 37530 451 37564 485
rect 37608 451 37642 485
rect 37692 443 37726 477
rect 37692 375 37726 409
rect 37827 451 37861 485
rect 37827 383 37861 417
rect 37924 451 37958 485
rect 37924 383 37958 417
rect 37692 307 37726 341
rect 37924 315 37958 349
rect 38008 415 38042 449
rect 38008 347 38042 381
rect 38123 443 38157 477
rect 38123 375 38157 409
rect 38207 427 38241 461
rect 38291 443 38325 477
rect 38474 451 38508 485
rect 38558 443 38592 477
rect 38651 449 38685 483
rect 38805 425 38839 459
rect 38902 441 38936 475
rect 38986 425 39020 459
rect 39099 451 39133 485
rect 38291 375 38325 409
rect 39187 443 39221 477
rect 39284 450 39318 484
rect 39476 451 39510 485
rect 39560 425 39594 459
rect 39646 451 39680 485
rect 39724 451 39758 485
rect 39808 443 39842 477
rect 39808 375 39842 409
rect 39943 451 39977 485
rect 39943 383 39977 417
rect 40040 451 40074 485
rect 40040 383 40074 417
rect 39808 307 39842 341
rect 40040 315 40074 349
rect 40124 415 40158 449
rect 40124 347 40158 381
rect 40239 443 40273 477
rect 40239 375 40273 409
rect 40323 427 40357 461
rect 40407 443 40441 477
rect 40590 451 40624 485
rect 40674 443 40708 477
rect 40767 449 40801 483
rect 40921 425 40955 459
rect 41018 441 41052 475
rect 41102 425 41136 459
rect 41215 451 41249 485
rect 40407 375 40441 409
rect 41303 443 41337 477
rect 41400 450 41434 484
rect 41592 451 41626 485
rect 41676 425 41710 459
rect 41762 451 41796 485
rect 41840 451 41874 485
rect 41924 443 41958 477
rect 41924 375 41958 409
rect 42059 451 42093 485
rect 42059 383 42093 417
rect 42156 451 42190 485
rect 42156 383 42190 417
rect 41924 307 41958 341
rect 42156 315 42190 349
rect 42240 415 42274 449
rect 42240 347 42274 381
<< psubdiff >>
rect 0 -41 29 -7
rect 63 -41 121 -7
rect 155 -41 213 -7
rect 247 -41 305 -7
rect 339 -41 397 -7
rect 431 -41 489 -7
rect 523 -41 581 -7
rect 615 -41 673 -7
rect 707 -41 765 -7
rect 799 -41 857 -7
rect 891 -41 949 -7
rect 983 -41 1041 -7
rect 1075 -41 1133 -7
rect 1167 -41 1225 -7
rect 1259 -41 1317 -7
rect 1351 -41 1409 -7
rect 1443 -41 1501 -7
rect 1535 -41 1593 -7
rect 1627 -41 1685 -7
rect 1719 -41 1777 -7
rect 1811 -41 1869 -7
rect 1903 -41 1961 -7
rect 1995 -41 2053 -7
rect 2087 -41 2145 -7
rect 2179 -41 2237 -7
rect 2271 -41 2329 -7
rect 2363 -41 2421 -7
rect 2455 -41 2513 -7
rect 2547 -41 2605 -7
rect 2639 -41 2697 -7
rect 2731 -41 2789 -7
rect 2823 -41 2881 -7
rect 2915 -41 2973 -7
rect 3007 -41 3065 -7
rect 3099 -41 3157 -7
rect 3191 -41 3249 -7
rect 3283 -41 3341 -7
rect 3375 -41 3433 -7
rect 3467 -41 3525 -7
rect 3559 -41 3617 -7
rect 3651 -41 3709 -7
rect 3743 -41 3801 -7
rect 3835 -41 3893 -7
rect 3927 -41 3985 -7
rect 4019 -41 4077 -7
rect 4111 -41 4169 -7
rect 4203 -41 4261 -7
rect 4295 -41 4353 -7
rect 4387 -41 4445 -7
rect 4479 -41 4537 -7
rect 4571 -41 4629 -7
rect 4663 -41 4721 -7
rect 4755 -41 4813 -7
rect 4847 -41 4905 -7
rect 4939 -41 4997 -7
rect 5031 -41 5089 -7
rect 5123 -41 5181 -7
rect 5215 -41 5273 -7
rect 5307 -41 5365 -7
rect 5399 -41 5457 -7
rect 5491 -41 5549 -7
rect 5583 -41 5641 -7
rect 5675 -41 5733 -7
rect 5767 -41 5825 -7
rect 5859 -41 5917 -7
rect 5951 -41 6009 -7
rect 6043 -41 6101 -7
rect 6135 -41 6193 -7
rect 6227 -41 6285 -7
rect 6319 -41 6377 -7
rect 6411 -41 6469 -7
rect 6503 -41 6561 -7
rect 6595 -41 6653 -7
rect 6687 -41 6745 -7
rect 6779 -41 6837 -7
rect 6871 -41 6929 -7
rect 6963 -41 7021 -7
rect 7055 -41 7113 -7
rect 7147 -41 7205 -7
rect 7239 -41 7297 -7
rect 7331 -41 7389 -7
rect 7423 -41 7481 -7
rect 7515 -41 7573 -7
rect 7607 -41 7665 -7
rect 7699 -41 7757 -7
rect 7791 -41 7849 -7
rect 7883 -41 7941 -7
rect 7975 -41 8033 -7
rect 8067 -41 8125 -7
rect 8159 -41 8217 -7
rect 8251 -41 8309 -7
rect 8343 -41 8401 -7
rect 8435 -41 8493 -7
rect 8527 -41 8585 -7
rect 8619 -41 8677 -7
rect 8711 -41 8769 -7
rect 8803 -41 8861 -7
rect 8895 -41 8953 -7
rect 8987 -41 9045 -7
rect 9079 -41 9137 -7
rect 9171 -41 9229 -7
rect 9263 -41 9321 -7
rect 9355 -41 9413 -7
rect 9447 -41 9505 -7
rect 9539 -41 9597 -7
rect 9631 -41 9689 -7
rect 9723 -41 9781 -7
rect 9815 -41 9873 -7
rect 9907 -41 9965 -7
rect 9999 -41 10057 -7
rect 10091 -41 10149 -7
rect 10183 -41 10241 -7
rect 10275 -41 10333 -7
rect 10367 -41 10425 -7
rect 10459 -41 10517 -7
rect 10551 -41 10609 -7
rect 10643 -41 10701 -7
rect 10735 -41 10793 -7
rect 10827 -41 10885 -7
rect 10919 -41 10977 -7
rect 11011 -41 11069 -7
rect 11103 -41 11161 -7
rect 11195 -41 11253 -7
rect 11287 -41 11345 -7
rect 11379 -41 11437 -7
rect 11471 -41 11529 -7
rect 11563 -41 11621 -7
rect 11655 -41 11713 -7
rect 11747 -41 11805 -7
rect 11839 -41 11897 -7
rect 11931 -41 11989 -7
rect 12023 -41 12081 -7
rect 12115 -41 12173 -7
rect 12207 -41 12265 -7
rect 12299 -41 12357 -7
rect 12391 -41 12449 -7
rect 12483 -41 12541 -7
rect 12575 -41 12633 -7
rect 12667 -41 12725 -7
rect 12759 -41 12817 -7
rect 12851 -41 12909 -7
rect 12943 -41 13001 -7
rect 13035 -41 13093 -7
rect 13127 -41 13185 -7
rect 13219 -41 13277 -7
rect 13311 -41 13369 -7
rect 13403 -41 13461 -7
rect 13495 -41 13553 -7
rect 13587 -41 13645 -7
rect 13679 -41 13737 -7
rect 13771 -41 13829 -7
rect 13863 -41 13921 -7
rect 13955 -41 14013 -7
rect 14047 -41 14105 -7
rect 14139 -41 14197 -7
rect 14231 -41 14289 -7
rect 14323 -41 14381 -7
rect 14415 -41 14473 -7
rect 14507 -41 14565 -7
rect 14599 -41 14657 -7
rect 14691 -41 14749 -7
rect 14783 -41 14841 -7
rect 14875 -41 14933 -7
rect 14967 -41 15025 -7
rect 15059 -41 15117 -7
rect 15151 -41 15209 -7
rect 15243 -41 15301 -7
rect 15335 -41 15393 -7
rect 15427 -41 15485 -7
rect 15519 -41 15577 -7
rect 15611 -41 15669 -7
rect 15703 -41 15761 -7
rect 15795 -41 15853 -7
rect 15887 -41 15945 -7
rect 15979 -41 16037 -7
rect 16071 -41 16129 -7
rect 16163 -41 16221 -7
rect 16255 -41 16313 -7
rect 16347 -41 16405 -7
rect 16439 -41 16497 -7
rect 16531 -41 16589 -7
rect 16623 -41 16681 -7
rect 16715 -41 16773 -7
rect 16807 -41 16865 -7
rect 16899 -41 16957 -7
rect 16991 -41 17049 -7
rect 17083 -41 17141 -7
rect 17175 -41 17233 -7
rect 17267 -41 17325 -7
rect 17359 -41 17417 -7
rect 17451 -41 17509 -7
rect 17543 -41 17601 -7
rect 17635 -41 17693 -7
rect 17727 -41 17785 -7
rect 17819 -41 17877 -7
rect 17911 -41 17969 -7
rect 18003 -41 18061 -7
rect 18095 -41 18153 -7
rect 18187 -41 18245 -7
rect 18279 -41 18337 -7
rect 18371 -41 18429 -7
rect 18463 -41 18521 -7
rect 18555 -41 18613 -7
rect 18647 -41 18705 -7
rect 18739 -41 18797 -7
rect 18831 -41 18889 -7
rect 18923 -41 18981 -7
rect 19015 -41 19073 -7
rect 19107 -41 19165 -7
rect 19199 -41 19257 -7
rect 19291 -41 19349 -7
rect 19383 -41 19441 -7
rect 19475 -41 19533 -7
rect 19567 -41 19625 -7
rect 19659 -41 19717 -7
rect 19751 -41 19809 -7
rect 19843 -41 19901 -7
rect 19935 -41 19993 -7
rect 20027 -41 20085 -7
rect 20119 -41 20177 -7
rect 20211 -41 20269 -7
rect 20303 -41 20361 -7
rect 20395 -41 20453 -7
rect 20487 -41 20545 -7
rect 20579 -41 20637 -7
rect 20671 -41 20729 -7
rect 20763 -41 20821 -7
rect 20855 -41 20913 -7
rect 20947 -41 21005 -7
rect 21039 -41 21097 -7
rect 21131 -41 21189 -7
rect 21223 -41 21281 -7
rect 21315 -41 21373 -7
rect 21407 -41 21465 -7
rect 21499 -41 21557 -7
rect 21591 -41 21649 -7
rect 21683 -41 21741 -7
rect 21775 -41 21833 -7
rect 21867 -41 21925 -7
rect 21959 -41 22017 -7
rect 22051 -41 22109 -7
rect 22143 -41 22201 -7
rect 22235 -41 22293 -7
rect 22327 -41 22385 -7
rect 22419 -41 22477 -7
rect 22511 -41 22569 -7
rect 22603 -41 22661 -7
rect 22695 -41 22753 -7
rect 22787 -41 22845 -7
rect 22879 -41 22937 -7
rect 22971 -41 23029 -7
rect 23063 -41 23121 -7
rect 23155 -41 23213 -7
rect 23247 -41 23305 -7
rect 23339 -41 23397 -7
rect 23431 -41 23489 -7
rect 23523 -41 23581 -7
rect 23615 -41 23673 -7
rect 23707 -41 23765 -7
rect 23799 -41 23857 -7
rect 23891 -41 23949 -7
rect 23983 -41 24041 -7
rect 24075 -41 24133 -7
rect 24167 -41 24225 -7
rect 24259 -41 24317 -7
rect 24351 -41 24409 -7
rect 24443 -41 24501 -7
rect 24535 -41 24593 -7
rect 24627 -41 24685 -7
rect 24719 -41 24777 -7
rect 24811 -41 24869 -7
rect 24903 -41 24961 -7
rect 24995 -41 25053 -7
rect 25087 -41 25145 -7
rect 25179 -41 25237 -7
rect 25271 -41 25329 -7
rect 25363 -41 25421 -7
rect 25455 -41 25513 -7
rect 25547 -41 25605 -7
rect 25639 -41 25697 -7
rect 25731 -41 25789 -7
rect 25823 -41 25881 -7
rect 25915 -41 25973 -7
rect 26007 -41 26065 -7
rect 26099 -41 26157 -7
rect 26191 -41 26249 -7
rect 26283 -41 26341 -7
rect 26375 -41 26433 -7
rect 26467 -41 26525 -7
rect 26559 -41 26617 -7
rect 26651 -41 26709 -7
rect 26743 -41 26801 -7
rect 26835 -41 26893 -7
rect 26927 -41 26985 -7
rect 27019 -41 27077 -7
rect 27111 -41 27169 -7
rect 27203 -41 27261 -7
rect 27295 -41 27353 -7
rect 27387 -41 27445 -7
rect 27479 -41 27537 -7
rect 27571 -41 27629 -7
rect 27663 -41 27721 -7
rect 27755 -41 27813 -7
rect 27847 -41 27905 -7
rect 27939 -41 27997 -7
rect 28031 -41 28089 -7
rect 28123 -41 28181 -7
rect 28215 -41 28273 -7
rect 28307 -41 28365 -7
rect 28399 -41 28457 -7
rect 28491 -41 28549 -7
rect 28583 -41 28641 -7
rect 28675 -41 28733 -7
rect 28767 -41 28825 -7
rect 28859 -41 28917 -7
rect 28951 -41 29009 -7
rect 29043 -41 29101 -7
rect 29135 -41 29193 -7
rect 29227 -41 29285 -7
rect 29319 -41 29377 -7
rect 29411 -41 29469 -7
rect 29503 -41 29561 -7
rect 29595 -41 29653 -7
rect 29687 -41 29745 -7
rect 29779 -41 29837 -7
rect 29871 -41 29929 -7
rect 29963 -41 30021 -7
rect 30055 -41 30113 -7
rect 30147 -41 30205 -7
rect 30239 -41 30297 -7
rect 30331 -41 30389 -7
rect 30423 -41 30481 -7
rect 30515 -41 30573 -7
rect 30607 -41 30665 -7
rect 30699 -41 30757 -7
rect 30791 -41 30849 -7
rect 30883 -41 30941 -7
rect 30975 -41 31033 -7
rect 31067 -41 31125 -7
rect 31159 -41 31217 -7
rect 31251 -41 31309 -7
rect 31343 -41 31401 -7
rect 31435 -41 31493 -7
rect 31527 -41 31585 -7
rect 31619 -41 31677 -7
rect 31711 -41 31769 -7
rect 31803 -41 31861 -7
rect 31895 -41 31953 -7
rect 31987 -41 32045 -7
rect 32079 -41 32137 -7
rect 32171 -41 32229 -7
rect 32263 -41 32321 -7
rect 32355 -41 32413 -7
rect 32447 -41 32505 -7
rect 32539 -41 32597 -7
rect 32631 -41 32689 -7
rect 32723 -41 32781 -7
rect 32815 -41 32873 -7
rect 32907 -41 32965 -7
rect 32999 -41 33057 -7
rect 33091 -41 33149 -7
rect 33183 -41 33241 -7
rect 33275 -41 33333 -7
rect 33367 -41 33425 -7
rect 33459 -41 33517 -7
rect 33551 -41 33609 -7
rect 33643 -41 33701 -7
rect 33735 -41 33793 -7
rect 33827 -41 33885 -7
rect 33919 -41 33977 -7
rect 34011 -41 34069 -7
rect 34103 -41 34161 -7
rect 34195 -41 34253 -7
rect 34287 -41 34345 -7
rect 34379 -41 34437 -7
rect 34471 -41 34529 -7
rect 34563 -41 34621 -7
rect 34655 -41 34713 -7
rect 34747 -41 34805 -7
rect 34839 -41 34897 -7
rect 34931 -41 34989 -7
rect 35023 -41 35081 -7
rect 35115 -41 35173 -7
rect 35207 -41 35265 -7
rect 35299 -41 35357 -7
rect 35391 -41 35449 -7
rect 35483 -41 35541 -7
rect 35575 -41 35633 -7
rect 35667 -41 35725 -7
rect 35759 -41 35817 -7
rect 35851 -41 35909 -7
rect 35943 -41 36001 -7
rect 36035 -41 36093 -7
rect 36127 -41 36185 -7
rect 36219 -41 36277 -7
rect 36311 -41 36369 -7
rect 36403 -41 36461 -7
rect 36495 -41 36553 -7
rect 36587 -41 36645 -7
rect 36679 -41 36737 -7
rect 36771 -41 36829 -7
rect 36863 -41 36921 -7
rect 36955 -41 37013 -7
rect 37047 -41 37105 -7
rect 37139 -41 37197 -7
rect 37231 -41 37289 -7
rect 37323 -41 37381 -7
rect 37415 -41 37473 -7
rect 37507 -41 37565 -7
rect 37599 -41 37657 -7
rect 37691 -41 37749 -7
rect 37783 -41 37841 -7
rect 37875 -41 37933 -7
rect 37967 -41 38025 -7
rect 38059 -41 38117 -7
rect 38151 -41 38209 -7
rect 38243 -41 38301 -7
rect 38335 -41 38393 -7
rect 38427 -41 38485 -7
rect 38519 -41 38577 -7
rect 38611 -41 38669 -7
rect 38703 -41 38761 -7
rect 38795 -41 38853 -7
rect 38887 -41 38945 -7
rect 38979 -41 39037 -7
rect 39071 -41 39129 -7
rect 39163 -41 39221 -7
rect 39255 -41 39313 -7
rect 39347 -41 39405 -7
rect 39439 -41 39497 -7
rect 39531 -41 39589 -7
rect 39623 -41 39681 -7
rect 39715 -41 39773 -7
rect 39807 -41 39865 -7
rect 39899 -41 39957 -7
rect 39991 -41 40049 -7
rect 40083 -41 40141 -7
rect 40175 -41 40233 -7
rect 40267 -41 40325 -7
rect 40359 -41 40417 -7
rect 40451 -41 40509 -7
rect 40543 -41 40601 -7
rect 40635 -41 40693 -7
rect 40727 -41 40785 -7
rect 40819 -41 40877 -7
rect 40911 -41 40969 -7
rect 41003 -41 41061 -7
rect 41095 -41 41153 -7
rect 41187 -41 41245 -7
rect 41279 -41 41337 -7
rect 41371 -41 41429 -7
rect 41463 -41 41521 -7
rect 41555 -41 41613 -7
rect 41647 -41 41705 -7
rect 41739 -41 41797 -7
rect 41831 -41 41889 -7
rect 41923 -41 41981 -7
rect 42015 -41 42073 -7
rect 42107 -41 42165 -7
rect 42199 -41 42257 -7
rect 42291 -41 42320 -7
<< nsubdiff >>
rect 0 551 29 585
rect 63 551 121 585
rect 155 551 213 585
rect 247 551 305 585
rect 339 551 397 585
rect 431 551 489 585
rect 523 551 581 585
rect 615 551 673 585
rect 707 551 765 585
rect 799 551 857 585
rect 891 551 949 585
rect 983 551 1041 585
rect 1075 551 1133 585
rect 1167 551 1225 585
rect 1259 551 1317 585
rect 1351 551 1409 585
rect 1443 551 1501 585
rect 1535 551 1593 585
rect 1627 551 1685 585
rect 1719 551 1777 585
rect 1811 551 1869 585
rect 1903 551 1961 585
rect 1995 551 2053 585
rect 2087 551 2145 585
rect 2179 551 2237 585
rect 2271 551 2329 585
rect 2363 551 2421 585
rect 2455 551 2513 585
rect 2547 551 2605 585
rect 2639 551 2697 585
rect 2731 551 2789 585
rect 2823 551 2881 585
rect 2915 551 2973 585
rect 3007 551 3065 585
rect 3099 551 3157 585
rect 3191 551 3249 585
rect 3283 551 3341 585
rect 3375 551 3433 585
rect 3467 551 3525 585
rect 3559 551 3617 585
rect 3651 551 3709 585
rect 3743 551 3801 585
rect 3835 551 3893 585
rect 3927 551 3985 585
rect 4019 551 4077 585
rect 4111 551 4169 585
rect 4203 551 4261 585
rect 4295 551 4353 585
rect 4387 551 4445 585
rect 4479 551 4537 585
rect 4571 551 4629 585
rect 4663 551 4721 585
rect 4755 551 4813 585
rect 4847 551 4905 585
rect 4939 551 4997 585
rect 5031 551 5089 585
rect 5123 551 5181 585
rect 5215 551 5273 585
rect 5307 551 5365 585
rect 5399 551 5457 585
rect 5491 551 5549 585
rect 5583 551 5641 585
rect 5675 551 5733 585
rect 5767 551 5825 585
rect 5859 551 5917 585
rect 5951 551 6009 585
rect 6043 551 6101 585
rect 6135 551 6193 585
rect 6227 551 6285 585
rect 6319 551 6377 585
rect 6411 551 6469 585
rect 6503 551 6561 585
rect 6595 551 6653 585
rect 6687 551 6745 585
rect 6779 551 6837 585
rect 6871 551 6929 585
rect 6963 551 7021 585
rect 7055 551 7113 585
rect 7147 551 7205 585
rect 7239 551 7297 585
rect 7331 551 7389 585
rect 7423 551 7481 585
rect 7515 551 7573 585
rect 7607 551 7665 585
rect 7699 551 7757 585
rect 7791 551 7849 585
rect 7883 551 7941 585
rect 7975 551 8033 585
rect 8067 551 8125 585
rect 8159 551 8217 585
rect 8251 551 8309 585
rect 8343 551 8401 585
rect 8435 551 8493 585
rect 8527 551 8585 585
rect 8619 551 8677 585
rect 8711 551 8769 585
rect 8803 551 8861 585
rect 8895 551 8953 585
rect 8987 551 9045 585
rect 9079 551 9137 585
rect 9171 551 9229 585
rect 9263 551 9321 585
rect 9355 551 9413 585
rect 9447 551 9505 585
rect 9539 551 9597 585
rect 9631 551 9689 585
rect 9723 551 9781 585
rect 9815 551 9873 585
rect 9907 551 9965 585
rect 9999 551 10057 585
rect 10091 551 10149 585
rect 10183 551 10241 585
rect 10275 551 10333 585
rect 10367 551 10425 585
rect 10459 551 10517 585
rect 10551 551 10609 585
rect 10643 551 10701 585
rect 10735 551 10793 585
rect 10827 551 10885 585
rect 10919 551 10977 585
rect 11011 551 11069 585
rect 11103 551 11161 585
rect 11195 551 11253 585
rect 11287 551 11345 585
rect 11379 551 11437 585
rect 11471 551 11529 585
rect 11563 551 11621 585
rect 11655 551 11713 585
rect 11747 551 11805 585
rect 11839 551 11897 585
rect 11931 551 11989 585
rect 12023 551 12081 585
rect 12115 551 12173 585
rect 12207 551 12265 585
rect 12299 551 12357 585
rect 12391 551 12449 585
rect 12483 551 12541 585
rect 12575 551 12633 585
rect 12667 551 12725 585
rect 12759 551 12817 585
rect 12851 551 12909 585
rect 12943 551 13001 585
rect 13035 551 13093 585
rect 13127 551 13185 585
rect 13219 551 13277 585
rect 13311 551 13369 585
rect 13403 551 13461 585
rect 13495 551 13553 585
rect 13587 551 13645 585
rect 13679 551 13737 585
rect 13771 551 13829 585
rect 13863 551 13921 585
rect 13955 551 14013 585
rect 14047 551 14105 585
rect 14139 551 14197 585
rect 14231 551 14289 585
rect 14323 551 14381 585
rect 14415 551 14473 585
rect 14507 551 14565 585
rect 14599 551 14657 585
rect 14691 551 14749 585
rect 14783 551 14841 585
rect 14875 551 14933 585
rect 14967 551 15025 585
rect 15059 551 15117 585
rect 15151 551 15209 585
rect 15243 551 15301 585
rect 15335 551 15393 585
rect 15427 551 15485 585
rect 15519 551 15577 585
rect 15611 551 15669 585
rect 15703 551 15761 585
rect 15795 551 15853 585
rect 15887 551 15945 585
rect 15979 551 16037 585
rect 16071 551 16129 585
rect 16163 551 16221 585
rect 16255 551 16313 585
rect 16347 551 16405 585
rect 16439 551 16497 585
rect 16531 551 16589 585
rect 16623 551 16681 585
rect 16715 551 16773 585
rect 16807 551 16865 585
rect 16899 551 16957 585
rect 16991 551 17049 585
rect 17083 551 17141 585
rect 17175 551 17233 585
rect 17267 551 17325 585
rect 17359 551 17417 585
rect 17451 551 17509 585
rect 17543 551 17601 585
rect 17635 551 17693 585
rect 17727 551 17785 585
rect 17819 551 17877 585
rect 17911 551 17969 585
rect 18003 551 18061 585
rect 18095 551 18153 585
rect 18187 551 18245 585
rect 18279 551 18337 585
rect 18371 551 18429 585
rect 18463 551 18521 585
rect 18555 551 18613 585
rect 18647 551 18705 585
rect 18739 551 18797 585
rect 18831 551 18889 585
rect 18923 551 18981 585
rect 19015 551 19073 585
rect 19107 551 19165 585
rect 19199 551 19257 585
rect 19291 551 19349 585
rect 19383 551 19441 585
rect 19475 551 19533 585
rect 19567 551 19625 585
rect 19659 551 19717 585
rect 19751 551 19809 585
rect 19843 551 19901 585
rect 19935 551 19993 585
rect 20027 551 20085 585
rect 20119 551 20177 585
rect 20211 551 20269 585
rect 20303 551 20361 585
rect 20395 551 20453 585
rect 20487 551 20545 585
rect 20579 551 20637 585
rect 20671 551 20729 585
rect 20763 551 20821 585
rect 20855 551 20913 585
rect 20947 551 21005 585
rect 21039 551 21097 585
rect 21131 551 21189 585
rect 21223 551 21281 585
rect 21315 551 21373 585
rect 21407 551 21465 585
rect 21499 551 21557 585
rect 21591 551 21649 585
rect 21683 551 21741 585
rect 21775 551 21833 585
rect 21867 551 21925 585
rect 21959 551 22017 585
rect 22051 551 22109 585
rect 22143 551 22201 585
rect 22235 551 22293 585
rect 22327 551 22385 585
rect 22419 551 22477 585
rect 22511 551 22569 585
rect 22603 551 22661 585
rect 22695 551 22753 585
rect 22787 551 22845 585
rect 22879 551 22937 585
rect 22971 551 23029 585
rect 23063 551 23121 585
rect 23155 551 23213 585
rect 23247 551 23305 585
rect 23339 551 23397 585
rect 23431 551 23489 585
rect 23523 551 23581 585
rect 23615 551 23673 585
rect 23707 551 23765 585
rect 23799 551 23857 585
rect 23891 551 23949 585
rect 23983 551 24041 585
rect 24075 551 24133 585
rect 24167 551 24225 585
rect 24259 551 24317 585
rect 24351 551 24409 585
rect 24443 551 24501 585
rect 24535 551 24593 585
rect 24627 551 24685 585
rect 24719 551 24777 585
rect 24811 551 24869 585
rect 24903 551 24961 585
rect 24995 551 25053 585
rect 25087 551 25145 585
rect 25179 551 25237 585
rect 25271 551 25329 585
rect 25363 551 25421 585
rect 25455 551 25513 585
rect 25547 551 25605 585
rect 25639 551 25697 585
rect 25731 551 25789 585
rect 25823 551 25881 585
rect 25915 551 25973 585
rect 26007 551 26065 585
rect 26099 551 26157 585
rect 26191 551 26249 585
rect 26283 551 26341 585
rect 26375 551 26433 585
rect 26467 551 26525 585
rect 26559 551 26617 585
rect 26651 551 26709 585
rect 26743 551 26801 585
rect 26835 551 26893 585
rect 26927 551 26985 585
rect 27019 551 27077 585
rect 27111 551 27169 585
rect 27203 551 27261 585
rect 27295 551 27353 585
rect 27387 551 27445 585
rect 27479 551 27537 585
rect 27571 551 27629 585
rect 27663 551 27721 585
rect 27755 551 27813 585
rect 27847 551 27905 585
rect 27939 551 27997 585
rect 28031 551 28089 585
rect 28123 551 28181 585
rect 28215 551 28273 585
rect 28307 551 28365 585
rect 28399 551 28457 585
rect 28491 551 28549 585
rect 28583 551 28641 585
rect 28675 551 28733 585
rect 28767 551 28825 585
rect 28859 551 28917 585
rect 28951 551 29009 585
rect 29043 551 29101 585
rect 29135 551 29193 585
rect 29227 551 29285 585
rect 29319 551 29377 585
rect 29411 551 29469 585
rect 29503 551 29561 585
rect 29595 551 29653 585
rect 29687 551 29745 585
rect 29779 551 29837 585
rect 29871 551 29929 585
rect 29963 551 30021 585
rect 30055 551 30113 585
rect 30147 551 30205 585
rect 30239 551 30297 585
rect 30331 551 30389 585
rect 30423 551 30481 585
rect 30515 551 30573 585
rect 30607 551 30665 585
rect 30699 551 30757 585
rect 30791 551 30849 585
rect 30883 551 30941 585
rect 30975 551 31033 585
rect 31067 551 31125 585
rect 31159 551 31217 585
rect 31251 551 31309 585
rect 31343 551 31401 585
rect 31435 551 31493 585
rect 31527 551 31585 585
rect 31619 551 31677 585
rect 31711 551 31769 585
rect 31803 551 31861 585
rect 31895 551 31953 585
rect 31987 551 32045 585
rect 32079 551 32137 585
rect 32171 551 32229 585
rect 32263 551 32321 585
rect 32355 551 32413 585
rect 32447 551 32505 585
rect 32539 551 32597 585
rect 32631 551 32689 585
rect 32723 551 32781 585
rect 32815 551 32873 585
rect 32907 551 32965 585
rect 32999 551 33057 585
rect 33091 551 33149 585
rect 33183 551 33241 585
rect 33275 551 33333 585
rect 33367 551 33425 585
rect 33459 551 33517 585
rect 33551 551 33609 585
rect 33643 551 33701 585
rect 33735 551 33793 585
rect 33827 551 33885 585
rect 33919 551 33977 585
rect 34011 551 34069 585
rect 34103 551 34161 585
rect 34195 551 34253 585
rect 34287 551 34345 585
rect 34379 551 34437 585
rect 34471 551 34529 585
rect 34563 551 34621 585
rect 34655 551 34713 585
rect 34747 551 34805 585
rect 34839 551 34897 585
rect 34931 551 34989 585
rect 35023 551 35081 585
rect 35115 551 35173 585
rect 35207 551 35265 585
rect 35299 551 35357 585
rect 35391 551 35449 585
rect 35483 551 35541 585
rect 35575 551 35633 585
rect 35667 551 35725 585
rect 35759 551 35817 585
rect 35851 551 35909 585
rect 35943 551 36001 585
rect 36035 551 36093 585
rect 36127 551 36185 585
rect 36219 551 36277 585
rect 36311 551 36369 585
rect 36403 551 36461 585
rect 36495 551 36553 585
rect 36587 551 36645 585
rect 36679 551 36737 585
rect 36771 551 36829 585
rect 36863 551 36921 585
rect 36955 551 37013 585
rect 37047 551 37105 585
rect 37139 551 37197 585
rect 37231 551 37289 585
rect 37323 551 37381 585
rect 37415 551 37473 585
rect 37507 551 37565 585
rect 37599 551 37657 585
rect 37691 551 37749 585
rect 37783 551 37841 585
rect 37875 551 37933 585
rect 37967 551 38025 585
rect 38059 551 38117 585
rect 38151 551 38209 585
rect 38243 551 38301 585
rect 38335 551 38393 585
rect 38427 551 38485 585
rect 38519 551 38577 585
rect 38611 551 38669 585
rect 38703 551 38761 585
rect 38795 551 38853 585
rect 38887 551 38945 585
rect 38979 551 39037 585
rect 39071 551 39129 585
rect 39163 551 39221 585
rect 39255 551 39313 585
rect 39347 551 39405 585
rect 39439 551 39497 585
rect 39531 551 39589 585
rect 39623 551 39681 585
rect 39715 551 39773 585
rect 39807 551 39865 585
rect 39899 551 39957 585
rect 39991 551 40049 585
rect 40083 551 40141 585
rect 40175 551 40233 585
rect 40267 551 40325 585
rect 40359 551 40417 585
rect 40451 551 40509 585
rect 40543 551 40601 585
rect 40635 551 40693 585
rect 40727 551 40785 585
rect 40819 551 40877 585
rect 40911 551 40969 585
rect 41003 551 41061 585
rect 41095 551 41153 585
rect 41187 551 41245 585
rect 41279 551 41337 585
rect 41371 551 41429 585
rect 41463 551 41521 585
rect 41555 551 41613 585
rect 41647 551 41705 585
rect 41739 551 41797 585
rect 41831 551 41889 585
rect 41923 551 41981 585
rect 42015 551 42073 585
rect 42107 551 42165 585
rect 42199 551 42257 585
rect 42291 551 42320 585
<< psubdiffcont >>
rect 29 -41 63 -7
rect 121 -41 155 -7
rect 213 -41 247 -7
rect 305 -41 339 -7
rect 397 -41 431 -7
rect 489 -41 523 -7
rect 581 -41 615 -7
rect 673 -41 707 -7
rect 765 -41 799 -7
rect 857 -41 891 -7
rect 949 -41 983 -7
rect 1041 -41 1075 -7
rect 1133 -41 1167 -7
rect 1225 -41 1259 -7
rect 1317 -41 1351 -7
rect 1409 -41 1443 -7
rect 1501 -41 1535 -7
rect 1593 -41 1627 -7
rect 1685 -41 1719 -7
rect 1777 -41 1811 -7
rect 1869 -41 1903 -7
rect 1961 -41 1995 -7
rect 2053 -41 2087 -7
rect 2145 -41 2179 -7
rect 2237 -41 2271 -7
rect 2329 -41 2363 -7
rect 2421 -41 2455 -7
rect 2513 -41 2547 -7
rect 2605 -41 2639 -7
rect 2697 -41 2731 -7
rect 2789 -41 2823 -7
rect 2881 -41 2915 -7
rect 2973 -41 3007 -7
rect 3065 -41 3099 -7
rect 3157 -41 3191 -7
rect 3249 -41 3283 -7
rect 3341 -41 3375 -7
rect 3433 -41 3467 -7
rect 3525 -41 3559 -7
rect 3617 -41 3651 -7
rect 3709 -41 3743 -7
rect 3801 -41 3835 -7
rect 3893 -41 3927 -7
rect 3985 -41 4019 -7
rect 4077 -41 4111 -7
rect 4169 -41 4203 -7
rect 4261 -41 4295 -7
rect 4353 -41 4387 -7
rect 4445 -41 4479 -7
rect 4537 -41 4571 -7
rect 4629 -41 4663 -7
rect 4721 -41 4755 -7
rect 4813 -41 4847 -7
rect 4905 -41 4939 -7
rect 4997 -41 5031 -7
rect 5089 -41 5123 -7
rect 5181 -41 5215 -7
rect 5273 -41 5307 -7
rect 5365 -41 5399 -7
rect 5457 -41 5491 -7
rect 5549 -41 5583 -7
rect 5641 -41 5675 -7
rect 5733 -41 5767 -7
rect 5825 -41 5859 -7
rect 5917 -41 5951 -7
rect 6009 -41 6043 -7
rect 6101 -41 6135 -7
rect 6193 -41 6227 -7
rect 6285 -41 6319 -7
rect 6377 -41 6411 -7
rect 6469 -41 6503 -7
rect 6561 -41 6595 -7
rect 6653 -41 6687 -7
rect 6745 -41 6779 -7
rect 6837 -41 6871 -7
rect 6929 -41 6963 -7
rect 7021 -41 7055 -7
rect 7113 -41 7147 -7
rect 7205 -41 7239 -7
rect 7297 -41 7331 -7
rect 7389 -41 7423 -7
rect 7481 -41 7515 -7
rect 7573 -41 7607 -7
rect 7665 -41 7699 -7
rect 7757 -41 7791 -7
rect 7849 -41 7883 -7
rect 7941 -41 7975 -7
rect 8033 -41 8067 -7
rect 8125 -41 8159 -7
rect 8217 -41 8251 -7
rect 8309 -41 8343 -7
rect 8401 -41 8435 -7
rect 8493 -41 8527 -7
rect 8585 -41 8619 -7
rect 8677 -41 8711 -7
rect 8769 -41 8803 -7
rect 8861 -41 8895 -7
rect 8953 -41 8987 -7
rect 9045 -41 9079 -7
rect 9137 -41 9171 -7
rect 9229 -41 9263 -7
rect 9321 -41 9355 -7
rect 9413 -41 9447 -7
rect 9505 -41 9539 -7
rect 9597 -41 9631 -7
rect 9689 -41 9723 -7
rect 9781 -41 9815 -7
rect 9873 -41 9907 -7
rect 9965 -41 9999 -7
rect 10057 -41 10091 -7
rect 10149 -41 10183 -7
rect 10241 -41 10275 -7
rect 10333 -41 10367 -7
rect 10425 -41 10459 -7
rect 10517 -41 10551 -7
rect 10609 -41 10643 -7
rect 10701 -41 10735 -7
rect 10793 -41 10827 -7
rect 10885 -41 10919 -7
rect 10977 -41 11011 -7
rect 11069 -41 11103 -7
rect 11161 -41 11195 -7
rect 11253 -41 11287 -7
rect 11345 -41 11379 -7
rect 11437 -41 11471 -7
rect 11529 -41 11563 -7
rect 11621 -41 11655 -7
rect 11713 -41 11747 -7
rect 11805 -41 11839 -7
rect 11897 -41 11931 -7
rect 11989 -41 12023 -7
rect 12081 -41 12115 -7
rect 12173 -41 12207 -7
rect 12265 -41 12299 -7
rect 12357 -41 12391 -7
rect 12449 -41 12483 -7
rect 12541 -41 12575 -7
rect 12633 -41 12667 -7
rect 12725 -41 12759 -7
rect 12817 -41 12851 -7
rect 12909 -41 12943 -7
rect 13001 -41 13035 -7
rect 13093 -41 13127 -7
rect 13185 -41 13219 -7
rect 13277 -41 13311 -7
rect 13369 -41 13403 -7
rect 13461 -41 13495 -7
rect 13553 -41 13587 -7
rect 13645 -41 13679 -7
rect 13737 -41 13771 -7
rect 13829 -41 13863 -7
rect 13921 -41 13955 -7
rect 14013 -41 14047 -7
rect 14105 -41 14139 -7
rect 14197 -41 14231 -7
rect 14289 -41 14323 -7
rect 14381 -41 14415 -7
rect 14473 -41 14507 -7
rect 14565 -41 14599 -7
rect 14657 -41 14691 -7
rect 14749 -41 14783 -7
rect 14841 -41 14875 -7
rect 14933 -41 14967 -7
rect 15025 -41 15059 -7
rect 15117 -41 15151 -7
rect 15209 -41 15243 -7
rect 15301 -41 15335 -7
rect 15393 -41 15427 -7
rect 15485 -41 15519 -7
rect 15577 -41 15611 -7
rect 15669 -41 15703 -7
rect 15761 -41 15795 -7
rect 15853 -41 15887 -7
rect 15945 -41 15979 -7
rect 16037 -41 16071 -7
rect 16129 -41 16163 -7
rect 16221 -41 16255 -7
rect 16313 -41 16347 -7
rect 16405 -41 16439 -7
rect 16497 -41 16531 -7
rect 16589 -41 16623 -7
rect 16681 -41 16715 -7
rect 16773 -41 16807 -7
rect 16865 -41 16899 -7
rect 16957 -41 16991 -7
rect 17049 -41 17083 -7
rect 17141 -41 17175 -7
rect 17233 -41 17267 -7
rect 17325 -41 17359 -7
rect 17417 -41 17451 -7
rect 17509 -41 17543 -7
rect 17601 -41 17635 -7
rect 17693 -41 17727 -7
rect 17785 -41 17819 -7
rect 17877 -41 17911 -7
rect 17969 -41 18003 -7
rect 18061 -41 18095 -7
rect 18153 -41 18187 -7
rect 18245 -41 18279 -7
rect 18337 -41 18371 -7
rect 18429 -41 18463 -7
rect 18521 -41 18555 -7
rect 18613 -41 18647 -7
rect 18705 -41 18739 -7
rect 18797 -41 18831 -7
rect 18889 -41 18923 -7
rect 18981 -41 19015 -7
rect 19073 -41 19107 -7
rect 19165 -41 19199 -7
rect 19257 -41 19291 -7
rect 19349 -41 19383 -7
rect 19441 -41 19475 -7
rect 19533 -41 19567 -7
rect 19625 -41 19659 -7
rect 19717 -41 19751 -7
rect 19809 -41 19843 -7
rect 19901 -41 19935 -7
rect 19993 -41 20027 -7
rect 20085 -41 20119 -7
rect 20177 -41 20211 -7
rect 20269 -41 20303 -7
rect 20361 -41 20395 -7
rect 20453 -41 20487 -7
rect 20545 -41 20579 -7
rect 20637 -41 20671 -7
rect 20729 -41 20763 -7
rect 20821 -41 20855 -7
rect 20913 -41 20947 -7
rect 21005 -41 21039 -7
rect 21097 -41 21131 -7
rect 21189 -41 21223 -7
rect 21281 -41 21315 -7
rect 21373 -41 21407 -7
rect 21465 -41 21499 -7
rect 21557 -41 21591 -7
rect 21649 -41 21683 -7
rect 21741 -41 21775 -7
rect 21833 -41 21867 -7
rect 21925 -41 21959 -7
rect 22017 -41 22051 -7
rect 22109 -41 22143 -7
rect 22201 -41 22235 -7
rect 22293 -41 22327 -7
rect 22385 -41 22419 -7
rect 22477 -41 22511 -7
rect 22569 -41 22603 -7
rect 22661 -41 22695 -7
rect 22753 -41 22787 -7
rect 22845 -41 22879 -7
rect 22937 -41 22971 -7
rect 23029 -41 23063 -7
rect 23121 -41 23155 -7
rect 23213 -41 23247 -7
rect 23305 -41 23339 -7
rect 23397 -41 23431 -7
rect 23489 -41 23523 -7
rect 23581 -41 23615 -7
rect 23673 -41 23707 -7
rect 23765 -41 23799 -7
rect 23857 -41 23891 -7
rect 23949 -41 23983 -7
rect 24041 -41 24075 -7
rect 24133 -41 24167 -7
rect 24225 -41 24259 -7
rect 24317 -41 24351 -7
rect 24409 -41 24443 -7
rect 24501 -41 24535 -7
rect 24593 -41 24627 -7
rect 24685 -41 24719 -7
rect 24777 -41 24811 -7
rect 24869 -41 24903 -7
rect 24961 -41 24995 -7
rect 25053 -41 25087 -7
rect 25145 -41 25179 -7
rect 25237 -41 25271 -7
rect 25329 -41 25363 -7
rect 25421 -41 25455 -7
rect 25513 -41 25547 -7
rect 25605 -41 25639 -7
rect 25697 -41 25731 -7
rect 25789 -41 25823 -7
rect 25881 -41 25915 -7
rect 25973 -41 26007 -7
rect 26065 -41 26099 -7
rect 26157 -41 26191 -7
rect 26249 -41 26283 -7
rect 26341 -41 26375 -7
rect 26433 -41 26467 -7
rect 26525 -41 26559 -7
rect 26617 -41 26651 -7
rect 26709 -41 26743 -7
rect 26801 -41 26835 -7
rect 26893 -41 26927 -7
rect 26985 -41 27019 -7
rect 27077 -41 27111 -7
rect 27169 -41 27203 -7
rect 27261 -41 27295 -7
rect 27353 -41 27387 -7
rect 27445 -41 27479 -7
rect 27537 -41 27571 -7
rect 27629 -41 27663 -7
rect 27721 -41 27755 -7
rect 27813 -41 27847 -7
rect 27905 -41 27939 -7
rect 27997 -41 28031 -7
rect 28089 -41 28123 -7
rect 28181 -41 28215 -7
rect 28273 -41 28307 -7
rect 28365 -41 28399 -7
rect 28457 -41 28491 -7
rect 28549 -41 28583 -7
rect 28641 -41 28675 -7
rect 28733 -41 28767 -7
rect 28825 -41 28859 -7
rect 28917 -41 28951 -7
rect 29009 -41 29043 -7
rect 29101 -41 29135 -7
rect 29193 -41 29227 -7
rect 29285 -41 29319 -7
rect 29377 -41 29411 -7
rect 29469 -41 29503 -7
rect 29561 -41 29595 -7
rect 29653 -41 29687 -7
rect 29745 -41 29779 -7
rect 29837 -41 29871 -7
rect 29929 -41 29963 -7
rect 30021 -41 30055 -7
rect 30113 -41 30147 -7
rect 30205 -41 30239 -7
rect 30297 -41 30331 -7
rect 30389 -41 30423 -7
rect 30481 -41 30515 -7
rect 30573 -41 30607 -7
rect 30665 -41 30699 -7
rect 30757 -41 30791 -7
rect 30849 -41 30883 -7
rect 30941 -41 30975 -7
rect 31033 -41 31067 -7
rect 31125 -41 31159 -7
rect 31217 -41 31251 -7
rect 31309 -41 31343 -7
rect 31401 -41 31435 -7
rect 31493 -41 31527 -7
rect 31585 -41 31619 -7
rect 31677 -41 31711 -7
rect 31769 -41 31803 -7
rect 31861 -41 31895 -7
rect 31953 -41 31987 -7
rect 32045 -41 32079 -7
rect 32137 -41 32171 -7
rect 32229 -41 32263 -7
rect 32321 -41 32355 -7
rect 32413 -41 32447 -7
rect 32505 -41 32539 -7
rect 32597 -41 32631 -7
rect 32689 -41 32723 -7
rect 32781 -41 32815 -7
rect 32873 -41 32907 -7
rect 32965 -41 32999 -7
rect 33057 -41 33091 -7
rect 33149 -41 33183 -7
rect 33241 -41 33275 -7
rect 33333 -41 33367 -7
rect 33425 -41 33459 -7
rect 33517 -41 33551 -7
rect 33609 -41 33643 -7
rect 33701 -41 33735 -7
rect 33793 -41 33827 -7
rect 33885 -41 33919 -7
rect 33977 -41 34011 -7
rect 34069 -41 34103 -7
rect 34161 -41 34195 -7
rect 34253 -41 34287 -7
rect 34345 -41 34379 -7
rect 34437 -41 34471 -7
rect 34529 -41 34563 -7
rect 34621 -41 34655 -7
rect 34713 -41 34747 -7
rect 34805 -41 34839 -7
rect 34897 -41 34931 -7
rect 34989 -41 35023 -7
rect 35081 -41 35115 -7
rect 35173 -41 35207 -7
rect 35265 -41 35299 -7
rect 35357 -41 35391 -7
rect 35449 -41 35483 -7
rect 35541 -41 35575 -7
rect 35633 -41 35667 -7
rect 35725 -41 35759 -7
rect 35817 -41 35851 -7
rect 35909 -41 35943 -7
rect 36001 -41 36035 -7
rect 36093 -41 36127 -7
rect 36185 -41 36219 -7
rect 36277 -41 36311 -7
rect 36369 -41 36403 -7
rect 36461 -41 36495 -7
rect 36553 -41 36587 -7
rect 36645 -41 36679 -7
rect 36737 -41 36771 -7
rect 36829 -41 36863 -7
rect 36921 -41 36955 -7
rect 37013 -41 37047 -7
rect 37105 -41 37139 -7
rect 37197 -41 37231 -7
rect 37289 -41 37323 -7
rect 37381 -41 37415 -7
rect 37473 -41 37507 -7
rect 37565 -41 37599 -7
rect 37657 -41 37691 -7
rect 37749 -41 37783 -7
rect 37841 -41 37875 -7
rect 37933 -41 37967 -7
rect 38025 -41 38059 -7
rect 38117 -41 38151 -7
rect 38209 -41 38243 -7
rect 38301 -41 38335 -7
rect 38393 -41 38427 -7
rect 38485 -41 38519 -7
rect 38577 -41 38611 -7
rect 38669 -41 38703 -7
rect 38761 -41 38795 -7
rect 38853 -41 38887 -7
rect 38945 -41 38979 -7
rect 39037 -41 39071 -7
rect 39129 -41 39163 -7
rect 39221 -41 39255 -7
rect 39313 -41 39347 -7
rect 39405 -41 39439 -7
rect 39497 -41 39531 -7
rect 39589 -41 39623 -7
rect 39681 -41 39715 -7
rect 39773 -41 39807 -7
rect 39865 -41 39899 -7
rect 39957 -41 39991 -7
rect 40049 -41 40083 -7
rect 40141 -41 40175 -7
rect 40233 -41 40267 -7
rect 40325 -41 40359 -7
rect 40417 -41 40451 -7
rect 40509 -41 40543 -7
rect 40601 -41 40635 -7
rect 40693 -41 40727 -7
rect 40785 -41 40819 -7
rect 40877 -41 40911 -7
rect 40969 -41 41003 -7
rect 41061 -41 41095 -7
rect 41153 -41 41187 -7
rect 41245 -41 41279 -7
rect 41337 -41 41371 -7
rect 41429 -41 41463 -7
rect 41521 -41 41555 -7
rect 41613 -41 41647 -7
rect 41705 -41 41739 -7
rect 41797 -41 41831 -7
rect 41889 -41 41923 -7
rect 41981 -41 42015 -7
rect 42073 -41 42107 -7
rect 42165 -41 42199 -7
rect 42257 -41 42291 -7
<< nsubdiffcont >>
rect 29 551 63 585
rect 121 551 155 585
rect 213 551 247 585
rect 305 551 339 585
rect 397 551 431 585
rect 489 551 523 585
rect 581 551 615 585
rect 673 551 707 585
rect 765 551 799 585
rect 857 551 891 585
rect 949 551 983 585
rect 1041 551 1075 585
rect 1133 551 1167 585
rect 1225 551 1259 585
rect 1317 551 1351 585
rect 1409 551 1443 585
rect 1501 551 1535 585
rect 1593 551 1627 585
rect 1685 551 1719 585
rect 1777 551 1811 585
rect 1869 551 1903 585
rect 1961 551 1995 585
rect 2053 551 2087 585
rect 2145 551 2179 585
rect 2237 551 2271 585
rect 2329 551 2363 585
rect 2421 551 2455 585
rect 2513 551 2547 585
rect 2605 551 2639 585
rect 2697 551 2731 585
rect 2789 551 2823 585
rect 2881 551 2915 585
rect 2973 551 3007 585
rect 3065 551 3099 585
rect 3157 551 3191 585
rect 3249 551 3283 585
rect 3341 551 3375 585
rect 3433 551 3467 585
rect 3525 551 3559 585
rect 3617 551 3651 585
rect 3709 551 3743 585
rect 3801 551 3835 585
rect 3893 551 3927 585
rect 3985 551 4019 585
rect 4077 551 4111 585
rect 4169 551 4203 585
rect 4261 551 4295 585
rect 4353 551 4387 585
rect 4445 551 4479 585
rect 4537 551 4571 585
rect 4629 551 4663 585
rect 4721 551 4755 585
rect 4813 551 4847 585
rect 4905 551 4939 585
rect 4997 551 5031 585
rect 5089 551 5123 585
rect 5181 551 5215 585
rect 5273 551 5307 585
rect 5365 551 5399 585
rect 5457 551 5491 585
rect 5549 551 5583 585
rect 5641 551 5675 585
rect 5733 551 5767 585
rect 5825 551 5859 585
rect 5917 551 5951 585
rect 6009 551 6043 585
rect 6101 551 6135 585
rect 6193 551 6227 585
rect 6285 551 6319 585
rect 6377 551 6411 585
rect 6469 551 6503 585
rect 6561 551 6595 585
rect 6653 551 6687 585
rect 6745 551 6779 585
rect 6837 551 6871 585
rect 6929 551 6963 585
rect 7021 551 7055 585
rect 7113 551 7147 585
rect 7205 551 7239 585
rect 7297 551 7331 585
rect 7389 551 7423 585
rect 7481 551 7515 585
rect 7573 551 7607 585
rect 7665 551 7699 585
rect 7757 551 7791 585
rect 7849 551 7883 585
rect 7941 551 7975 585
rect 8033 551 8067 585
rect 8125 551 8159 585
rect 8217 551 8251 585
rect 8309 551 8343 585
rect 8401 551 8435 585
rect 8493 551 8527 585
rect 8585 551 8619 585
rect 8677 551 8711 585
rect 8769 551 8803 585
rect 8861 551 8895 585
rect 8953 551 8987 585
rect 9045 551 9079 585
rect 9137 551 9171 585
rect 9229 551 9263 585
rect 9321 551 9355 585
rect 9413 551 9447 585
rect 9505 551 9539 585
rect 9597 551 9631 585
rect 9689 551 9723 585
rect 9781 551 9815 585
rect 9873 551 9907 585
rect 9965 551 9999 585
rect 10057 551 10091 585
rect 10149 551 10183 585
rect 10241 551 10275 585
rect 10333 551 10367 585
rect 10425 551 10459 585
rect 10517 551 10551 585
rect 10609 551 10643 585
rect 10701 551 10735 585
rect 10793 551 10827 585
rect 10885 551 10919 585
rect 10977 551 11011 585
rect 11069 551 11103 585
rect 11161 551 11195 585
rect 11253 551 11287 585
rect 11345 551 11379 585
rect 11437 551 11471 585
rect 11529 551 11563 585
rect 11621 551 11655 585
rect 11713 551 11747 585
rect 11805 551 11839 585
rect 11897 551 11931 585
rect 11989 551 12023 585
rect 12081 551 12115 585
rect 12173 551 12207 585
rect 12265 551 12299 585
rect 12357 551 12391 585
rect 12449 551 12483 585
rect 12541 551 12575 585
rect 12633 551 12667 585
rect 12725 551 12759 585
rect 12817 551 12851 585
rect 12909 551 12943 585
rect 13001 551 13035 585
rect 13093 551 13127 585
rect 13185 551 13219 585
rect 13277 551 13311 585
rect 13369 551 13403 585
rect 13461 551 13495 585
rect 13553 551 13587 585
rect 13645 551 13679 585
rect 13737 551 13771 585
rect 13829 551 13863 585
rect 13921 551 13955 585
rect 14013 551 14047 585
rect 14105 551 14139 585
rect 14197 551 14231 585
rect 14289 551 14323 585
rect 14381 551 14415 585
rect 14473 551 14507 585
rect 14565 551 14599 585
rect 14657 551 14691 585
rect 14749 551 14783 585
rect 14841 551 14875 585
rect 14933 551 14967 585
rect 15025 551 15059 585
rect 15117 551 15151 585
rect 15209 551 15243 585
rect 15301 551 15335 585
rect 15393 551 15427 585
rect 15485 551 15519 585
rect 15577 551 15611 585
rect 15669 551 15703 585
rect 15761 551 15795 585
rect 15853 551 15887 585
rect 15945 551 15979 585
rect 16037 551 16071 585
rect 16129 551 16163 585
rect 16221 551 16255 585
rect 16313 551 16347 585
rect 16405 551 16439 585
rect 16497 551 16531 585
rect 16589 551 16623 585
rect 16681 551 16715 585
rect 16773 551 16807 585
rect 16865 551 16899 585
rect 16957 551 16991 585
rect 17049 551 17083 585
rect 17141 551 17175 585
rect 17233 551 17267 585
rect 17325 551 17359 585
rect 17417 551 17451 585
rect 17509 551 17543 585
rect 17601 551 17635 585
rect 17693 551 17727 585
rect 17785 551 17819 585
rect 17877 551 17911 585
rect 17969 551 18003 585
rect 18061 551 18095 585
rect 18153 551 18187 585
rect 18245 551 18279 585
rect 18337 551 18371 585
rect 18429 551 18463 585
rect 18521 551 18555 585
rect 18613 551 18647 585
rect 18705 551 18739 585
rect 18797 551 18831 585
rect 18889 551 18923 585
rect 18981 551 19015 585
rect 19073 551 19107 585
rect 19165 551 19199 585
rect 19257 551 19291 585
rect 19349 551 19383 585
rect 19441 551 19475 585
rect 19533 551 19567 585
rect 19625 551 19659 585
rect 19717 551 19751 585
rect 19809 551 19843 585
rect 19901 551 19935 585
rect 19993 551 20027 585
rect 20085 551 20119 585
rect 20177 551 20211 585
rect 20269 551 20303 585
rect 20361 551 20395 585
rect 20453 551 20487 585
rect 20545 551 20579 585
rect 20637 551 20671 585
rect 20729 551 20763 585
rect 20821 551 20855 585
rect 20913 551 20947 585
rect 21005 551 21039 585
rect 21097 551 21131 585
rect 21189 551 21223 585
rect 21281 551 21315 585
rect 21373 551 21407 585
rect 21465 551 21499 585
rect 21557 551 21591 585
rect 21649 551 21683 585
rect 21741 551 21775 585
rect 21833 551 21867 585
rect 21925 551 21959 585
rect 22017 551 22051 585
rect 22109 551 22143 585
rect 22201 551 22235 585
rect 22293 551 22327 585
rect 22385 551 22419 585
rect 22477 551 22511 585
rect 22569 551 22603 585
rect 22661 551 22695 585
rect 22753 551 22787 585
rect 22845 551 22879 585
rect 22937 551 22971 585
rect 23029 551 23063 585
rect 23121 551 23155 585
rect 23213 551 23247 585
rect 23305 551 23339 585
rect 23397 551 23431 585
rect 23489 551 23523 585
rect 23581 551 23615 585
rect 23673 551 23707 585
rect 23765 551 23799 585
rect 23857 551 23891 585
rect 23949 551 23983 585
rect 24041 551 24075 585
rect 24133 551 24167 585
rect 24225 551 24259 585
rect 24317 551 24351 585
rect 24409 551 24443 585
rect 24501 551 24535 585
rect 24593 551 24627 585
rect 24685 551 24719 585
rect 24777 551 24811 585
rect 24869 551 24903 585
rect 24961 551 24995 585
rect 25053 551 25087 585
rect 25145 551 25179 585
rect 25237 551 25271 585
rect 25329 551 25363 585
rect 25421 551 25455 585
rect 25513 551 25547 585
rect 25605 551 25639 585
rect 25697 551 25731 585
rect 25789 551 25823 585
rect 25881 551 25915 585
rect 25973 551 26007 585
rect 26065 551 26099 585
rect 26157 551 26191 585
rect 26249 551 26283 585
rect 26341 551 26375 585
rect 26433 551 26467 585
rect 26525 551 26559 585
rect 26617 551 26651 585
rect 26709 551 26743 585
rect 26801 551 26835 585
rect 26893 551 26927 585
rect 26985 551 27019 585
rect 27077 551 27111 585
rect 27169 551 27203 585
rect 27261 551 27295 585
rect 27353 551 27387 585
rect 27445 551 27479 585
rect 27537 551 27571 585
rect 27629 551 27663 585
rect 27721 551 27755 585
rect 27813 551 27847 585
rect 27905 551 27939 585
rect 27997 551 28031 585
rect 28089 551 28123 585
rect 28181 551 28215 585
rect 28273 551 28307 585
rect 28365 551 28399 585
rect 28457 551 28491 585
rect 28549 551 28583 585
rect 28641 551 28675 585
rect 28733 551 28767 585
rect 28825 551 28859 585
rect 28917 551 28951 585
rect 29009 551 29043 585
rect 29101 551 29135 585
rect 29193 551 29227 585
rect 29285 551 29319 585
rect 29377 551 29411 585
rect 29469 551 29503 585
rect 29561 551 29595 585
rect 29653 551 29687 585
rect 29745 551 29779 585
rect 29837 551 29871 585
rect 29929 551 29963 585
rect 30021 551 30055 585
rect 30113 551 30147 585
rect 30205 551 30239 585
rect 30297 551 30331 585
rect 30389 551 30423 585
rect 30481 551 30515 585
rect 30573 551 30607 585
rect 30665 551 30699 585
rect 30757 551 30791 585
rect 30849 551 30883 585
rect 30941 551 30975 585
rect 31033 551 31067 585
rect 31125 551 31159 585
rect 31217 551 31251 585
rect 31309 551 31343 585
rect 31401 551 31435 585
rect 31493 551 31527 585
rect 31585 551 31619 585
rect 31677 551 31711 585
rect 31769 551 31803 585
rect 31861 551 31895 585
rect 31953 551 31987 585
rect 32045 551 32079 585
rect 32137 551 32171 585
rect 32229 551 32263 585
rect 32321 551 32355 585
rect 32413 551 32447 585
rect 32505 551 32539 585
rect 32597 551 32631 585
rect 32689 551 32723 585
rect 32781 551 32815 585
rect 32873 551 32907 585
rect 32965 551 32999 585
rect 33057 551 33091 585
rect 33149 551 33183 585
rect 33241 551 33275 585
rect 33333 551 33367 585
rect 33425 551 33459 585
rect 33517 551 33551 585
rect 33609 551 33643 585
rect 33701 551 33735 585
rect 33793 551 33827 585
rect 33885 551 33919 585
rect 33977 551 34011 585
rect 34069 551 34103 585
rect 34161 551 34195 585
rect 34253 551 34287 585
rect 34345 551 34379 585
rect 34437 551 34471 585
rect 34529 551 34563 585
rect 34621 551 34655 585
rect 34713 551 34747 585
rect 34805 551 34839 585
rect 34897 551 34931 585
rect 34989 551 35023 585
rect 35081 551 35115 585
rect 35173 551 35207 585
rect 35265 551 35299 585
rect 35357 551 35391 585
rect 35449 551 35483 585
rect 35541 551 35575 585
rect 35633 551 35667 585
rect 35725 551 35759 585
rect 35817 551 35851 585
rect 35909 551 35943 585
rect 36001 551 36035 585
rect 36093 551 36127 585
rect 36185 551 36219 585
rect 36277 551 36311 585
rect 36369 551 36403 585
rect 36461 551 36495 585
rect 36553 551 36587 585
rect 36645 551 36679 585
rect 36737 551 36771 585
rect 36829 551 36863 585
rect 36921 551 36955 585
rect 37013 551 37047 585
rect 37105 551 37139 585
rect 37197 551 37231 585
rect 37289 551 37323 585
rect 37381 551 37415 585
rect 37473 551 37507 585
rect 37565 551 37599 585
rect 37657 551 37691 585
rect 37749 551 37783 585
rect 37841 551 37875 585
rect 37933 551 37967 585
rect 38025 551 38059 585
rect 38117 551 38151 585
rect 38209 551 38243 585
rect 38301 551 38335 585
rect 38393 551 38427 585
rect 38485 551 38519 585
rect 38577 551 38611 585
rect 38669 551 38703 585
rect 38761 551 38795 585
rect 38853 551 38887 585
rect 38945 551 38979 585
rect 39037 551 39071 585
rect 39129 551 39163 585
rect 39221 551 39255 585
rect 39313 551 39347 585
rect 39405 551 39439 585
rect 39497 551 39531 585
rect 39589 551 39623 585
rect 39681 551 39715 585
rect 39773 551 39807 585
rect 39865 551 39899 585
rect 39957 551 39991 585
rect 40049 551 40083 585
rect 40141 551 40175 585
rect 40233 551 40267 585
rect 40325 551 40359 585
rect 40417 551 40451 585
rect 40509 551 40543 585
rect 40601 551 40635 585
rect 40693 551 40727 585
rect 40785 551 40819 585
rect 40877 551 40911 585
rect 40969 551 41003 585
rect 41061 551 41095 585
rect 41153 551 41187 585
rect 41245 551 41279 585
rect 41337 551 41371 585
rect 41429 551 41463 585
rect 41521 551 41555 585
rect 41613 551 41647 585
rect 41705 551 41739 585
rect 41797 551 41831 585
rect 41889 551 41923 585
rect 41981 551 42015 585
rect 42073 551 42107 585
rect 42165 551 42199 585
rect 42257 551 42291 585
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 430 497 460 523
rect 522 497 552 523
rect 621 497 651 523
rect 761 497 791 523
rect 858 497 888 523
rect 1055 497 1085 523
rect 1154 497 1184 523
rect 1240 497 1270 523
rect 1324 497 1354 523
rect 1432 497 1462 523
rect 1516 497 1546 523
rect 1680 497 1710 523
rect 1899 497 1929 523
rect 1996 497 2026 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 265 76 318
rect 163 274 193 363
rect 430 326 460 413
rect 522 375 552 413
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 331 310 460 326
rect 506 365 572 375
rect 506 331 522 365
rect 556 331 572 365
rect 506 321 572 331
rect 331 276 341 310
rect 375 296 460 310
rect 375 276 448 296
rect 621 279 651 413
rect 761 355 791 413
rect 761 339 816 355
rect 761 305 771 339
rect 805 305 816 339
rect 761 289 816 305
rect 331 260 448 276
rect 118 220 193 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 418 131 448 260
rect 513 249 651 279
rect 513 219 544 249
rect 490 203 544 219
rect 490 169 500 203
rect 534 169 544 203
rect 490 153 544 169
rect 586 197 652 207
rect 586 163 602 197
rect 636 163 652 197
rect 586 153 652 163
rect 513 119 543 153
rect 609 119 639 153
rect 775 131 805 289
rect 858 219 888 413
rect 1055 314 1085 329
rect 979 284 1085 314
rect 979 267 1009 284
rect 943 251 1009 267
rect 847 203 901 219
rect 847 169 857 203
rect 891 169 901 203
rect 943 217 953 251
rect 987 217 1009 251
rect 1154 279 1184 413
rect 1240 381 1270 413
rect 1226 365 1280 381
rect 1226 331 1236 365
rect 1270 331 1280 365
rect 1226 315 1280 331
rect 1154 267 1204 279
rect 1154 255 1217 267
rect 1154 249 1241 255
rect 1175 239 1241 249
rect 1175 237 1197 239
rect 943 201 1009 217
rect 979 175 1009 201
rect 1078 191 1145 207
rect 847 153 901 169
rect 847 131 877 153
rect 1078 157 1101 191
rect 1135 157 1145 191
rect 1078 141 1145 157
rect 1187 205 1197 237
rect 1231 205 1241 239
rect 1187 189 1241 205
rect 1324 229 1354 413
rect 1432 257 1462 413
rect 1516 365 1546 413
rect 1504 349 1558 365
rect 1504 315 1514 349
rect 1548 315 1558 349
rect 1504 299 1558 315
rect 1427 241 1481 257
rect 1324 213 1385 229
rect 1324 193 1341 213
rect 1078 119 1108 141
rect 1187 119 1217 189
rect 1283 179 1341 193
rect 1375 179 1385 213
rect 1427 207 1437 241
rect 1471 207 1481 241
rect 1427 191 1481 207
rect 1283 163 1385 179
rect 1283 131 1313 163
rect 1432 131 1462 191
rect 1523 131 1553 299
rect 1899 333 1929 369
rect 1888 303 1929 333
rect 1680 265 1710 297
rect 1888 265 1918 303
rect 2195 491 2225 517
rect 2279 491 2309 517
rect 2546 497 2576 523
rect 2638 497 2668 523
rect 2737 497 2767 523
rect 2877 497 2907 523
rect 2974 497 3004 523
rect 3171 497 3201 523
rect 3270 497 3300 523
rect 3356 497 3386 523
rect 3440 497 3470 523
rect 3548 497 3578 523
rect 3632 497 3662 523
rect 3796 497 3826 523
rect 4015 497 4045 523
rect 4112 497 4142 523
rect 2195 348 2225 363
rect 2162 318 2225 348
rect 1996 265 2026 297
rect 2162 265 2192 318
rect 2279 274 2309 363
rect 2546 326 2576 413
rect 2638 375 2668 413
rect 1609 249 1918 265
rect 1609 215 1637 249
rect 1671 215 1918 249
rect 1609 199 1918 215
rect 1967 249 2026 265
rect 1967 215 1977 249
rect 2011 215 2026 249
rect 1967 199 2026 215
rect 2138 249 2192 265
rect 2138 215 2148 249
rect 2182 215 2192 249
rect 2234 264 2309 274
rect 2234 230 2250 264
rect 2284 230 2309 264
rect 2447 310 2576 326
rect 2622 365 2688 375
rect 2622 331 2638 365
rect 2672 331 2688 365
rect 2622 321 2688 331
rect 2447 276 2457 310
rect 2491 296 2576 310
rect 2491 276 2564 296
rect 2737 279 2767 413
rect 2877 355 2907 413
rect 2877 339 2932 355
rect 2877 305 2887 339
rect 2921 305 2932 339
rect 2877 289 2932 305
rect 2447 260 2564 276
rect 2234 220 2309 230
rect 2138 199 2192 215
rect 1711 177 1741 199
rect 1888 176 1918 199
rect 1996 177 2026 199
rect 1888 146 1929 176
rect 1899 131 1929 146
rect 2162 176 2192 199
rect 2162 146 2225 176
rect 2195 131 2225 146
rect 2279 131 2309 220
rect 2534 131 2564 260
rect 2629 249 2767 279
rect 2629 219 2660 249
rect 2606 203 2660 219
rect 2606 169 2616 203
rect 2650 169 2660 203
rect 2606 153 2660 169
rect 2702 197 2768 207
rect 2702 163 2718 197
rect 2752 163 2768 197
rect 2702 153 2768 163
rect 2629 119 2659 153
rect 2725 119 2755 153
rect 2891 131 2921 289
rect 2974 219 3004 413
rect 3171 314 3201 329
rect 3095 284 3201 314
rect 3095 267 3125 284
rect 3059 251 3125 267
rect 2963 203 3017 219
rect 2963 169 2973 203
rect 3007 169 3017 203
rect 3059 217 3069 251
rect 3103 217 3125 251
rect 3270 279 3300 413
rect 3356 381 3386 413
rect 3342 365 3396 381
rect 3342 331 3352 365
rect 3386 331 3396 365
rect 3342 315 3396 331
rect 3270 267 3320 279
rect 3270 255 3333 267
rect 3270 249 3357 255
rect 3291 239 3357 249
rect 3291 237 3313 239
rect 3059 201 3125 217
rect 3095 175 3125 201
rect 3194 191 3261 207
rect 2963 153 3017 169
rect 2963 131 2993 153
rect 3194 157 3217 191
rect 3251 157 3261 191
rect 3194 141 3261 157
rect 3303 205 3313 237
rect 3347 205 3357 239
rect 3303 189 3357 205
rect 3440 229 3470 413
rect 3548 257 3578 413
rect 3632 365 3662 413
rect 3620 349 3674 365
rect 3620 315 3630 349
rect 3664 315 3674 349
rect 3620 299 3674 315
rect 3543 241 3597 257
rect 3440 213 3501 229
rect 3440 193 3457 213
rect 3194 119 3224 141
rect 3303 119 3333 189
rect 3399 179 3457 193
rect 3491 179 3501 213
rect 3543 207 3553 241
rect 3587 207 3597 241
rect 3543 191 3597 207
rect 3399 163 3501 179
rect 3399 131 3429 163
rect 3548 131 3578 191
rect 3639 131 3669 299
rect 4015 333 4045 369
rect 4004 303 4045 333
rect 3796 265 3826 297
rect 4004 265 4034 303
rect 4311 491 4341 517
rect 4395 491 4425 517
rect 4662 497 4692 523
rect 4754 497 4784 523
rect 4853 497 4883 523
rect 4993 497 5023 523
rect 5090 497 5120 523
rect 5287 497 5317 523
rect 5386 497 5416 523
rect 5472 497 5502 523
rect 5556 497 5586 523
rect 5664 497 5694 523
rect 5748 497 5778 523
rect 5912 497 5942 523
rect 6131 497 6161 523
rect 6228 497 6258 523
rect 4311 348 4341 363
rect 4278 318 4341 348
rect 4112 265 4142 297
rect 4278 265 4308 318
rect 4395 274 4425 363
rect 4662 326 4692 413
rect 4754 375 4784 413
rect 3725 249 4034 265
rect 3725 215 3753 249
rect 3787 215 4034 249
rect 3725 199 4034 215
rect 4083 249 4142 265
rect 4083 215 4093 249
rect 4127 215 4142 249
rect 4083 199 4142 215
rect 4254 249 4308 265
rect 4254 215 4264 249
rect 4298 215 4308 249
rect 4350 264 4425 274
rect 4350 230 4366 264
rect 4400 230 4425 264
rect 4563 310 4692 326
rect 4738 365 4804 375
rect 4738 331 4754 365
rect 4788 331 4804 365
rect 4738 321 4804 331
rect 4563 276 4573 310
rect 4607 296 4692 310
rect 4607 276 4680 296
rect 4853 279 4883 413
rect 4993 355 5023 413
rect 4993 339 5048 355
rect 4993 305 5003 339
rect 5037 305 5048 339
rect 4993 289 5048 305
rect 4563 260 4680 276
rect 4350 220 4425 230
rect 4254 199 4308 215
rect 3827 177 3857 199
rect 4004 176 4034 199
rect 4112 177 4142 199
rect 4004 146 4045 176
rect 4015 131 4045 146
rect 4278 176 4308 199
rect 4278 146 4341 176
rect 4311 131 4341 146
rect 4395 131 4425 220
rect 4650 131 4680 260
rect 4745 249 4883 279
rect 4745 219 4776 249
rect 4722 203 4776 219
rect 4722 169 4732 203
rect 4766 169 4776 203
rect 4722 153 4776 169
rect 4818 197 4884 207
rect 4818 163 4834 197
rect 4868 163 4884 197
rect 4818 153 4884 163
rect 4745 119 4775 153
rect 4841 119 4871 153
rect 5007 131 5037 289
rect 5090 219 5120 413
rect 5287 314 5317 329
rect 5211 284 5317 314
rect 5211 267 5241 284
rect 5175 251 5241 267
rect 5079 203 5133 219
rect 5079 169 5089 203
rect 5123 169 5133 203
rect 5175 217 5185 251
rect 5219 217 5241 251
rect 5386 279 5416 413
rect 5472 381 5502 413
rect 5458 365 5512 381
rect 5458 331 5468 365
rect 5502 331 5512 365
rect 5458 315 5512 331
rect 5386 267 5436 279
rect 5386 255 5449 267
rect 5386 249 5473 255
rect 5407 239 5473 249
rect 5407 237 5429 239
rect 5175 201 5241 217
rect 5211 175 5241 201
rect 5310 191 5377 207
rect 5079 153 5133 169
rect 5079 131 5109 153
rect 5310 157 5333 191
rect 5367 157 5377 191
rect 5310 141 5377 157
rect 5419 205 5429 237
rect 5463 205 5473 239
rect 5419 189 5473 205
rect 5556 229 5586 413
rect 5664 257 5694 413
rect 5748 365 5778 413
rect 5736 349 5790 365
rect 5736 315 5746 349
rect 5780 315 5790 349
rect 5736 299 5790 315
rect 5659 241 5713 257
rect 5556 213 5617 229
rect 5556 193 5573 213
rect 5310 119 5340 141
rect 5419 119 5449 189
rect 5515 179 5573 193
rect 5607 179 5617 213
rect 5659 207 5669 241
rect 5703 207 5713 241
rect 5659 191 5713 207
rect 5515 163 5617 179
rect 5515 131 5545 163
rect 5664 131 5694 191
rect 5755 131 5785 299
rect 6131 333 6161 369
rect 6120 303 6161 333
rect 5912 265 5942 297
rect 6120 265 6150 303
rect 6427 491 6457 517
rect 6511 491 6541 517
rect 6778 497 6808 523
rect 6870 497 6900 523
rect 6969 497 6999 523
rect 7109 497 7139 523
rect 7206 497 7236 523
rect 7403 497 7433 523
rect 7502 497 7532 523
rect 7588 497 7618 523
rect 7672 497 7702 523
rect 7780 497 7810 523
rect 7864 497 7894 523
rect 8028 497 8058 523
rect 8247 497 8277 523
rect 8344 497 8374 523
rect 6427 348 6457 363
rect 6394 318 6457 348
rect 6228 265 6258 297
rect 6394 265 6424 318
rect 6511 274 6541 363
rect 6778 326 6808 413
rect 6870 375 6900 413
rect 5841 249 6150 265
rect 5841 215 5869 249
rect 5903 215 6150 249
rect 5841 199 6150 215
rect 6199 249 6258 265
rect 6199 215 6209 249
rect 6243 215 6258 249
rect 6199 199 6258 215
rect 6370 249 6424 265
rect 6370 215 6380 249
rect 6414 215 6424 249
rect 6466 264 6541 274
rect 6466 230 6482 264
rect 6516 230 6541 264
rect 6679 310 6808 326
rect 6854 365 6920 375
rect 6854 331 6870 365
rect 6904 331 6920 365
rect 6854 321 6920 331
rect 6679 276 6689 310
rect 6723 296 6808 310
rect 6723 276 6796 296
rect 6969 279 6999 413
rect 7109 355 7139 413
rect 7109 339 7164 355
rect 7109 305 7119 339
rect 7153 305 7164 339
rect 7109 289 7164 305
rect 6679 260 6796 276
rect 6466 220 6541 230
rect 6370 199 6424 215
rect 5943 177 5973 199
rect 6120 176 6150 199
rect 6228 177 6258 199
rect 6120 146 6161 176
rect 6131 131 6161 146
rect 6394 176 6424 199
rect 6394 146 6457 176
rect 6427 131 6457 146
rect 6511 131 6541 220
rect 6766 131 6796 260
rect 6861 249 6999 279
rect 6861 219 6892 249
rect 6838 203 6892 219
rect 6838 169 6848 203
rect 6882 169 6892 203
rect 6838 153 6892 169
rect 6934 197 7000 207
rect 6934 163 6950 197
rect 6984 163 7000 197
rect 6934 153 7000 163
rect 6861 119 6891 153
rect 6957 119 6987 153
rect 7123 131 7153 289
rect 7206 219 7236 413
rect 7403 314 7433 329
rect 7327 284 7433 314
rect 7327 267 7357 284
rect 7291 251 7357 267
rect 7195 203 7249 219
rect 7195 169 7205 203
rect 7239 169 7249 203
rect 7291 217 7301 251
rect 7335 217 7357 251
rect 7502 279 7532 413
rect 7588 381 7618 413
rect 7574 365 7628 381
rect 7574 331 7584 365
rect 7618 331 7628 365
rect 7574 315 7628 331
rect 7502 267 7552 279
rect 7502 255 7565 267
rect 7502 249 7589 255
rect 7523 239 7589 249
rect 7523 237 7545 239
rect 7291 201 7357 217
rect 7327 175 7357 201
rect 7426 191 7493 207
rect 7195 153 7249 169
rect 7195 131 7225 153
rect 7426 157 7449 191
rect 7483 157 7493 191
rect 7426 141 7493 157
rect 7535 205 7545 237
rect 7579 205 7589 239
rect 7535 189 7589 205
rect 7672 229 7702 413
rect 7780 257 7810 413
rect 7864 365 7894 413
rect 7852 349 7906 365
rect 7852 315 7862 349
rect 7896 315 7906 349
rect 7852 299 7906 315
rect 7775 241 7829 257
rect 7672 213 7733 229
rect 7672 193 7689 213
rect 7426 119 7456 141
rect 7535 119 7565 189
rect 7631 179 7689 193
rect 7723 179 7733 213
rect 7775 207 7785 241
rect 7819 207 7829 241
rect 7775 191 7829 207
rect 7631 163 7733 179
rect 7631 131 7661 163
rect 7780 131 7810 191
rect 7871 131 7901 299
rect 8247 333 8277 369
rect 8236 303 8277 333
rect 8028 265 8058 297
rect 8236 265 8266 303
rect 8543 491 8573 517
rect 8627 491 8657 517
rect 8894 497 8924 523
rect 8986 497 9016 523
rect 9085 497 9115 523
rect 9225 497 9255 523
rect 9322 497 9352 523
rect 9519 497 9549 523
rect 9618 497 9648 523
rect 9704 497 9734 523
rect 9788 497 9818 523
rect 9896 497 9926 523
rect 9980 497 10010 523
rect 10144 497 10174 523
rect 10363 497 10393 523
rect 10460 497 10490 523
rect 8543 348 8573 363
rect 8510 318 8573 348
rect 8344 265 8374 297
rect 8510 265 8540 318
rect 8627 274 8657 363
rect 8894 326 8924 413
rect 8986 375 9016 413
rect 7957 249 8266 265
rect 7957 215 7985 249
rect 8019 215 8266 249
rect 7957 199 8266 215
rect 8315 249 8374 265
rect 8315 215 8325 249
rect 8359 215 8374 249
rect 8315 199 8374 215
rect 8486 249 8540 265
rect 8486 215 8496 249
rect 8530 215 8540 249
rect 8582 264 8657 274
rect 8582 230 8598 264
rect 8632 230 8657 264
rect 8795 310 8924 326
rect 8970 365 9036 375
rect 8970 331 8986 365
rect 9020 331 9036 365
rect 8970 321 9036 331
rect 8795 276 8805 310
rect 8839 296 8924 310
rect 8839 276 8912 296
rect 9085 279 9115 413
rect 9225 355 9255 413
rect 9225 339 9280 355
rect 9225 305 9235 339
rect 9269 305 9280 339
rect 9225 289 9280 305
rect 8795 260 8912 276
rect 8582 220 8657 230
rect 8486 199 8540 215
rect 8059 177 8089 199
rect 8236 176 8266 199
rect 8344 177 8374 199
rect 8236 146 8277 176
rect 8247 131 8277 146
rect 8510 176 8540 199
rect 8510 146 8573 176
rect 8543 131 8573 146
rect 8627 131 8657 220
rect 8882 131 8912 260
rect 8977 249 9115 279
rect 8977 219 9008 249
rect 8954 203 9008 219
rect 8954 169 8964 203
rect 8998 169 9008 203
rect 8954 153 9008 169
rect 9050 197 9116 207
rect 9050 163 9066 197
rect 9100 163 9116 197
rect 9050 153 9116 163
rect 8977 119 9007 153
rect 9073 119 9103 153
rect 9239 131 9269 289
rect 9322 219 9352 413
rect 9519 314 9549 329
rect 9443 284 9549 314
rect 9443 267 9473 284
rect 9407 251 9473 267
rect 9311 203 9365 219
rect 9311 169 9321 203
rect 9355 169 9365 203
rect 9407 217 9417 251
rect 9451 217 9473 251
rect 9618 279 9648 413
rect 9704 381 9734 413
rect 9690 365 9744 381
rect 9690 331 9700 365
rect 9734 331 9744 365
rect 9690 315 9744 331
rect 9618 267 9668 279
rect 9618 255 9681 267
rect 9618 249 9705 255
rect 9639 239 9705 249
rect 9639 237 9661 239
rect 9407 201 9473 217
rect 9443 175 9473 201
rect 9542 191 9609 207
rect 9311 153 9365 169
rect 9311 131 9341 153
rect 9542 157 9565 191
rect 9599 157 9609 191
rect 9542 141 9609 157
rect 9651 205 9661 237
rect 9695 205 9705 239
rect 9651 189 9705 205
rect 9788 229 9818 413
rect 9896 257 9926 413
rect 9980 365 10010 413
rect 9968 349 10022 365
rect 9968 315 9978 349
rect 10012 315 10022 349
rect 9968 299 10022 315
rect 9891 241 9945 257
rect 9788 213 9849 229
rect 9788 193 9805 213
rect 9542 119 9572 141
rect 9651 119 9681 189
rect 9747 179 9805 193
rect 9839 179 9849 213
rect 9891 207 9901 241
rect 9935 207 9945 241
rect 9891 191 9945 207
rect 9747 163 9849 179
rect 9747 131 9777 163
rect 9896 131 9926 191
rect 9987 131 10017 299
rect 10363 333 10393 369
rect 10352 303 10393 333
rect 10144 265 10174 297
rect 10352 265 10382 303
rect 10659 491 10689 517
rect 10743 491 10773 517
rect 11010 497 11040 523
rect 11102 497 11132 523
rect 11201 497 11231 523
rect 11341 497 11371 523
rect 11438 497 11468 523
rect 11635 497 11665 523
rect 11734 497 11764 523
rect 11820 497 11850 523
rect 11904 497 11934 523
rect 12012 497 12042 523
rect 12096 497 12126 523
rect 12260 497 12290 523
rect 12479 497 12509 523
rect 12576 497 12606 523
rect 10659 348 10689 363
rect 10626 318 10689 348
rect 10460 265 10490 297
rect 10626 265 10656 318
rect 10743 274 10773 363
rect 11010 326 11040 413
rect 11102 375 11132 413
rect 10073 249 10382 265
rect 10073 215 10101 249
rect 10135 215 10382 249
rect 10073 199 10382 215
rect 10431 249 10490 265
rect 10431 215 10441 249
rect 10475 215 10490 249
rect 10431 199 10490 215
rect 10602 249 10656 265
rect 10602 215 10612 249
rect 10646 215 10656 249
rect 10698 264 10773 274
rect 10698 230 10714 264
rect 10748 230 10773 264
rect 10911 310 11040 326
rect 11086 365 11152 375
rect 11086 331 11102 365
rect 11136 331 11152 365
rect 11086 321 11152 331
rect 10911 276 10921 310
rect 10955 296 11040 310
rect 10955 276 11028 296
rect 11201 279 11231 413
rect 11341 355 11371 413
rect 11341 339 11396 355
rect 11341 305 11351 339
rect 11385 305 11396 339
rect 11341 289 11396 305
rect 10911 260 11028 276
rect 10698 220 10773 230
rect 10602 199 10656 215
rect 10175 177 10205 199
rect 10352 176 10382 199
rect 10460 177 10490 199
rect 10352 146 10393 176
rect 10363 131 10393 146
rect 10626 176 10656 199
rect 10626 146 10689 176
rect 10659 131 10689 146
rect 10743 131 10773 220
rect 10998 131 11028 260
rect 11093 249 11231 279
rect 11093 219 11124 249
rect 11070 203 11124 219
rect 11070 169 11080 203
rect 11114 169 11124 203
rect 11070 153 11124 169
rect 11166 197 11232 207
rect 11166 163 11182 197
rect 11216 163 11232 197
rect 11166 153 11232 163
rect 11093 119 11123 153
rect 11189 119 11219 153
rect 11355 131 11385 289
rect 11438 219 11468 413
rect 11635 314 11665 329
rect 11559 284 11665 314
rect 11559 267 11589 284
rect 11523 251 11589 267
rect 11427 203 11481 219
rect 11427 169 11437 203
rect 11471 169 11481 203
rect 11523 217 11533 251
rect 11567 217 11589 251
rect 11734 279 11764 413
rect 11820 381 11850 413
rect 11806 365 11860 381
rect 11806 331 11816 365
rect 11850 331 11860 365
rect 11806 315 11860 331
rect 11734 267 11784 279
rect 11734 255 11797 267
rect 11734 249 11821 255
rect 11755 239 11821 249
rect 11755 237 11777 239
rect 11523 201 11589 217
rect 11559 175 11589 201
rect 11658 191 11725 207
rect 11427 153 11481 169
rect 11427 131 11457 153
rect 11658 157 11681 191
rect 11715 157 11725 191
rect 11658 141 11725 157
rect 11767 205 11777 237
rect 11811 205 11821 239
rect 11767 189 11821 205
rect 11904 229 11934 413
rect 12012 257 12042 413
rect 12096 365 12126 413
rect 12084 349 12138 365
rect 12084 315 12094 349
rect 12128 315 12138 349
rect 12084 299 12138 315
rect 12007 241 12061 257
rect 11904 213 11965 229
rect 11904 193 11921 213
rect 11658 119 11688 141
rect 11767 119 11797 189
rect 11863 179 11921 193
rect 11955 179 11965 213
rect 12007 207 12017 241
rect 12051 207 12061 241
rect 12007 191 12061 207
rect 11863 163 11965 179
rect 11863 131 11893 163
rect 12012 131 12042 191
rect 12103 131 12133 299
rect 12479 333 12509 369
rect 12468 303 12509 333
rect 12260 265 12290 297
rect 12468 265 12498 303
rect 12775 491 12805 517
rect 12859 491 12889 517
rect 13126 497 13156 523
rect 13218 497 13248 523
rect 13317 497 13347 523
rect 13457 497 13487 523
rect 13554 497 13584 523
rect 13751 497 13781 523
rect 13850 497 13880 523
rect 13936 497 13966 523
rect 14020 497 14050 523
rect 14128 497 14158 523
rect 14212 497 14242 523
rect 14376 497 14406 523
rect 14595 497 14625 523
rect 14692 497 14722 523
rect 12775 348 12805 363
rect 12742 318 12805 348
rect 12576 265 12606 297
rect 12742 265 12772 318
rect 12859 274 12889 363
rect 13126 326 13156 413
rect 13218 375 13248 413
rect 12189 249 12498 265
rect 12189 215 12217 249
rect 12251 215 12498 249
rect 12189 199 12498 215
rect 12547 249 12606 265
rect 12547 215 12557 249
rect 12591 215 12606 249
rect 12547 199 12606 215
rect 12718 249 12772 265
rect 12718 215 12728 249
rect 12762 215 12772 249
rect 12814 264 12889 274
rect 12814 230 12830 264
rect 12864 230 12889 264
rect 13027 310 13156 326
rect 13202 365 13268 375
rect 13202 331 13218 365
rect 13252 331 13268 365
rect 13202 321 13268 331
rect 13027 276 13037 310
rect 13071 296 13156 310
rect 13071 276 13144 296
rect 13317 279 13347 413
rect 13457 355 13487 413
rect 13457 339 13512 355
rect 13457 305 13467 339
rect 13501 305 13512 339
rect 13457 289 13512 305
rect 13027 260 13144 276
rect 12814 220 12889 230
rect 12718 199 12772 215
rect 12291 177 12321 199
rect 12468 176 12498 199
rect 12576 177 12606 199
rect 12468 146 12509 176
rect 12479 131 12509 146
rect 12742 176 12772 199
rect 12742 146 12805 176
rect 12775 131 12805 146
rect 12859 131 12889 220
rect 13114 131 13144 260
rect 13209 249 13347 279
rect 13209 219 13240 249
rect 13186 203 13240 219
rect 13186 169 13196 203
rect 13230 169 13240 203
rect 13186 153 13240 169
rect 13282 197 13348 207
rect 13282 163 13298 197
rect 13332 163 13348 197
rect 13282 153 13348 163
rect 13209 119 13239 153
rect 13305 119 13335 153
rect 13471 131 13501 289
rect 13554 219 13584 413
rect 13751 314 13781 329
rect 13675 284 13781 314
rect 13675 267 13705 284
rect 13639 251 13705 267
rect 13543 203 13597 219
rect 13543 169 13553 203
rect 13587 169 13597 203
rect 13639 217 13649 251
rect 13683 217 13705 251
rect 13850 279 13880 413
rect 13936 381 13966 413
rect 13922 365 13976 381
rect 13922 331 13932 365
rect 13966 331 13976 365
rect 13922 315 13976 331
rect 13850 267 13900 279
rect 13850 255 13913 267
rect 13850 249 13937 255
rect 13871 239 13937 249
rect 13871 237 13893 239
rect 13639 201 13705 217
rect 13675 175 13705 201
rect 13774 191 13841 207
rect 13543 153 13597 169
rect 13543 131 13573 153
rect 13774 157 13797 191
rect 13831 157 13841 191
rect 13774 141 13841 157
rect 13883 205 13893 237
rect 13927 205 13937 239
rect 13883 189 13937 205
rect 14020 229 14050 413
rect 14128 257 14158 413
rect 14212 365 14242 413
rect 14200 349 14254 365
rect 14200 315 14210 349
rect 14244 315 14254 349
rect 14200 299 14254 315
rect 14123 241 14177 257
rect 14020 213 14081 229
rect 14020 193 14037 213
rect 13774 119 13804 141
rect 13883 119 13913 189
rect 13979 179 14037 193
rect 14071 179 14081 213
rect 14123 207 14133 241
rect 14167 207 14177 241
rect 14123 191 14177 207
rect 13979 163 14081 179
rect 13979 131 14009 163
rect 14128 131 14158 191
rect 14219 131 14249 299
rect 14595 333 14625 369
rect 14584 303 14625 333
rect 14376 265 14406 297
rect 14584 265 14614 303
rect 14891 491 14921 517
rect 14975 491 15005 517
rect 15242 497 15272 523
rect 15334 497 15364 523
rect 15433 497 15463 523
rect 15573 497 15603 523
rect 15670 497 15700 523
rect 15867 497 15897 523
rect 15966 497 15996 523
rect 16052 497 16082 523
rect 16136 497 16166 523
rect 16244 497 16274 523
rect 16328 497 16358 523
rect 16492 497 16522 523
rect 16711 497 16741 523
rect 16808 497 16838 523
rect 14891 348 14921 363
rect 14858 318 14921 348
rect 14692 265 14722 297
rect 14858 265 14888 318
rect 14975 274 15005 363
rect 15242 326 15272 413
rect 15334 375 15364 413
rect 14305 249 14614 265
rect 14305 215 14333 249
rect 14367 215 14614 249
rect 14305 199 14614 215
rect 14663 249 14722 265
rect 14663 215 14673 249
rect 14707 215 14722 249
rect 14663 199 14722 215
rect 14834 249 14888 265
rect 14834 215 14844 249
rect 14878 215 14888 249
rect 14930 264 15005 274
rect 14930 230 14946 264
rect 14980 230 15005 264
rect 15143 310 15272 326
rect 15318 365 15384 375
rect 15318 331 15334 365
rect 15368 331 15384 365
rect 15318 321 15384 331
rect 15143 276 15153 310
rect 15187 296 15272 310
rect 15187 276 15260 296
rect 15433 279 15463 413
rect 15573 355 15603 413
rect 15573 339 15628 355
rect 15573 305 15583 339
rect 15617 305 15628 339
rect 15573 289 15628 305
rect 15143 260 15260 276
rect 14930 220 15005 230
rect 14834 199 14888 215
rect 14407 177 14437 199
rect 14584 176 14614 199
rect 14692 177 14722 199
rect 14584 146 14625 176
rect 14595 131 14625 146
rect 14858 176 14888 199
rect 14858 146 14921 176
rect 14891 131 14921 146
rect 14975 131 15005 220
rect 15230 131 15260 260
rect 15325 249 15463 279
rect 15325 219 15356 249
rect 15302 203 15356 219
rect 15302 169 15312 203
rect 15346 169 15356 203
rect 15302 153 15356 169
rect 15398 197 15464 207
rect 15398 163 15414 197
rect 15448 163 15464 197
rect 15398 153 15464 163
rect 15325 119 15355 153
rect 15421 119 15451 153
rect 15587 131 15617 289
rect 15670 219 15700 413
rect 15867 314 15897 329
rect 15791 284 15897 314
rect 15791 267 15821 284
rect 15755 251 15821 267
rect 15659 203 15713 219
rect 15659 169 15669 203
rect 15703 169 15713 203
rect 15755 217 15765 251
rect 15799 217 15821 251
rect 15966 279 15996 413
rect 16052 381 16082 413
rect 16038 365 16092 381
rect 16038 331 16048 365
rect 16082 331 16092 365
rect 16038 315 16092 331
rect 15966 267 16016 279
rect 15966 255 16029 267
rect 15966 249 16053 255
rect 15987 239 16053 249
rect 15987 237 16009 239
rect 15755 201 15821 217
rect 15791 175 15821 201
rect 15890 191 15957 207
rect 15659 153 15713 169
rect 15659 131 15689 153
rect 15890 157 15913 191
rect 15947 157 15957 191
rect 15890 141 15957 157
rect 15999 205 16009 237
rect 16043 205 16053 239
rect 15999 189 16053 205
rect 16136 229 16166 413
rect 16244 257 16274 413
rect 16328 365 16358 413
rect 16316 349 16370 365
rect 16316 315 16326 349
rect 16360 315 16370 349
rect 16316 299 16370 315
rect 16239 241 16293 257
rect 16136 213 16197 229
rect 16136 193 16153 213
rect 15890 119 15920 141
rect 15999 119 16029 189
rect 16095 179 16153 193
rect 16187 179 16197 213
rect 16239 207 16249 241
rect 16283 207 16293 241
rect 16239 191 16293 207
rect 16095 163 16197 179
rect 16095 131 16125 163
rect 16244 131 16274 191
rect 16335 131 16365 299
rect 16711 333 16741 369
rect 16700 303 16741 333
rect 16492 265 16522 297
rect 16700 265 16730 303
rect 17007 491 17037 517
rect 17091 491 17121 517
rect 17358 497 17388 523
rect 17450 497 17480 523
rect 17549 497 17579 523
rect 17689 497 17719 523
rect 17786 497 17816 523
rect 17983 497 18013 523
rect 18082 497 18112 523
rect 18168 497 18198 523
rect 18252 497 18282 523
rect 18360 497 18390 523
rect 18444 497 18474 523
rect 18608 497 18638 523
rect 18827 497 18857 523
rect 18924 497 18954 523
rect 17007 348 17037 363
rect 16974 318 17037 348
rect 16808 265 16838 297
rect 16974 265 17004 318
rect 17091 274 17121 363
rect 17358 326 17388 413
rect 17450 375 17480 413
rect 16421 249 16730 265
rect 16421 215 16449 249
rect 16483 215 16730 249
rect 16421 199 16730 215
rect 16779 249 16838 265
rect 16779 215 16789 249
rect 16823 215 16838 249
rect 16779 199 16838 215
rect 16950 249 17004 265
rect 16950 215 16960 249
rect 16994 215 17004 249
rect 17046 264 17121 274
rect 17046 230 17062 264
rect 17096 230 17121 264
rect 17259 310 17388 326
rect 17434 365 17500 375
rect 17434 331 17450 365
rect 17484 331 17500 365
rect 17434 321 17500 331
rect 17259 276 17269 310
rect 17303 296 17388 310
rect 17303 276 17376 296
rect 17549 279 17579 413
rect 17689 355 17719 413
rect 17689 339 17744 355
rect 17689 305 17699 339
rect 17733 305 17744 339
rect 17689 289 17744 305
rect 17259 260 17376 276
rect 17046 220 17121 230
rect 16950 199 17004 215
rect 16523 177 16553 199
rect 16700 176 16730 199
rect 16808 177 16838 199
rect 16700 146 16741 176
rect 16711 131 16741 146
rect 16974 176 17004 199
rect 16974 146 17037 176
rect 17007 131 17037 146
rect 17091 131 17121 220
rect 17346 131 17376 260
rect 17441 249 17579 279
rect 17441 219 17472 249
rect 17418 203 17472 219
rect 17418 169 17428 203
rect 17462 169 17472 203
rect 17418 153 17472 169
rect 17514 197 17580 207
rect 17514 163 17530 197
rect 17564 163 17580 197
rect 17514 153 17580 163
rect 17441 119 17471 153
rect 17537 119 17567 153
rect 17703 131 17733 289
rect 17786 219 17816 413
rect 17983 314 18013 329
rect 17907 284 18013 314
rect 17907 267 17937 284
rect 17871 251 17937 267
rect 17775 203 17829 219
rect 17775 169 17785 203
rect 17819 169 17829 203
rect 17871 217 17881 251
rect 17915 217 17937 251
rect 18082 279 18112 413
rect 18168 381 18198 413
rect 18154 365 18208 381
rect 18154 331 18164 365
rect 18198 331 18208 365
rect 18154 315 18208 331
rect 18082 267 18132 279
rect 18082 255 18145 267
rect 18082 249 18169 255
rect 18103 239 18169 249
rect 18103 237 18125 239
rect 17871 201 17937 217
rect 17907 175 17937 201
rect 18006 191 18073 207
rect 17775 153 17829 169
rect 17775 131 17805 153
rect 18006 157 18029 191
rect 18063 157 18073 191
rect 18006 141 18073 157
rect 18115 205 18125 237
rect 18159 205 18169 239
rect 18115 189 18169 205
rect 18252 229 18282 413
rect 18360 257 18390 413
rect 18444 365 18474 413
rect 18432 349 18486 365
rect 18432 315 18442 349
rect 18476 315 18486 349
rect 18432 299 18486 315
rect 18355 241 18409 257
rect 18252 213 18313 229
rect 18252 193 18269 213
rect 18006 119 18036 141
rect 18115 119 18145 189
rect 18211 179 18269 193
rect 18303 179 18313 213
rect 18355 207 18365 241
rect 18399 207 18409 241
rect 18355 191 18409 207
rect 18211 163 18313 179
rect 18211 131 18241 163
rect 18360 131 18390 191
rect 18451 131 18481 299
rect 18827 333 18857 369
rect 18816 303 18857 333
rect 18608 265 18638 297
rect 18816 265 18846 303
rect 19123 491 19153 517
rect 19207 491 19237 517
rect 19474 497 19504 523
rect 19566 497 19596 523
rect 19665 497 19695 523
rect 19805 497 19835 523
rect 19902 497 19932 523
rect 20099 497 20129 523
rect 20198 497 20228 523
rect 20284 497 20314 523
rect 20368 497 20398 523
rect 20476 497 20506 523
rect 20560 497 20590 523
rect 20724 497 20754 523
rect 20943 497 20973 523
rect 21040 497 21070 523
rect 19123 348 19153 363
rect 19090 318 19153 348
rect 18924 265 18954 297
rect 19090 265 19120 318
rect 19207 274 19237 363
rect 19474 326 19504 413
rect 19566 375 19596 413
rect 18537 249 18846 265
rect 18537 215 18565 249
rect 18599 215 18846 249
rect 18537 199 18846 215
rect 18895 249 18954 265
rect 18895 215 18905 249
rect 18939 215 18954 249
rect 18895 199 18954 215
rect 19066 249 19120 265
rect 19066 215 19076 249
rect 19110 215 19120 249
rect 19162 264 19237 274
rect 19162 230 19178 264
rect 19212 230 19237 264
rect 19375 310 19504 326
rect 19550 365 19616 375
rect 19550 331 19566 365
rect 19600 331 19616 365
rect 19550 321 19616 331
rect 19375 276 19385 310
rect 19419 296 19504 310
rect 19419 276 19492 296
rect 19665 279 19695 413
rect 19805 355 19835 413
rect 19805 339 19860 355
rect 19805 305 19815 339
rect 19849 305 19860 339
rect 19805 289 19860 305
rect 19375 260 19492 276
rect 19162 220 19237 230
rect 19066 199 19120 215
rect 18639 177 18669 199
rect 18816 176 18846 199
rect 18924 177 18954 199
rect 18816 146 18857 176
rect 18827 131 18857 146
rect 19090 176 19120 199
rect 19090 146 19153 176
rect 19123 131 19153 146
rect 19207 131 19237 220
rect 19462 131 19492 260
rect 19557 249 19695 279
rect 19557 219 19588 249
rect 19534 203 19588 219
rect 19534 169 19544 203
rect 19578 169 19588 203
rect 19534 153 19588 169
rect 19630 197 19696 207
rect 19630 163 19646 197
rect 19680 163 19696 197
rect 19630 153 19696 163
rect 19557 119 19587 153
rect 19653 119 19683 153
rect 19819 131 19849 289
rect 19902 219 19932 413
rect 20099 314 20129 329
rect 20023 284 20129 314
rect 20023 267 20053 284
rect 19987 251 20053 267
rect 19891 203 19945 219
rect 19891 169 19901 203
rect 19935 169 19945 203
rect 19987 217 19997 251
rect 20031 217 20053 251
rect 20198 279 20228 413
rect 20284 381 20314 413
rect 20270 365 20324 381
rect 20270 331 20280 365
rect 20314 331 20324 365
rect 20270 315 20324 331
rect 20198 267 20248 279
rect 20198 255 20261 267
rect 20198 249 20285 255
rect 20219 239 20285 249
rect 20219 237 20241 239
rect 19987 201 20053 217
rect 20023 175 20053 201
rect 20122 191 20189 207
rect 19891 153 19945 169
rect 19891 131 19921 153
rect 20122 157 20145 191
rect 20179 157 20189 191
rect 20122 141 20189 157
rect 20231 205 20241 237
rect 20275 205 20285 239
rect 20231 189 20285 205
rect 20368 229 20398 413
rect 20476 257 20506 413
rect 20560 365 20590 413
rect 20548 349 20602 365
rect 20548 315 20558 349
rect 20592 315 20602 349
rect 20548 299 20602 315
rect 20471 241 20525 257
rect 20368 213 20429 229
rect 20368 193 20385 213
rect 20122 119 20152 141
rect 20231 119 20261 189
rect 20327 179 20385 193
rect 20419 179 20429 213
rect 20471 207 20481 241
rect 20515 207 20525 241
rect 20471 191 20525 207
rect 20327 163 20429 179
rect 20327 131 20357 163
rect 20476 131 20506 191
rect 20567 131 20597 299
rect 20943 333 20973 369
rect 20932 303 20973 333
rect 20724 265 20754 297
rect 20932 265 20962 303
rect 21239 491 21269 517
rect 21323 491 21353 517
rect 21590 497 21620 523
rect 21682 497 21712 523
rect 21781 497 21811 523
rect 21921 497 21951 523
rect 22018 497 22048 523
rect 22215 497 22245 523
rect 22314 497 22344 523
rect 22400 497 22430 523
rect 22484 497 22514 523
rect 22592 497 22622 523
rect 22676 497 22706 523
rect 22840 497 22870 523
rect 23059 497 23089 523
rect 23156 497 23186 523
rect 21239 348 21269 363
rect 21206 318 21269 348
rect 21040 265 21070 297
rect 21206 265 21236 318
rect 21323 274 21353 363
rect 21590 326 21620 413
rect 21682 375 21712 413
rect 20653 249 20962 265
rect 20653 215 20681 249
rect 20715 215 20962 249
rect 20653 199 20962 215
rect 21011 249 21070 265
rect 21011 215 21021 249
rect 21055 215 21070 249
rect 21011 199 21070 215
rect 21182 249 21236 265
rect 21182 215 21192 249
rect 21226 215 21236 249
rect 21278 264 21353 274
rect 21278 230 21294 264
rect 21328 230 21353 264
rect 21491 310 21620 326
rect 21666 365 21732 375
rect 21666 331 21682 365
rect 21716 331 21732 365
rect 21666 321 21732 331
rect 21491 276 21501 310
rect 21535 296 21620 310
rect 21535 276 21608 296
rect 21781 279 21811 413
rect 21921 355 21951 413
rect 21921 339 21976 355
rect 21921 305 21931 339
rect 21965 305 21976 339
rect 21921 289 21976 305
rect 21491 260 21608 276
rect 21278 220 21353 230
rect 21182 199 21236 215
rect 20755 177 20785 199
rect 20932 176 20962 199
rect 21040 177 21070 199
rect 20932 146 20973 176
rect 20943 131 20973 146
rect 21206 176 21236 199
rect 21206 146 21269 176
rect 21239 131 21269 146
rect 21323 131 21353 220
rect 21578 131 21608 260
rect 21673 249 21811 279
rect 21673 219 21704 249
rect 21650 203 21704 219
rect 21650 169 21660 203
rect 21694 169 21704 203
rect 21650 153 21704 169
rect 21746 197 21812 207
rect 21746 163 21762 197
rect 21796 163 21812 197
rect 21746 153 21812 163
rect 21673 119 21703 153
rect 21769 119 21799 153
rect 21935 131 21965 289
rect 22018 219 22048 413
rect 22215 314 22245 329
rect 22139 284 22245 314
rect 22139 267 22169 284
rect 22103 251 22169 267
rect 22007 203 22061 219
rect 22007 169 22017 203
rect 22051 169 22061 203
rect 22103 217 22113 251
rect 22147 217 22169 251
rect 22314 279 22344 413
rect 22400 381 22430 413
rect 22386 365 22440 381
rect 22386 331 22396 365
rect 22430 331 22440 365
rect 22386 315 22440 331
rect 22314 267 22364 279
rect 22314 255 22377 267
rect 22314 249 22401 255
rect 22335 239 22401 249
rect 22335 237 22357 239
rect 22103 201 22169 217
rect 22139 175 22169 201
rect 22238 191 22305 207
rect 22007 153 22061 169
rect 22007 131 22037 153
rect 22238 157 22261 191
rect 22295 157 22305 191
rect 22238 141 22305 157
rect 22347 205 22357 237
rect 22391 205 22401 239
rect 22347 189 22401 205
rect 22484 229 22514 413
rect 22592 257 22622 413
rect 22676 365 22706 413
rect 22664 349 22718 365
rect 22664 315 22674 349
rect 22708 315 22718 349
rect 22664 299 22718 315
rect 22587 241 22641 257
rect 22484 213 22545 229
rect 22484 193 22501 213
rect 22238 119 22268 141
rect 22347 119 22377 189
rect 22443 179 22501 193
rect 22535 179 22545 213
rect 22587 207 22597 241
rect 22631 207 22641 241
rect 22587 191 22641 207
rect 22443 163 22545 179
rect 22443 131 22473 163
rect 22592 131 22622 191
rect 22683 131 22713 299
rect 23059 333 23089 369
rect 23048 303 23089 333
rect 22840 265 22870 297
rect 23048 265 23078 303
rect 23355 491 23385 517
rect 23439 491 23469 517
rect 23706 497 23736 523
rect 23798 497 23828 523
rect 23897 497 23927 523
rect 24037 497 24067 523
rect 24134 497 24164 523
rect 24331 497 24361 523
rect 24430 497 24460 523
rect 24516 497 24546 523
rect 24600 497 24630 523
rect 24708 497 24738 523
rect 24792 497 24822 523
rect 24956 497 24986 523
rect 25175 497 25205 523
rect 25272 497 25302 523
rect 23355 348 23385 363
rect 23322 318 23385 348
rect 23156 265 23186 297
rect 23322 265 23352 318
rect 23439 274 23469 363
rect 23706 326 23736 413
rect 23798 375 23828 413
rect 22769 249 23078 265
rect 22769 215 22797 249
rect 22831 215 23078 249
rect 22769 199 23078 215
rect 23127 249 23186 265
rect 23127 215 23137 249
rect 23171 215 23186 249
rect 23127 199 23186 215
rect 23298 249 23352 265
rect 23298 215 23308 249
rect 23342 215 23352 249
rect 23394 264 23469 274
rect 23394 230 23410 264
rect 23444 230 23469 264
rect 23607 310 23736 326
rect 23782 365 23848 375
rect 23782 331 23798 365
rect 23832 331 23848 365
rect 23782 321 23848 331
rect 23607 276 23617 310
rect 23651 296 23736 310
rect 23651 276 23724 296
rect 23897 279 23927 413
rect 24037 355 24067 413
rect 24037 339 24092 355
rect 24037 305 24047 339
rect 24081 305 24092 339
rect 24037 289 24092 305
rect 23607 260 23724 276
rect 23394 220 23469 230
rect 23298 199 23352 215
rect 22871 177 22901 199
rect 23048 176 23078 199
rect 23156 177 23186 199
rect 23048 146 23089 176
rect 23059 131 23089 146
rect 23322 176 23352 199
rect 23322 146 23385 176
rect 23355 131 23385 146
rect 23439 131 23469 220
rect 23694 131 23724 260
rect 23789 249 23927 279
rect 23789 219 23820 249
rect 23766 203 23820 219
rect 23766 169 23776 203
rect 23810 169 23820 203
rect 23766 153 23820 169
rect 23862 197 23928 207
rect 23862 163 23878 197
rect 23912 163 23928 197
rect 23862 153 23928 163
rect 23789 119 23819 153
rect 23885 119 23915 153
rect 24051 131 24081 289
rect 24134 219 24164 413
rect 24331 314 24361 329
rect 24255 284 24361 314
rect 24255 267 24285 284
rect 24219 251 24285 267
rect 24123 203 24177 219
rect 24123 169 24133 203
rect 24167 169 24177 203
rect 24219 217 24229 251
rect 24263 217 24285 251
rect 24430 279 24460 413
rect 24516 381 24546 413
rect 24502 365 24556 381
rect 24502 331 24512 365
rect 24546 331 24556 365
rect 24502 315 24556 331
rect 24430 267 24480 279
rect 24430 255 24493 267
rect 24430 249 24517 255
rect 24451 239 24517 249
rect 24451 237 24473 239
rect 24219 201 24285 217
rect 24255 175 24285 201
rect 24354 191 24421 207
rect 24123 153 24177 169
rect 24123 131 24153 153
rect 24354 157 24377 191
rect 24411 157 24421 191
rect 24354 141 24421 157
rect 24463 205 24473 237
rect 24507 205 24517 239
rect 24463 189 24517 205
rect 24600 229 24630 413
rect 24708 257 24738 413
rect 24792 365 24822 413
rect 24780 349 24834 365
rect 24780 315 24790 349
rect 24824 315 24834 349
rect 24780 299 24834 315
rect 24703 241 24757 257
rect 24600 213 24661 229
rect 24600 193 24617 213
rect 24354 119 24384 141
rect 24463 119 24493 189
rect 24559 179 24617 193
rect 24651 179 24661 213
rect 24703 207 24713 241
rect 24747 207 24757 241
rect 24703 191 24757 207
rect 24559 163 24661 179
rect 24559 131 24589 163
rect 24708 131 24738 191
rect 24799 131 24829 299
rect 25175 333 25205 369
rect 25164 303 25205 333
rect 24956 265 24986 297
rect 25164 265 25194 303
rect 25471 491 25501 517
rect 25555 491 25585 517
rect 25822 497 25852 523
rect 25914 497 25944 523
rect 26013 497 26043 523
rect 26153 497 26183 523
rect 26250 497 26280 523
rect 26447 497 26477 523
rect 26546 497 26576 523
rect 26632 497 26662 523
rect 26716 497 26746 523
rect 26824 497 26854 523
rect 26908 497 26938 523
rect 27072 497 27102 523
rect 27291 497 27321 523
rect 27388 497 27418 523
rect 25471 348 25501 363
rect 25438 318 25501 348
rect 25272 265 25302 297
rect 25438 265 25468 318
rect 25555 274 25585 363
rect 25822 326 25852 413
rect 25914 375 25944 413
rect 24885 249 25194 265
rect 24885 215 24913 249
rect 24947 215 25194 249
rect 24885 199 25194 215
rect 25243 249 25302 265
rect 25243 215 25253 249
rect 25287 215 25302 249
rect 25243 199 25302 215
rect 25414 249 25468 265
rect 25414 215 25424 249
rect 25458 215 25468 249
rect 25510 264 25585 274
rect 25510 230 25526 264
rect 25560 230 25585 264
rect 25723 310 25852 326
rect 25898 365 25964 375
rect 25898 331 25914 365
rect 25948 331 25964 365
rect 25898 321 25964 331
rect 25723 276 25733 310
rect 25767 296 25852 310
rect 25767 276 25840 296
rect 26013 279 26043 413
rect 26153 355 26183 413
rect 26153 339 26208 355
rect 26153 305 26163 339
rect 26197 305 26208 339
rect 26153 289 26208 305
rect 25723 260 25840 276
rect 25510 220 25585 230
rect 25414 199 25468 215
rect 24987 177 25017 199
rect 25164 176 25194 199
rect 25272 177 25302 199
rect 25164 146 25205 176
rect 25175 131 25205 146
rect 25438 176 25468 199
rect 25438 146 25501 176
rect 25471 131 25501 146
rect 25555 131 25585 220
rect 25810 131 25840 260
rect 25905 249 26043 279
rect 25905 219 25936 249
rect 25882 203 25936 219
rect 25882 169 25892 203
rect 25926 169 25936 203
rect 25882 153 25936 169
rect 25978 197 26044 207
rect 25978 163 25994 197
rect 26028 163 26044 197
rect 25978 153 26044 163
rect 25905 119 25935 153
rect 26001 119 26031 153
rect 26167 131 26197 289
rect 26250 219 26280 413
rect 26447 314 26477 329
rect 26371 284 26477 314
rect 26371 267 26401 284
rect 26335 251 26401 267
rect 26239 203 26293 219
rect 26239 169 26249 203
rect 26283 169 26293 203
rect 26335 217 26345 251
rect 26379 217 26401 251
rect 26546 279 26576 413
rect 26632 381 26662 413
rect 26618 365 26672 381
rect 26618 331 26628 365
rect 26662 331 26672 365
rect 26618 315 26672 331
rect 26546 267 26596 279
rect 26546 255 26609 267
rect 26546 249 26633 255
rect 26567 239 26633 249
rect 26567 237 26589 239
rect 26335 201 26401 217
rect 26371 175 26401 201
rect 26470 191 26537 207
rect 26239 153 26293 169
rect 26239 131 26269 153
rect 26470 157 26493 191
rect 26527 157 26537 191
rect 26470 141 26537 157
rect 26579 205 26589 237
rect 26623 205 26633 239
rect 26579 189 26633 205
rect 26716 229 26746 413
rect 26824 257 26854 413
rect 26908 365 26938 413
rect 26896 349 26950 365
rect 26896 315 26906 349
rect 26940 315 26950 349
rect 26896 299 26950 315
rect 26819 241 26873 257
rect 26716 213 26777 229
rect 26716 193 26733 213
rect 26470 119 26500 141
rect 26579 119 26609 189
rect 26675 179 26733 193
rect 26767 179 26777 213
rect 26819 207 26829 241
rect 26863 207 26873 241
rect 26819 191 26873 207
rect 26675 163 26777 179
rect 26675 131 26705 163
rect 26824 131 26854 191
rect 26915 131 26945 299
rect 27291 333 27321 369
rect 27280 303 27321 333
rect 27072 265 27102 297
rect 27280 265 27310 303
rect 27587 491 27617 517
rect 27671 491 27701 517
rect 27938 497 27968 523
rect 28030 497 28060 523
rect 28129 497 28159 523
rect 28269 497 28299 523
rect 28366 497 28396 523
rect 28563 497 28593 523
rect 28662 497 28692 523
rect 28748 497 28778 523
rect 28832 497 28862 523
rect 28940 497 28970 523
rect 29024 497 29054 523
rect 29188 497 29218 523
rect 29407 497 29437 523
rect 29504 497 29534 523
rect 27587 348 27617 363
rect 27554 318 27617 348
rect 27388 265 27418 297
rect 27554 265 27584 318
rect 27671 274 27701 363
rect 27938 326 27968 413
rect 28030 375 28060 413
rect 27001 249 27310 265
rect 27001 215 27029 249
rect 27063 215 27310 249
rect 27001 199 27310 215
rect 27359 249 27418 265
rect 27359 215 27369 249
rect 27403 215 27418 249
rect 27359 199 27418 215
rect 27530 249 27584 265
rect 27530 215 27540 249
rect 27574 215 27584 249
rect 27626 264 27701 274
rect 27626 230 27642 264
rect 27676 230 27701 264
rect 27839 310 27968 326
rect 28014 365 28080 375
rect 28014 331 28030 365
rect 28064 331 28080 365
rect 28014 321 28080 331
rect 27839 276 27849 310
rect 27883 296 27968 310
rect 27883 276 27956 296
rect 28129 279 28159 413
rect 28269 355 28299 413
rect 28269 339 28324 355
rect 28269 305 28279 339
rect 28313 305 28324 339
rect 28269 289 28324 305
rect 27839 260 27956 276
rect 27626 220 27701 230
rect 27530 199 27584 215
rect 27103 177 27133 199
rect 27280 176 27310 199
rect 27388 177 27418 199
rect 27280 146 27321 176
rect 27291 131 27321 146
rect 27554 176 27584 199
rect 27554 146 27617 176
rect 27587 131 27617 146
rect 27671 131 27701 220
rect 27926 131 27956 260
rect 28021 249 28159 279
rect 28021 219 28052 249
rect 27998 203 28052 219
rect 27998 169 28008 203
rect 28042 169 28052 203
rect 27998 153 28052 169
rect 28094 197 28160 207
rect 28094 163 28110 197
rect 28144 163 28160 197
rect 28094 153 28160 163
rect 28021 119 28051 153
rect 28117 119 28147 153
rect 28283 131 28313 289
rect 28366 219 28396 413
rect 28563 314 28593 329
rect 28487 284 28593 314
rect 28487 267 28517 284
rect 28451 251 28517 267
rect 28355 203 28409 219
rect 28355 169 28365 203
rect 28399 169 28409 203
rect 28451 217 28461 251
rect 28495 217 28517 251
rect 28662 279 28692 413
rect 28748 381 28778 413
rect 28734 365 28788 381
rect 28734 331 28744 365
rect 28778 331 28788 365
rect 28734 315 28788 331
rect 28662 267 28712 279
rect 28662 255 28725 267
rect 28662 249 28749 255
rect 28683 239 28749 249
rect 28683 237 28705 239
rect 28451 201 28517 217
rect 28487 175 28517 201
rect 28586 191 28653 207
rect 28355 153 28409 169
rect 28355 131 28385 153
rect 28586 157 28609 191
rect 28643 157 28653 191
rect 28586 141 28653 157
rect 28695 205 28705 237
rect 28739 205 28749 239
rect 28695 189 28749 205
rect 28832 229 28862 413
rect 28940 257 28970 413
rect 29024 365 29054 413
rect 29012 349 29066 365
rect 29012 315 29022 349
rect 29056 315 29066 349
rect 29012 299 29066 315
rect 28935 241 28989 257
rect 28832 213 28893 229
rect 28832 193 28849 213
rect 28586 119 28616 141
rect 28695 119 28725 189
rect 28791 179 28849 193
rect 28883 179 28893 213
rect 28935 207 28945 241
rect 28979 207 28989 241
rect 28935 191 28989 207
rect 28791 163 28893 179
rect 28791 131 28821 163
rect 28940 131 28970 191
rect 29031 131 29061 299
rect 29407 333 29437 369
rect 29396 303 29437 333
rect 29188 265 29218 297
rect 29396 265 29426 303
rect 29703 491 29733 517
rect 29787 491 29817 517
rect 30054 497 30084 523
rect 30146 497 30176 523
rect 30245 497 30275 523
rect 30385 497 30415 523
rect 30482 497 30512 523
rect 30679 497 30709 523
rect 30778 497 30808 523
rect 30864 497 30894 523
rect 30948 497 30978 523
rect 31056 497 31086 523
rect 31140 497 31170 523
rect 31304 497 31334 523
rect 31523 497 31553 523
rect 31620 497 31650 523
rect 29703 348 29733 363
rect 29670 318 29733 348
rect 29504 265 29534 297
rect 29670 265 29700 318
rect 29787 274 29817 363
rect 30054 326 30084 413
rect 30146 375 30176 413
rect 29117 249 29426 265
rect 29117 215 29145 249
rect 29179 215 29426 249
rect 29117 199 29426 215
rect 29475 249 29534 265
rect 29475 215 29485 249
rect 29519 215 29534 249
rect 29475 199 29534 215
rect 29646 249 29700 265
rect 29646 215 29656 249
rect 29690 215 29700 249
rect 29742 264 29817 274
rect 29742 230 29758 264
rect 29792 230 29817 264
rect 29955 310 30084 326
rect 30130 365 30196 375
rect 30130 331 30146 365
rect 30180 331 30196 365
rect 30130 321 30196 331
rect 29955 276 29965 310
rect 29999 296 30084 310
rect 29999 276 30072 296
rect 30245 279 30275 413
rect 30385 355 30415 413
rect 30385 339 30440 355
rect 30385 305 30395 339
rect 30429 305 30440 339
rect 30385 289 30440 305
rect 29955 260 30072 276
rect 29742 220 29817 230
rect 29646 199 29700 215
rect 29219 177 29249 199
rect 29396 176 29426 199
rect 29504 177 29534 199
rect 29396 146 29437 176
rect 29407 131 29437 146
rect 29670 176 29700 199
rect 29670 146 29733 176
rect 29703 131 29733 146
rect 29787 131 29817 220
rect 30042 131 30072 260
rect 30137 249 30275 279
rect 30137 219 30168 249
rect 30114 203 30168 219
rect 30114 169 30124 203
rect 30158 169 30168 203
rect 30114 153 30168 169
rect 30210 197 30276 207
rect 30210 163 30226 197
rect 30260 163 30276 197
rect 30210 153 30276 163
rect 30137 119 30167 153
rect 30233 119 30263 153
rect 30399 131 30429 289
rect 30482 219 30512 413
rect 30679 314 30709 329
rect 30603 284 30709 314
rect 30603 267 30633 284
rect 30567 251 30633 267
rect 30471 203 30525 219
rect 30471 169 30481 203
rect 30515 169 30525 203
rect 30567 217 30577 251
rect 30611 217 30633 251
rect 30778 279 30808 413
rect 30864 381 30894 413
rect 30850 365 30904 381
rect 30850 331 30860 365
rect 30894 331 30904 365
rect 30850 315 30904 331
rect 30778 267 30828 279
rect 30778 255 30841 267
rect 30778 249 30865 255
rect 30799 239 30865 249
rect 30799 237 30821 239
rect 30567 201 30633 217
rect 30603 175 30633 201
rect 30702 191 30769 207
rect 30471 153 30525 169
rect 30471 131 30501 153
rect 30702 157 30725 191
rect 30759 157 30769 191
rect 30702 141 30769 157
rect 30811 205 30821 237
rect 30855 205 30865 239
rect 30811 189 30865 205
rect 30948 229 30978 413
rect 31056 257 31086 413
rect 31140 365 31170 413
rect 31128 349 31182 365
rect 31128 315 31138 349
rect 31172 315 31182 349
rect 31128 299 31182 315
rect 31051 241 31105 257
rect 30948 213 31009 229
rect 30948 193 30965 213
rect 30702 119 30732 141
rect 30811 119 30841 189
rect 30907 179 30965 193
rect 30999 179 31009 213
rect 31051 207 31061 241
rect 31095 207 31105 241
rect 31051 191 31105 207
rect 30907 163 31009 179
rect 30907 131 30937 163
rect 31056 131 31086 191
rect 31147 131 31177 299
rect 31523 333 31553 369
rect 31512 303 31553 333
rect 31304 265 31334 297
rect 31512 265 31542 303
rect 31819 491 31849 517
rect 31903 491 31933 517
rect 32170 497 32200 523
rect 32262 497 32292 523
rect 32361 497 32391 523
rect 32501 497 32531 523
rect 32598 497 32628 523
rect 32795 497 32825 523
rect 32894 497 32924 523
rect 32980 497 33010 523
rect 33064 497 33094 523
rect 33172 497 33202 523
rect 33256 497 33286 523
rect 33420 497 33450 523
rect 33639 497 33669 523
rect 33736 497 33766 523
rect 31819 348 31849 363
rect 31786 318 31849 348
rect 31620 265 31650 297
rect 31786 265 31816 318
rect 31903 274 31933 363
rect 32170 326 32200 413
rect 32262 375 32292 413
rect 31233 249 31542 265
rect 31233 215 31261 249
rect 31295 215 31542 249
rect 31233 199 31542 215
rect 31591 249 31650 265
rect 31591 215 31601 249
rect 31635 215 31650 249
rect 31591 199 31650 215
rect 31762 249 31816 265
rect 31762 215 31772 249
rect 31806 215 31816 249
rect 31858 264 31933 274
rect 31858 230 31874 264
rect 31908 230 31933 264
rect 32071 310 32200 326
rect 32246 365 32312 375
rect 32246 331 32262 365
rect 32296 331 32312 365
rect 32246 321 32312 331
rect 32071 276 32081 310
rect 32115 296 32200 310
rect 32115 276 32188 296
rect 32361 279 32391 413
rect 32501 355 32531 413
rect 32501 339 32556 355
rect 32501 305 32511 339
rect 32545 305 32556 339
rect 32501 289 32556 305
rect 32071 260 32188 276
rect 31858 220 31933 230
rect 31762 199 31816 215
rect 31335 177 31365 199
rect 31512 176 31542 199
rect 31620 177 31650 199
rect 31512 146 31553 176
rect 31523 131 31553 146
rect 31786 176 31816 199
rect 31786 146 31849 176
rect 31819 131 31849 146
rect 31903 131 31933 220
rect 32158 131 32188 260
rect 32253 249 32391 279
rect 32253 219 32284 249
rect 32230 203 32284 219
rect 32230 169 32240 203
rect 32274 169 32284 203
rect 32230 153 32284 169
rect 32326 197 32392 207
rect 32326 163 32342 197
rect 32376 163 32392 197
rect 32326 153 32392 163
rect 32253 119 32283 153
rect 32349 119 32379 153
rect 32515 131 32545 289
rect 32598 219 32628 413
rect 32795 314 32825 329
rect 32719 284 32825 314
rect 32719 267 32749 284
rect 32683 251 32749 267
rect 32587 203 32641 219
rect 32587 169 32597 203
rect 32631 169 32641 203
rect 32683 217 32693 251
rect 32727 217 32749 251
rect 32894 279 32924 413
rect 32980 381 33010 413
rect 32966 365 33020 381
rect 32966 331 32976 365
rect 33010 331 33020 365
rect 32966 315 33020 331
rect 32894 267 32944 279
rect 32894 255 32957 267
rect 32894 249 32981 255
rect 32915 239 32981 249
rect 32915 237 32937 239
rect 32683 201 32749 217
rect 32719 175 32749 201
rect 32818 191 32885 207
rect 32587 153 32641 169
rect 32587 131 32617 153
rect 32818 157 32841 191
rect 32875 157 32885 191
rect 32818 141 32885 157
rect 32927 205 32937 237
rect 32971 205 32981 239
rect 32927 189 32981 205
rect 33064 229 33094 413
rect 33172 257 33202 413
rect 33256 365 33286 413
rect 33244 349 33298 365
rect 33244 315 33254 349
rect 33288 315 33298 349
rect 33244 299 33298 315
rect 33167 241 33221 257
rect 33064 213 33125 229
rect 33064 193 33081 213
rect 32818 119 32848 141
rect 32927 119 32957 189
rect 33023 179 33081 193
rect 33115 179 33125 213
rect 33167 207 33177 241
rect 33211 207 33221 241
rect 33167 191 33221 207
rect 33023 163 33125 179
rect 33023 131 33053 163
rect 33172 131 33202 191
rect 33263 131 33293 299
rect 33639 333 33669 369
rect 33628 303 33669 333
rect 33420 265 33450 297
rect 33628 265 33658 303
rect 33935 491 33965 517
rect 34019 491 34049 517
rect 34286 497 34316 523
rect 34378 497 34408 523
rect 34477 497 34507 523
rect 34617 497 34647 523
rect 34714 497 34744 523
rect 34911 497 34941 523
rect 35010 497 35040 523
rect 35096 497 35126 523
rect 35180 497 35210 523
rect 35288 497 35318 523
rect 35372 497 35402 523
rect 35536 497 35566 523
rect 35755 497 35785 523
rect 35852 497 35882 523
rect 33935 348 33965 363
rect 33902 318 33965 348
rect 33736 265 33766 297
rect 33902 265 33932 318
rect 34019 274 34049 363
rect 34286 326 34316 413
rect 34378 375 34408 413
rect 33349 249 33658 265
rect 33349 215 33377 249
rect 33411 215 33658 249
rect 33349 199 33658 215
rect 33707 249 33766 265
rect 33707 215 33717 249
rect 33751 215 33766 249
rect 33707 199 33766 215
rect 33878 249 33932 265
rect 33878 215 33888 249
rect 33922 215 33932 249
rect 33974 264 34049 274
rect 33974 230 33990 264
rect 34024 230 34049 264
rect 34187 310 34316 326
rect 34362 365 34428 375
rect 34362 331 34378 365
rect 34412 331 34428 365
rect 34362 321 34428 331
rect 34187 276 34197 310
rect 34231 296 34316 310
rect 34231 276 34304 296
rect 34477 279 34507 413
rect 34617 355 34647 413
rect 34617 339 34672 355
rect 34617 305 34627 339
rect 34661 305 34672 339
rect 34617 289 34672 305
rect 34187 260 34304 276
rect 33974 220 34049 230
rect 33878 199 33932 215
rect 33451 177 33481 199
rect 33628 176 33658 199
rect 33736 177 33766 199
rect 33628 146 33669 176
rect 33639 131 33669 146
rect 33902 176 33932 199
rect 33902 146 33965 176
rect 33935 131 33965 146
rect 34019 131 34049 220
rect 34274 131 34304 260
rect 34369 249 34507 279
rect 34369 219 34400 249
rect 34346 203 34400 219
rect 34346 169 34356 203
rect 34390 169 34400 203
rect 34346 153 34400 169
rect 34442 197 34508 207
rect 34442 163 34458 197
rect 34492 163 34508 197
rect 34442 153 34508 163
rect 34369 119 34399 153
rect 34465 119 34495 153
rect 34631 131 34661 289
rect 34714 219 34744 413
rect 34911 314 34941 329
rect 34835 284 34941 314
rect 34835 267 34865 284
rect 34799 251 34865 267
rect 34703 203 34757 219
rect 34703 169 34713 203
rect 34747 169 34757 203
rect 34799 217 34809 251
rect 34843 217 34865 251
rect 35010 279 35040 413
rect 35096 381 35126 413
rect 35082 365 35136 381
rect 35082 331 35092 365
rect 35126 331 35136 365
rect 35082 315 35136 331
rect 35010 267 35060 279
rect 35010 255 35073 267
rect 35010 249 35097 255
rect 35031 239 35097 249
rect 35031 237 35053 239
rect 34799 201 34865 217
rect 34835 175 34865 201
rect 34934 191 35001 207
rect 34703 153 34757 169
rect 34703 131 34733 153
rect 34934 157 34957 191
rect 34991 157 35001 191
rect 34934 141 35001 157
rect 35043 205 35053 237
rect 35087 205 35097 239
rect 35043 189 35097 205
rect 35180 229 35210 413
rect 35288 257 35318 413
rect 35372 365 35402 413
rect 35360 349 35414 365
rect 35360 315 35370 349
rect 35404 315 35414 349
rect 35360 299 35414 315
rect 35283 241 35337 257
rect 35180 213 35241 229
rect 35180 193 35197 213
rect 34934 119 34964 141
rect 35043 119 35073 189
rect 35139 179 35197 193
rect 35231 179 35241 213
rect 35283 207 35293 241
rect 35327 207 35337 241
rect 35283 191 35337 207
rect 35139 163 35241 179
rect 35139 131 35169 163
rect 35288 131 35318 191
rect 35379 131 35409 299
rect 35755 333 35785 369
rect 35744 303 35785 333
rect 35536 265 35566 297
rect 35744 265 35774 303
rect 36051 491 36081 517
rect 36135 491 36165 517
rect 36402 497 36432 523
rect 36494 497 36524 523
rect 36593 497 36623 523
rect 36733 497 36763 523
rect 36830 497 36860 523
rect 37027 497 37057 523
rect 37126 497 37156 523
rect 37212 497 37242 523
rect 37296 497 37326 523
rect 37404 497 37434 523
rect 37488 497 37518 523
rect 37652 497 37682 523
rect 37871 497 37901 523
rect 37968 497 37998 523
rect 36051 348 36081 363
rect 36018 318 36081 348
rect 35852 265 35882 297
rect 36018 265 36048 318
rect 36135 274 36165 363
rect 36402 326 36432 413
rect 36494 375 36524 413
rect 35465 249 35774 265
rect 35465 215 35493 249
rect 35527 215 35774 249
rect 35465 199 35774 215
rect 35823 249 35882 265
rect 35823 215 35833 249
rect 35867 215 35882 249
rect 35823 199 35882 215
rect 35994 249 36048 265
rect 35994 215 36004 249
rect 36038 215 36048 249
rect 36090 264 36165 274
rect 36090 230 36106 264
rect 36140 230 36165 264
rect 36303 310 36432 326
rect 36478 365 36544 375
rect 36478 331 36494 365
rect 36528 331 36544 365
rect 36478 321 36544 331
rect 36303 276 36313 310
rect 36347 296 36432 310
rect 36347 276 36420 296
rect 36593 279 36623 413
rect 36733 355 36763 413
rect 36733 339 36788 355
rect 36733 305 36743 339
rect 36777 305 36788 339
rect 36733 289 36788 305
rect 36303 260 36420 276
rect 36090 220 36165 230
rect 35994 199 36048 215
rect 35567 177 35597 199
rect 35744 176 35774 199
rect 35852 177 35882 199
rect 35744 146 35785 176
rect 35755 131 35785 146
rect 36018 176 36048 199
rect 36018 146 36081 176
rect 36051 131 36081 146
rect 36135 131 36165 220
rect 36390 131 36420 260
rect 36485 249 36623 279
rect 36485 219 36516 249
rect 36462 203 36516 219
rect 36462 169 36472 203
rect 36506 169 36516 203
rect 36462 153 36516 169
rect 36558 197 36624 207
rect 36558 163 36574 197
rect 36608 163 36624 197
rect 36558 153 36624 163
rect 36485 119 36515 153
rect 36581 119 36611 153
rect 36747 131 36777 289
rect 36830 219 36860 413
rect 37027 314 37057 329
rect 36951 284 37057 314
rect 36951 267 36981 284
rect 36915 251 36981 267
rect 36819 203 36873 219
rect 36819 169 36829 203
rect 36863 169 36873 203
rect 36915 217 36925 251
rect 36959 217 36981 251
rect 37126 279 37156 413
rect 37212 381 37242 413
rect 37198 365 37252 381
rect 37198 331 37208 365
rect 37242 331 37252 365
rect 37198 315 37252 331
rect 37126 267 37176 279
rect 37126 255 37189 267
rect 37126 249 37213 255
rect 37147 239 37213 249
rect 37147 237 37169 239
rect 36915 201 36981 217
rect 36951 175 36981 201
rect 37050 191 37117 207
rect 36819 153 36873 169
rect 36819 131 36849 153
rect 37050 157 37073 191
rect 37107 157 37117 191
rect 37050 141 37117 157
rect 37159 205 37169 237
rect 37203 205 37213 239
rect 37159 189 37213 205
rect 37296 229 37326 413
rect 37404 257 37434 413
rect 37488 365 37518 413
rect 37476 349 37530 365
rect 37476 315 37486 349
rect 37520 315 37530 349
rect 37476 299 37530 315
rect 37399 241 37453 257
rect 37296 213 37357 229
rect 37296 193 37313 213
rect 37050 119 37080 141
rect 37159 119 37189 189
rect 37255 179 37313 193
rect 37347 179 37357 213
rect 37399 207 37409 241
rect 37443 207 37453 241
rect 37399 191 37453 207
rect 37255 163 37357 179
rect 37255 131 37285 163
rect 37404 131 37434 191
rect 37495 131 37525 299
rect 37871 333 37901 369
rect 37860 303 37901 333
rect 37652 265 37682 297
rect 37860 265 37890 303
rect 38167 491 38197 517
rect 38251 491 38281 517
rect 38518 497 38548 523
rect 38610 497 38640 523
rect 38709 497 38739 523
rect 38849 497 38879 523
rect 38946 497 38976 523
rect 39143 497 39173 523
rect 39242 497 39272 523
rect 39328 497 39358 523
rect 39412 497 39442 523
rect 39520 497 39550 523
rect 39604 497 39634 523
rect 39768 497 39798 523
rect 39987 497 40017 523
rect 40084 497 40114 523
rect 38167 348 38197 363
rect 38134 318 38197 348
rect 37968 265 37998 297
rect 38134 265 38164 318
rect 38251 274 38281 363
rect 38518 326 38548 413
rect 38610 375 38640 413
rect 37581 249 37890 265
rect 37581 215 37609 249
rect 37643 215 37890 249
rect 37581 199 37890 215
rect 37939 249 37998 265
rect 37939 215 37949 249
rect 37983 215 37998 249
rect 37939 199 37998 215
rect 38110 249 38164 265
rect 38110 215 38120 249
rect 38154 215 38164 249
rect 38206 264 38281 274
rect 38206 230 38222 264
rect 38256 230 38281 264
rect 38419 310 38548 326
rect 38594 365 38660 375
rect 38594 331 38610 365
rect 38644 331 38660 365
rect 38594 321 38660 331
rect 38419 276 38429 310
rect 38463 296 38548 310
rect 38463 276 38536 296
rect 38709 279 38739 413
rect 38849 355 38879 413
rect 38849 339 38904 355
rect 38849 305 38859 339
rect 38893 305 38904 339
rect 38849 289 38904 305
rect 38419 260 38536 276
rect 38206 220 38281 230
rect 38110 199 38164 215
rect 37683 177 37713 199
rect 37860 176 37890 199
rect 37968 177 37998 199
rect 37860 146 37901 176
rect 37871 131 37901 146
rect 38134 176 38164 199
rect 38134 146 38197 176
rect 38167 131 38197 146
rect 38251 131 38281 220
rect 38506 131 38536 260
rect 38601 249 38739 279
rect 38601 219 38632 249
rect 38578 203 38632 219
rect 38578 169 38588 203
rect 38622 169 38632 203
rect 38578 153 38632 169
rect 38674 197 38740 207
rect 38674 163 38690 197
rect 38724 163 38740 197
rect 38674 153 38740 163
rect 38601 119 38631 153
rect 38697 119 38727 153
rect 38863 131 38893 289
rect 38946 219 38976 413
rect 39143 314 39173 329
rect 39067 284 39173 314
rect 39067 267 39097 284
rect 39031 251 39097 267
rect 38935 203 38989 219
rect 38935 169 38945 203
rect 38979 169 38989 203
rect 39031 217 39041 251
rect 39075 217 39097 251
rect 39242 279 39272 413
rect 39328 381 39358 413
rect 39314 365 39368 381
rect 39314 331 39324 365
rect 39358 331 39368 365
rect 39314 315 39368 331
rect 39242 267 39292 279
rect 39242 255 39305 267
rect 39242 249 39329 255
rect 39263 239 39329 249
rect 39263 237 39285 239
rect 39031 201 39097 217
rect 39067 175 39097 201
rect 39166 191 39233 207
rect 38935 153 38989 169
rect 38935 131 38965 153
rect 39166 157 39189 191
rect 39223 157 39233 191
rect 39166 141 39233 157
rect 39275 205 39285 237
rect 39319 205 39329 239
rect 39275 189 39329 205
rect 39412 229 39442 413
rect 39520 257 39550 413
rect 39604 365 39634 413
rect 39592 349 39646 365
rect 39592 315 39602 349
rect 39636 315 39646 349
rect 39592 299 39646 315
rect 39515 241 39569 257
rect 39412 213 39473 229
rect 39412 193 39429 213
rect 39166 119 39196 141
rect 39275 119 39305 189
rect 39371 179 39429 193
rect 39463 179 39473 213
rect 39515 207 39525 241
rect 39559 207 39569 241
rect 39515 191 39569 207
rect 39371 163 39473 179
rect 39371 131 39401 163
rect 39520 131 39550 191
rect 39611 131 39641 299
rect 39987 333 40017 369
rect 39976 303 40017 333
rect 39768 265 39798 297
rect 39976 265 40006 303
rect 40283 491 40313 517
rect 40367 491 40397 517
rect 40634 497 40664 523
rect 40726 497 40756 523
rect 40825 497 40855 523
rect 40965 497 40995 523
rect 41062 497 41092 523
rect 41259 497 41289 523
rect 41358 497 41388 523
rect 41444 497 41474 523
rect 41528 497 41558 523
rect 41636 497 41666 523
rect 41720 497 41750 523
rect 41884 497 41914 523
rect 42103 497 42133 523
rect 42200 497 42230 523
rect 40283 348 40313 363
rect 40250 318 40313 348
rect 40084 265 40114 297
rect 40250 265 40280 318
rect 40367 274 40397 363
rect 40634 326 40664 413
rect 40726 375 40756 413
rect 39697 249 40006 265
rect 39697 215 39725 249
rect 39759 215 40006 249
rect 39697 199 40006 215
rect 40055 249 40114 265
rect 40055 215 40065 249
rect 40099 215 40114 249
rect 40055 199 40114 215
rect 40226 249 40280 265
rect 40226 215 40236 249
rect 40270 215 40280 249
rect 40322 264 40397 274
rect 40322 230 40338 264
rect 40372 230 40397 264
rect 40535 310 40664 326
rect 40710 365 40776 375
rect 40710 331 40726 365
rect 40760 331 40776 365
rect 40710 321 40776 331
rect 40535 276 40545 310
rect 40579 296 40664 310
rect 40579 276 40652 296
rect 40825 279 40855 413
rect 40965 355 40995 413
rect 40965 339 41020 355
rect 40965 305 40975 339
rect 41009 305 41020 339
rect 40965 289 41020 305
rect 40535 260 40652 276
rect 40322 220 40397 230
rect 40226 199 40280 215
rect 39799 177 39829 199
rect 39976 176 40006 199
rect 40084 177 40114 199
rect 39976 146 40017 176
rect 39987 131 40017 146
rect 40250 176 40280 199
rect 40250 146 40313 176
rect 40283 131 40313 146
rect 40367 131 40397 220
rect 40622 131 40652 260
rect 40717 249 40855 279
rect 40717 219 40748 249
rect 40694 203 40748 219
rect 40694 169 40704 203
rect 40738 169 40748 203
rect 40694 153 40748 169
rect 40790 197 40856 207
rect 40790 163 40806 197
rect 40840 163 40856 197
rect 40790 153 40856 163
rect 40717 119 40747 153
rect 40813 119 40843 153
rect 40979 131 41009 289
rect 41062 219 41092 413
rect 41259 314 41289 329
rect 41183 284 41289 314
rect 41183 267 41213 284
rect 41147 251 41213 267
rect 41051 203 41105 219
rect 41051 169 41061 203
rect 41095 169 41105 203
rect 41147 217 41157 251
rect 41191 217 41213 251
rect 41358 279 41388 413
rect 41444 381 41474 413
rect 41430 365 41484 381
rect 41430 331 41440 365
rect 41474 331 41484 365
rect 41430 315 41484 331
rect 41358 267 41408 279
rect 41358 255 41421 267
rect 41358 249 41445 255
rect 41379 239 41445 249
rect 41379 237 41401 239
rect 41147 201 41213 217
rect 41183 175 41213 201
rect 41282 191 41349 207
rect 41051 153 41105 169
rect 41051 131 41081 153
rect 41282 157 41305 191
rect 41339 157 41349 191
rect 41282 141 41349 157
rect 41391 205 41401 237
rect 41435 205 41445 239
rect 41391 189 41445 205
rect 41528 229 41558 413
rect 41636 257 41666 413
rect 41720 365 41750 413
rect 41708 349 41762 365
rect 41708 315 41718 349
rect 41752 315 41762 349
rect 41708 299 41762 315
rect 41631 241 41685 257
rect 41528 213 41589 229
rect 41528 193 41545 213
rect 41282 119 41312 141
rect 41391 119 41421 189
rect 41487 179 41545 193
rect 41579 179 41589 213
rect 41631 207 41641 241
rect 41675 207 41685 241
rect 41631 191 41685 207
rect 41487 163 41589 179
rect 41487 131 41517 163
rect 41636 131 41666 191
rect 41727 131 41757 299
rect 42103 333 42133 369
rect 42092 303 42133 333
rect 41884 265 41914 297
rect 42092 265 42122 303
rect 42200 265 42230 297
rect 41813 249 42122 265
rect 41813 215 41841 249
rect 41875 215 42122 249
rect 41813 199 42122 215
rect 42171 249 42230 265
rect 42171 215 42181 249
rect 42215 215 42230 249
rect 42171 199 42230 215
rect 41915 177 41945 199
rect 42092 176 42122 199
rect 42200 177 42230 199
rect 42092 146 42133 176
rect 42103 131 42133 146
rect 79 21 109 47
rect 163 21 193 47
rect 418 21 448 47
rect 513 21 543 47
rect 609 21 639 47
rect 775 21 805 47
rect 847 21 877 47
rect 979 21 1009 47
rect 1078 21 1108 47
rect 1187 21 1217 47
rect 1283 21 1313 47
rect 1432 21 1462 47
rect 1523 21 1553 47
rect 1711 21 1741 47
rect 1899 21 1929 47
rect 1996 21 2026 47
rect 2195 21 2225 47
rect 2279 21 2309 47
rect 2534 21 2564 47
rect 2629 21 2659 47
rect 2725 21 2755 47
rect 2891 21 2921 47
rect 2963 21 2993 47
rect 3095 21 3125 47
rect 3194 21 3224 47
rect 3303 21 3333 47
rect 3399 21 3429 47
rect 3548 21 3578 47
rect 3639 21 3669 47
rect 3827 21 3857 47
rect 4015 21 4045 47
rect 4112 21 4142 47
rect 4311 21 4341 47
rect 4395 21 4425 47
rect 4650 21 4680 47
rect 4745 21 4775 47
rect 4841 21 4871 47
rect 5007 21 5037 47
rect 5079 21 5109 47
rect 5211 21 5241 47
rect 5310 21 5340 47
rect 5419 21 5449 47
rect 5515 21 5545 47
rect 5664 21 5694 47
rect 5755 21 5785 47
rect 5943 21 5973 47
rect 6131 21 6161 47
rect 6228 21 6258 47
rect 6427 21 6457 47
rect 6511 21 6541 47
rect 6766 21 6796 47
rect 6861 21 6891 47
rect 6957 21 6987 47
rect 7123 21 7153 47
rect 7195 21 7225 47
rect 7327 21 7357 47
rect 7426 21 7456 47
rect 7535 21 7565 47
rect 7631 21 7661 47
rect 7780 21 7810 47
rect 7871 21 7901 47
rect 8059 21 8089 47
rect 8247 21 8277 47
rect 8344 21 8374 47
rect 8543 21 8573 47
rect 8627 21 8657 47
rect 8882 21 8912 47
rect 8977 21 9007 47
rect 9073 21 9103 47
rect 9239 21 9269 47
rect 9311 21 9341 47
rect 9443 21 9473 47
rect 9542 21 9572 47
rect 9651 21 9681 47
rect 9747 21 9777 47
rect 9896 21 9926 47
rect 9987 21 10017 47
rect 10175 21 10205 47
rect 10363 21 10393 47
rect 10460 21 10490 47
rect 10659 21 10689 47
rect 10743 21 10773 47
rect 10998 21 11028 47
rect 11093 21 11123 47
rect 11189 21 11219 47
rect 11355 21 11385 47
rect 11427 21 11457 47
rect 11559 21 11589 47
rect 11658 21 11688 47
rect 11767 21 11797 47
rect 11863 21 11893 47
rect 12012 21 12042 47
rect 12103 21 12133 47
rect 12291 21 12321 47
rect 12479 21 12509 47
rect 12576 21 12606 47
rect 12775 21 12805 47
rect 12859 21 12889 47
rect 13114 21 13144 47
rect 13209 21 13239 47
rect 13305 21 13335 47
rect 13471 21 13501 47
rect 13543 21 13573 47
rect 13675 21 13705 47
rect 13774 21 13804 47
rect 13883 21 13913 47
rect 13979 21 14009 47
rect 14128 21 14158 47
rect 14219 21 14249 47
rect 14407 21 14437 47
rect 14595 21 14625 47
rect 14692 21 14722 47
rect 14891 21 14921 47
rect 14975 21 15005 47
rect 15230 21 15260 47
rect 15325 21 15355 47
rect 15421 21 15451 47
rect 15587 21 15617 47
rect 15659 21 15689 47
rect 15791 21 15821 47
rect 15890 21 15920 47
rect 15999 21 16029 47
rect 16095 21 16125 47
rect 16244 21 16274 47
rect 16335 21 16365 47
rect 16523 21 16553 47
rect 16711 21 16741 47
rect 16808 21 16838 47
rect 17007 21 17037 47
rect 17091 21 17121 47
rect 17346 21 17376 47
rect 17441 21 17471 47
rect 17537 21 17567 47
rect 17703 21 17733 47
rect 17775 21 17805 47
rect 17907 21 17937 47
rect 18006 21 18036 47
rect 18115 21 18145 47
rect 18211 21 18241 47
rect 18360 21 18390 47
rect 18451 21 18481 47
rect 18639 21 18669 47
rect 18827 21 18857 47
rect 18924 21 18954 47
rect 19123 21 19153 47
rect 19207 21 19237 47
rect 19462 21 19492 47
rect 19557 21 19587 47
rect 19653 21 19683 47
rect 19819 21 19849 47
rect 19891 21 19921 47
rect 20023 21 20053 47
rect 20122 21 20152 47
rect 20231 21 20261 47
rect 20327 21 20357 47
rect 20476 21 20506 47
rect 20567 21 20597 47
rect 20755 21 20785 47
rect 20943 21 20973 47
rect 21040 21 21070 47
rect 21239 21 21269 47
rect 21323 21 21353 47
rect 21578 21 21608 47
rect 21673 21 21703 47
rect 21769 21 21799 47
rect 21935 21 21965 47
rect 22007 21 22037 47
rect 22139 21 22169 47
rect 22238 21 22268 47
rect 22347 21 22377 47
rect 22443 21 22473 47
rect 22592 21 22622 47
rect 22683 21 22713 47
rect 22871 21 22901 47
rect 23059 21 23089 47
rect 23156 21 23186 47
rect 23355 21 23385 47
rect 23439 21 23469 47
rect 23694 21 23724 47
rect 23789 21 23819 47
rect 23885 21 23915 47
rect 24051 21 24081 47
rect 24123 21 24153 47
rect 24255 21 24285 47
rect 24354 21 24384 47
rect 24463 21 24493 47
rect 24559 21 24589 47
rect 24708 21 24738 47
rect 24799 21 24829 47
rect 24987 21 25017 47
rect 25175 21 25205 47
rect 25272 21 25302 47
rect 25471 21 25501 47
rect 25555 21 25585 47
rect 25810 21 25840 47
rect 25905 21 25935 47
rect 26001 21 26031 47
rect 26167 21 26197 47
rect 26239 21 26269 47
rect 26371 21 26401 47
rect 26470 21 26500 47
rect 26579 21 26609 47
rect 26675 21 26705 47
rect 26824 21 26854 47
rect 26915 21 26945 47
rect 27103 21 27133 47
rect 27291 21 27321 47
rect 27388 21 27418 47
rect 27587 21 27617 47
rect 27671 21 27701 47
rect 27926 21 27956 47
rect 28021 21 28051 47
rect 28117 21 28147 47
rect 28283 21 28313 47
rect 28355 21 28385 47
rect 28487 21 28517 47
rect 28586 21 28616 47
rect 28695 21 28725 47
rect 28791 21 28821 47
rect 28940 21 28970 47
rect 29031 21 29061 47
rect 29219 21 29249 47
rect 29407 21 29437 47
rect 29504 21 29534 47
rect 29703 21 29733 47
rect 29787 21 29817 47
rect 30042 21 30072 47
rect 30137 21 30167 47
rect 30233 21 30263 47
rect 30399 21 30429 47
rect 30471 21 30501 47
rect 30603 21 30633 47
rect 30702 21 30732 47
rect 30811 21 30841 47
rect 30907 21 30937 47
rect 31056 21 31086 47
rect 31147 21 31177 47
rect 31335 21 31365 47
rect 31523 21 31553 47
rect 31620 21 31650 47
rect 31819 21 31849 47
rect 31903 21 31933 47
rect 32158 21 32188 47
rect 32253 21 32283 47
rect 32349 21 32379 47
rect 32515 21 32545 47
rect 32587 21 32617 47
rect 32719 21 32749 47
rect 32818 21 32848 47
rect 32927 21 32957 47
rect 33023 21 33053 47
rect 33172 21 33202 47
rect 33263 21 33293 47
rect 33451 21 33481 47
rect 33639 21 33669 47
rect 33736 21 33766 47
rect 33935 21 33965 47
rect 34019 21 34049 47
rect 34274 21 34304 47
rect 34369 21 34399 47
rect 34465 21 34495 47
rect 34631 21 34661 47
rect 34703 21 34733 47
rect 34835 21 34865 47
rect 34934 21 34964 47
rect 35043 21 35073 47
rect 35139 21 35169 47
rect 35288 21 35318 47
rect 35379 21 35409 47
rect 35567 21 35597 47
rect 35755 21 35785 47
rect 35852 21 35882 47
rect 36051 21 36081 47
rect 36135 21 36165 47
rect 36390 21 36420 47
rect 36485 21 36515 47
rect 36581 21 36611 47
rect 36747 21 36777 47
rect 36819 21 36849 47
rect 36951 21 36981 47
rect 37050 21 37080 47
rect 37159 21 37189 47
rect 37255 21 37285 47
rect 37404 21 37434 47
rect 37495 21 37525 47
rect 37683 21 37713 47
rect 37871 21 37901 47
rect 37968 21 37998 47
rect 38167 21 38197 47
rect 38251 21 38281 47
rect 38506 21 38536 47
rect 38601 21 38631 47
rect 38697 21 38727 47
rect 38863 21 38893 47
rect 38935 21 38965 47
rect 39067 21 39097 47
rect 39166 21 39196 47
rect 39275 21 39305 47
rect 39371 21 39401 47
rect 39520 21 39550 47
rect 39611 21 39641 47
rect 39799 21 39829 47
rect 39987 21 40017 47
rect 40084 21 40114 47
rect 40283 21 40313 47
rect 40367 21 40397 47
rect 40622 21 40652 47
rect 40717 21 40747 47
rect 40813 21 40843 47
rect 40979 21 41009 47
rect 41051 21 41081 47
rect 41183 21 41213 47
rect 41282 21 41312 47
rect 41391 21 41421 47
rect 41487 21 41517 47
rect 41636 21 41666 47
rect 41727 21 41757 47
rect 41915 21 41945 47
rect 42103 21 42133 47
rect 42200 21 42230 47
<< polycont >>
rect 32 215 66 249
rect 134 230 168 264
rect 522 331 556 365
rect 341 276 375 310
rect 771 305 805 339
rect 500 169 534 203
rect 602 163 636 197
rect 857 169 891 203
rect 953 217 987 251
rect 1236 331 1270 365
rect 1101 157 1135 191
rect 1197 205 1231 239
rect 1514 315 1548 349
rect 1341 179 1375 213
rect 1437 207 1471 241
rect 1637 215 1671 249
rect 1977 215 2011 249
rect 2148 215 2182 249
rect 2250 230 2284 264
rect 2638 331 2672 365
rect 2457 276 2491 310
rect 2887 305 2921 339
rect 2616 169 2650 203
rect 2718 163 2752 197
rect 2973 169 3007 203
rect 3069 217 3103 251
rect 3352 331 3386 365
rect 3217 157 3251 191
rect 3313 205 3347 239
rect 3630 315 3664 349
rect 3457 179 3491 213
rect 3553 207 3587 241
rect 3753 215 3787 249
rect 4093 215 4127 249
rect 4264 215 4298 249
rect 4366 230 4400 264
rect 4754 331 4788 365
rect 4573 276 4607 310
rect 5003 305 5037 339
rect 4732 169 4766 203
rect 4834 163 4868 197
rect 5089 169 5123 203
rect 5185 217 5219 251
rect 5468 331 5502 365
rect 5333 157 5367 191
rect 5429 205 5463 239
rect 5746 315 5780 349
rect 5573 179 5607 213
rect 5669 207 5703 241
rect 5869 215 5903 249
rect 6209 215 6243 249
rect 6380 215 6414 249
rect 6482 230 6516 264
rect 6870 331 6904 365
rect 6689 276 6723 310
rect 7119 305 7153 339
rect 6848 169 6882 203
rect 6950 163 6984 197
rect 7205 169 7239 203
rect 7301 217 7335 251
rect 7584 331 7618 365
rect 7449 157 7483 191
rect 7545 205 7579 239
rect 7862 315 7896 349
rect 7689 179 7723 213
rect 7785 207 7819 241
rect 7985 215 8019 249
rect 8325 215 8359 249
rect 8496 215 8530 249
rect 8598 230 8632 264
rect 8986 331 9020 365
rect 8805 276 8839 310
rect 9235 305 9269 339
rect 8964 169 8998 203
rect 9066 163 9100 197
rect 9321 169 9355 203
rect 9417 217 9451 251
rect 9700 331 9734 365
rect 9565 157 9599 191
rect 9661 205 9695 239
rect 9978 315 10012 349
rect 9805 179 9839 213
rect 9901 207 9935 241
rect 10101 215 10135 249
rect 10441 215 10475 249
rect 10612 215 10646 249
rect 10714 230 10748 264
rect 11102 331 11136 365
rect 10921 276 10955 310
rect 11351 305 11385 339
rect 11080 169 11114 203
rect 11182 163 11216 197
rect 11437 169 11471 203
rect 11533 217 11567 251
rect 11816 331 11850 365
rect 11681 157 11715 191
rect 11777 205 11811 239
rect 12094 315 12128 349
rect 11921 179 11955 213
rect 12017 207 12051 241
rect 12217 215 12251 249
rect 12557 215 12591 249
rect 12728 215 12762 249
rect 12830 230 12864 264
rect 13218 331 13252 365
rect 13037 276 13071 310
rect 13467 305 13501 339
rect 13196 169 13230 203
rect 13298 163 13332 197
rect 13553 169 13587 203
rect 13649 217 13683 251
rect 13932 331 13966 365
rect 13797 157 13831 191
rect 13893 205 13927 239
rect 14210 315 14244 349
rect 14037 179 14071 213
rect 14133 207 14167 241
rect 14333 215 14367 249
rect 14673 215 14707 249
rect 14844 215 14878 249
rect 14946 230 14980 264
rect 15334 331 15368 365
rect 15153 276 15187 310
rect 15583 305 15617 339
rect 15312 169 15346 203
rect 15414 163 15448 197
rect 15669 169 15703 203
rect 15765 217 15799 251
rect 16048 331 16082 365
rect 15913 157 15947 191
rect 16009 205 16043 239
rect 16326 315 16360 349
rect 16153 179 16187 213
rect 16249 207 16283 241
rect 16449 215 16483 249
rect 16789 215 16823 249
rect 16960 215 16994 249
rect 17062 230 17096 264
rect 17450 331 17484 365
rect 17269 276 17303 310
rect 17699 305 17733 339
rect 17428 169 17462 203
rect 17530 163 17564 197
rect 17785 169 17819 203
rect 17881 217 17915 251
rect 18164 331 18198 365
rect 18029 157 18063 191
rect 18125 205 18159 239
rect 18442 315 18476 349
rect 18269 179 18303 213
rect 18365 207 18399 241
rect 18565 215 18599 249
rect 18905 215 18939 249
rect 19076 215 19110 249
rect 19178 230 19212 264
rect 19566 331 19600 365
rect 19385 276 19419 310
rect 19815 305 19849 339
rect 19544 169 19578 203
rect 19646 163 19680 197
rect 19901 169 19935 203
rect 19997 217 20031 251
rect 20280 331 20314 365
rect 20145 157 20179 191
rect 20241 205 20275 239
rect 20558 315 20592 349
rect 20385 179 20419 213
rect 20481 207 20515 241
rect 20681 215 20715 249
rect 21021 215 21055 249
rect 21192 215 21226 249
rect 21294 230 21328 264
rect 21682 331 21716 365
rect 21501 276 21535 310
rect 21931 305 21965 339
rect 21660 169 21694 203
rect 21762 163 21796 197
rect 22017 169 22051 203
rect 22113 217 22147 251
rect 22396 331 22430 365
rect 22261 157 22295 191
rect 22357 205 22391 239
rect 22674 315 22708 349
rect 22501 179 22535 213
rect 22597 207 22631 241
rect 22797 215 22831 249
rect 23137 215 23171 249
rect 23308 215 23342 249
rect 23410 230 23444 264
rect 23798 331 23832 365
rect 23617 276 23651 310
rect 24047 305 24081 339
rect 23776 169 23810 203
rect 23878 163 23912 197
rect 24133 169 24167 203
rect 24229 217 24263 251
rect 24512 331 24546 365
rect 24377 157 24411 191
rect 24473 205 24507 239
rect 24790 315 24824 349
rect 24617 179 24651 213
rect 24713 207 24747 241
rect 24913 215 24947 249
rect 25253 215 25287 249
rect 25424 215 25458 249
rect 25526 230 25560 264
rect 25914 331 25948 365
rect 25733 276 25767 310
rect 26163 305 26197 339
rect 25892 169 25926 203
rect 25994 163 26028 197
rect 26249 169 26283 203
rect 26345 217 26379 251
rect 26628 331 26662 365
rect 26493 157 26527 191
rect 26589 205 26623 239
rect 26906 315 26940 349
rect 26733 179 26767 213
rect 26829 207 26863 241
rect 27029 215 27063 249
rect 27369 215 27403 249
rect 27540 215 27574 249
rect 27642 230 27676 264
rect 28030 331 28064 365
rect 27849 276 27883 310
rect 28279 305 28313 339
rect 28008 169 28042 203
rect 28110 163 28144 197
rect 28365 169 28399 203
rect 28461 217 28495 251
rect 28744 331 28778 365
rect 28609 157 28643 191
rect 28705 205 28739 239
rect 29022 315 29056 349
rect 28849 179 28883 213
rect 28945 207 28979 241
rect 29145 215 29179 249
rect 29485 215 29519 249
rect 29656 215 29690 249
rect 29758 230 29792 264
rect 30146 331 30180 365
rect 29965 276 29999 310
rect 30395 305 30429 339
rect 30124 169 30158 203
rect 30226 163 30260 197
rect 30481 169 30515 203
rect 30577 217 30611 251
rect 30860 331 30894 365
rect 30725 157 30759 191
rect 30821 205 30855 239
rect 31138 315 31172 349
rect 30965 179 30999 213
rect 31061 207 31095 241
rect 31261 215 31295 249
rect 31601 215 31635 249
rect 31772 215 31806 249
rect 31874 230 31908 264
rect 32262 331 32296 365
rect 32081 276 32115 310
rect 32511 305 32545 339
rect 32240 169 32274 203
rect 32342 163 32376 197
rect 32597 169 32631 203
rect 32693 217 32727 251
rect 32976 331 33010 365
rect 32841 157 32875 191
rect 32937 205 32971 239
rect 33254 315 33288 349
rect 33081 179 33115 213
rect 33177 207 33211 241
rect 33377 215 33411 249
rect 33717 215 33751 249
rect 33888 215 33922 249
rect 33990 230 34024 264
rect 34378 331 34412 365
rect 34197 276 34231 310
rect 34627 305 34661 339
rect 34356 169 34390 203
rect 34458 163 34492 197
rect 34713 169 34747 203
rect 34809 217 34843 251
rect 35092 331 35126 365
rect 34957 157 34991 191
rect 35053 205 35087 239
rect 35370 315 35404 349
rect 35197 179 35231 213
rect 35293 207 35327 241
rect 35493 215 35527 249
rect 35833 215 35867 249
rect 36004 215 36038 249
rect 36106 230 36140 264
rect 36494 331 36528 365
rect 36313 276 36347 310
rect 36743 305 36777 339
rect 36472 169 36506 203
rect 36574 163 36608 197
rect 36829 169 36863 203
rect 36925 217 36959 251
rect 37208 331 37242 365
rect 37073 157 37107 191
rect 37169 205 37203 239
rect 37486 315 37520 349
rect 37313 179 37347 213
rect 37409 207 37443 241
rect 37609 215 37643 249
rect 37949 215 37983 249
rect 38120 215 38154 249
rect 38222 230 38256 264
rect 38610 331 38644 365
rect 38429 276 38463 310
rect 38859 305 38893 339
rect 38588 169 38622 203
rect 38690 163 38724 197
rect 38945 169 38979 203
rect 39041 217 39075 251
rect 39324 331 39358 365
rect 39189 157 39223 191
rect 39285 205 39319 239
rect 39602 315 39636 349
rect 39429 179 39463 213
rect 39525 207 39559 241
rect 39725 215 39759 249
rect 40065 215 40099 249
rect 40236 215 40270 249
rect 40338 230 40372 264
rect 40726 331 40760 365
rect 40545 276 40579 310
rect 40975 305 41009 339
rect 40704 169 40738 203
rect 40806 163 40840 197
rect 41061 169 41095 203
rect 41157 217 41191 251
rect 41440 331 41474 365
rect 41305 157 41339 191
rect 41401 205 41435 239
rect 41718 315 41752 349
rect 41545 179 41579 213
rect 41641 207 41675 241
rect 41841 215 41875 249
rect 42181 215 42215 249
<< locali >>
rect 0 585 42320 601
rect 0 527 29 585
rect 63 527 121 585
rect 155 527 213 585
rect 247 527 305 585
rect 339 527 397 585
rect 431 527 489 585
rect 523 527 581 585
rect 615 527 673 585
rect 707 527 765 585
rect 799 527 857 585
rect 891 527 949 585
rect 983 527 1041 585
rect 1075 527 1133 585
rect 1167 527 1225 585
rect 1259 527 1317 585
rect 1351 527 1409 585
rect 1443 527 1501 585
rect 1535 527 1593 585
rect 1627 527 1685 585
rect 1719 527 1777 585
rect 1811 527 1869 585
rect 1903 527 1961 585
rect 1995 527 2053 585
rect 2087 527 2145 585
rect 2179 527 2237 585
rect 2271 527 2329 585
rect 2363 527 2421 585
rect 2455 527 2513 585
rect 2547 527 2605 585
rect 2639 527 2697 585
rect 2731 527 2789 585
rect 2823 527 2881 585
rect 2915 527 2973 585
rect 3007 527 3065 585
rect 3099 527 3157 585
rect 3191 527 3249 585
rect 3283 527 3341 585
rect 3375 527 3433 585
rect 3467 527 3525 585
rect 3559 527 3617 585
rect 3651 527 3709 585
rect 3743 527 3801 585
rect 3835 527 3893 585
rect 3927 527 3985 585
rect 4019 527 4077 585
rect 4111 527 4169 585
rect 4203 527 4261 585
rect 4295 527 4353 585
rect 4387 527 4445 585
rect 4479 527 4537 585
rect 4571 527 4629 585
rect 4663 527 4721 585
rect 4755 527 4813 585
rect 4847 527 4905 585
rect 4939 527 4997 585
rect 5031 527 5089 585
rect 5123 527 5181 585
rect 5215 527 5273 585
rect 5307 527 5365 585
rect 5399 527 5457 585
rect 5491 527 5549 585
rect 5583 527 5641 585
rect 5675 527 5733 585
rect 5767 527 5825 585
rect 5859 527 5917 585
rect 5951 527 6009 585
rect 6043 527 6101 585
rect 6135 527 6193 585
rect 6227 527 6285 585
rect 6319 527 6377 585
rect 6411 527 6469 585
rect 6503 527 6561 585
rect 6595 527 6653 585
rect 6687 527 6745 585
rect 6779 527 6837 585
rect 6871 527 6929 585
rect 6963 527 7021 585
rect 7055 527 7113 585
rect 7147 527 7205 585
rect 7239 527 7297 585
rect 7331 527 7389 585
rect 7423 527 7481 585
rect 7515 527 7573 585
rect 7607 527 7665 585
rect 7699 527 7757 585
rect 7791 527 7849 585
rect 7883 527 7941 585
rect 7975 527 8033 585
rect 8067 527 8125 585
rect 8159 527 8217 585
rect 8251 527 8309 585
rect 8343 527 8401 585
rect 8435 527 8493 585
rect 8527 527 8585 585
rect 8619 527 8677 585
rect 8711 527 8769 585
rect 8803 527 8861 585
rect 8895 527 8953 585
rect 8987 527 9045 585
rect 9079 527 9137 585
rect 9171 527 9229 585
rect 9263 527 9321 585
rect 9355 527 9413 585
rect 9447 527 9505 585
rect 9539 527 9597 585
rect 9631 527 9689 585
rect 9723 527 9781 585
rect 9815 527 9873 585
rect 9907 527 9965 585
rect 9999 527 10057 585
rect 10091 527 10149 585
rect 10183 527 10241 585
rect 10275 527 10333 585
rect 10367 527 10425 585
rect 10459 527 10517 585
rect 10551 527 10609 585
rect 10643 527 10701 585
rect 10735 527 10793 585
rect 10827 527 10885 585
rect 10919 527 10977 585
rect 11011 527 11069 585
rect 11103 527 11161 585
rect 11195 527 11253 585
rect 11287 527 11345 585
rect 11379 527 11437 585
rect 11471 527 11529 585
rect 11563 527 11621 585
rect 11655 527 11713 585
rect 11747 527 11805 585
rect 11839 527 11897 585
rect 11931 527 11989 585
rect 12023 527 12081 585
rect 12115 527 12173 585
rect 12207 527 12265 585
rect 12299 527 12357 585
rect 12391 527 12449 585
rect 12483 527 12541 585
rect 12575 527 12633 585
rect 12667 527 12725 585
rect 12759 527 12817 585
rect 12851 527 12909 585
rect 12943 527 13001 585
rect 13035 527 13093 585
rect 13127 527 13185 585
rect 13219 527 13277 585
rect 13311 527 13369 585
rect 13403 527 13461 585
rect 13495 527 13553 585
rect 13587 527 13645 585
rect 13679 527 13737 585
rect 13771 527 13829 585
rect 13863 527 13921 585
rect 13955 527 14013 585
rect 14047 527 14105 585
rect 14139 527 14197 585
rect 14231 527 14289 585
rect 14323 527 14381 585
rect 14415 527 14473 585
rect 14507 527 14565 585
rect 14599 527 14657 585
rect 14691 527 14749 585
rect 14783 527 14841 585
rect 14875 527 14933 585
rect 14967 527 15025 585
rect 15059 527 15117 585
rect 15151 527 15209 585
rect 15243 527 15301 585
rect 15335 527 15393 585
rect 15427 527 15485 585
rect 15519 527 15577 585
rect 15611 527 15669 585
rect 15703 527 15761 585
rect 15795 527 15853 585
rect 15887 527 15945 585
rect 15979 527 16037 585
rect 16071 527 16129 585
rect 16163 527 16221 585
rect 16255 527 16313 585
rect 16347 527 16405 585
rect 16439 527 16497 585
rect 16531 527 16589 585
rect 16623 527 16681 585
rect 16715 527 16773 585
rect 16807 527 16865 585
rect 16899 527 16957 585
rect 16991 527 17049 585
rect 17083 527 17141 585
rect 17175 527 17233 585
rect 17267 527 17325 585
rect 17359 527 17417 585
rect 17451 527 17509 585
rect 17543 527 17601 585
rect 17635 527 17693 585
rect 17727 527 17785 585
rect 17819 527 17877 585
rect 17911 527 17969 585
rect 18003 527 18061 585
rect 18095 527 18153 585
rect 18187 527 18245 585
rect 18279 527 18337 585
rect 18371 527 18429 585
rect 18463 527 18521 585
rect 18555 527 18613 585
rect 18647 527 18705 585
rect 18739 527 18797 585
rect 18831 527 18889 585
rect 18923 527 18981 585
rect 19015 527 19073 585
rect 19107 527 19165 585
rect 19199 527 19257 585
rect 19291 527 19349 585
rect 19383 527 19441 585
rect 19475 527 19533 585
rect 19567 527 19625 585
rect 19659 527 19717 585
rect 19751 527 19809 585
rect 19843 527 19901 585
rect 19935 527 19993 585
rect 20027 527 20085 585
rect 20119 527 20177 585
rect 20211 527 20269 585
rect 20303 527 20361 585
rect 20395 527 20453 585
rect 20487 527 20545 585
rect 20579 527 20637 585
rect 20671 527 20729 585
rect 20763 527 20821 585
rect 20855 527 20913 585
rect 20947 527 21005 585
rect 21039 527 21097 585
rect 21131 527 21189 585
rect 21223 527 21281 585
rect 21315 527 21373 585
rect 21407 527 21465 585
rect 21499 527 21557 585
rect 21591 527 21649 585
rect 21683 527 21741 585
rect 21775 527 21833 585
rect 21867 527 21925 585
rect 21959 527 22017 585
rect 22051 527 22109 585
rect 22143 527 22201 585
rect 22235 527 22293 585
rect 22327 527 22385 585
rect 22419 527 22477 585
rect 22511 527 22569 585
rect 22603 527 22661 585
rect 22695 527 22753 585
rect 22787 527 22845 585
rect 22879 527 22937 585
rect 22971 527 23029 585
rect 23063 527 23121 585
rect 23155 527 23213 585
rect 23247 527 23305 585
rect 23339 527 23397 585
rect 23431 527 23489 585
rect 23523 527 23581 585
rect 23615 527 23673 585
rect 23707 527 23765 585
rect 23799 527 23857 585
rect 23891 527 23949 585
rect 23983 527 24041 585
rect 24075 527 24133 585
rect 24167 527 24225 585
rect 24259 527 24317 585
rect 24351 527 24409 585
rect 24443 527 24501 585
rect 24535 527 24593 585
rect 24627 527 24685 585
rect 24719 527 24777 585
rect 24811 527 24869 585
rect 24903 527 24961 585
rect 24995 527 25053 585
rect 25087 527 25145 585
rect 25179 527 25237 585
rect 25271 527 25329 585
rect 25363 527 25421 585
rect 25455 527 25513 585
rect 25547 527 25605 585
rect 25639 527 25697 585
rect 25731 527 25789 585
rect 25823 527 25881 585
rect 25915 527 25973 585
rect 26007 527 26065 585
rect 26099 527 26157 585
rect 26191 527 26249 585
rect 26283 527 26341 585
rect 26375 527 26433 585
rect 26467 527 26525 585
rect 26559 527 26617 585
rect 26651 527 26709 585
rect 26743 527 26801 585
rect 26835 527 26893 585
rect 26927 527 26985 585
rect 27019 527 27077 585
rect 27111 527 27169 585
rect 27203 527 27261 585
rect 27295 527 27353 585
rect 27387 527 27445 585
rect 27479 527 27537 585
rect 27571 527 27629 585
rect 27663 527 27721 585
rect 27755 527 27813 585
rect 27847 527 27905 585
rect 27939 527 27997 585
rect 28031 527 28089 585
rect 28123 527 28181 585
rect 28215 527 28273 585
rect 28307 527 28365 585
rect 28399 527 28457 585
rect 28491 527 28549 585
rect 28583 527 28641 585
rect 28675 527 28733 585
rect 28767 527 28825 585
rect 28859 527 28917 585
rect 28951 527 29009 585
rect 29043 527 29101 585
rect 29135 527 29193 585
rect 29227 527 29285 585
rect 29319 527 29377 585
rect 29411 527 29469 585
rect 29503 527 29561 585
rect 29595 527 29653 585
rect 29687 527 29745 585
rect 29779 527 29837 585
rect 29871 527 29929 585
rect 29963 527 30021 585
rect 30055 527 30113 585
rect 30147 527 30205 585
rect 30239 527 30297 585
rect 30331 527 30389 585
rect 30423 527 30481 585
rect 30515 527 30573 585
rect 30607 527 30665 585
rect 30699 527 30757 585
rect 30791 527 30849 585
rect 30883 527 30941 585
rect 30975 527 31033 585
rect 31067 527 31125 585
rect 31159 527 31217 585
rect 31251 527 31309 585
rect 31343 527 31401 585
rect 31435 527 31493 585
rect 31527 527 31585 585
rect 31619 527 31677 585
rect 31711 527 31769 585
rect 31803 527 31861 585
rect 31895 527 31953 585
rect 31987 527 32045 585
rect 32079 527 32137 585
rect 32171 527 32229 585
rect 32263 527 32321 585
rect 32355 527 32413 585
rect 32447 527 32505 585
rect 32539 527 32597 585
rect 32631 527 32689 585
rect 32723 527 32781 585
rect 32815 527 32873 585
rect 32907 527 32965 585
rect 32999 527 33057 585
rect 33091 527 33149 585
rect 33183 527 33241 585
rect 33275 527 33333 585
rect 33367 527 33425 585
rect 33459 527 33517 585
rect 33551 527 33609 585
rect 33643 527 33701 585
rect 33735 527 33793 585
rect 33827 527 33885 585
rect 33919 527 33977 585
rect 34011 527 34069 585
rect 34103 527 34161 585
rect 34195 527 34253 585
rect 34287 527 34345 585
rect 34379 527 34437 585
rect 34471 527 34529 585
rect 34563 527 34621 585
rect 34655 527 34713 585
rect 34747 527 34805 585
rect 34839 527 34897 585
rect 34931 527 34989 585
rect 35023 527 35081 585
rect 35115 527 35173 585
rect 35207 527 35265 585
rect 35299 527 35357 585
rect 35391 527 35449 585
rect 35483 527 35541 585
rect 35575 527 35633 585
rect 35667 527 35725 585
rect 35759 527 35817 585
rect 35851 527 35909 585
rect 35943 527 36001 585
rect 36035 527 36093 585
rect 36127 527 36185 585
rect 36219 527 36277 585
rect 36311 527 36369 585
rect 36403 527 36461 585
rect 36495 527 36553 585
rect 36587 527 36645 585
rect 36679 527 36737 585
rect 36771 527 36829 585
rect 36863 527 36921 585
rect 36955 527 37013 585
rect 37047 527 37105 585
rect 37139 527 37197 585
rect 37231 527 37289 585
rect 37323 527 37381 585
rect 37415 527 37473 585
rect 37507 527 37565 585
rect 37599 527 37657 585
rect 37691 527 37749 585
rect 37783 527 37841 585
rect 37875 527 37933 585
rect 37967 527 38025 585
rect 38059 527 38117 585
rect 38151 527 38209 585
rect 38243 527 38301 585
rect 38335 527 38393 585
rect 38427 527 38485 585
rect 38519 527 38577 585
rect 38611 527 38669 585
rect 38703 527 38761 585
rect 38795 527 38853 585
rect 38887 527 38945 585
rect 38979 527 39037 585
rect 39071 527 39129 585
rect 39163 527 39221 585
rect 39255 527 39313 585
rect 39347 527 39405 585
rect 39439 527 39497 585
rect 39531 527 39589 585
rect 39623 527 39681 585
rect 39715 527 39773 585
rect 39807 527 39865 585
rect 39899 527 39957 585
rect 39991 527 40049 585
rect 40083 527 40141 585
rect 40175 527 40233 585
rect 40267 527 40325 585
rect 40359 527 40417 585
rect 40451 527 40509 585
rect 40543 527 40601 585
rect 40635 527 40693 585
rect 40727 527 40785 585
rect 40819 527 40877 585
rect 40911 527 40969 585
rect 41003 527 41061 585
rect 41095 527 41153 585
rect 41187 527 41245 585
rect 41279 527 41337 585
rect 41371 527 41429 585
rect 41463 527 41521 585
rect 41555 527 41613 585
rect 41647 527 41705 585
rect 41739 527 41797 585
rect 41831 527 41889 585
rect 41923 527 41981 585
rect 42015 527 42073 585
rect 42107 527 42165 585
rect 42199 527 42257 585
rect 42291 527 42320 585
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 18 375 35 409
rect 203 409 237 443
rect 69 375 168 393
rect 18 359 168 375
rect 0 249 88 325
rect 0 215 32 249
rect 66 215 88 249
rect 0 195 88 215
rect 122 264 168 359
rect 122 255 134 264
rect 156 221 168 230
rect 122 161 168 221
rect 18 127 168 161
rect 18 119 69 127
rect 18 85 35 119
rect 203 119 237 357
rect 271 333 336 490
rect 370 485 420 527
rect 370 451 386 485
rect 370 435 420 451
rect 454 477 504 493
rect 454 443 470 477
rect 454 427 504 443
rect 547 483 683 493
rect 547 449 563 483
rect 597 449 683 483
rect 798 475 864 527
rect 991 485 1065 527
rect 547 427 683 449
rect 454 401 488 427
rect 409 367 488 401
rect 522 391 615 393
rect 283 310 375 333
rect 283 276 341 310
rect 283 175 375 276
rect 283 141 307 175
rect 345 141 375 175
rect 283 123 375 141
rect 18 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 409 95 443 367
rect 522 365 581 391
rect 556 357 581 365
rect 556 331 615 357
rect 522 315 615 331
rect 477 255 547 277
rect 477 221 489 255
rect 523 221 547 255
rect 477 203 547 221
rect 477 169 500 203
rect 534 169 547 203
rect 477 153 547 169
rect 581 197 615 315
rect 649 271 683 427
rect 717 459 751 475
rect 798 441 814 475
rect 848 441 864 475
rect 898 459 932 475
rect 717 407 751 425
rect 991 451 1011 485
rect 1045 451 1065 485
rect 991 435 1065 451
rect 1099 477 1133 493
rect 898 407 932 425
rect 717 373 932 407
rect 1099 401 1133 443
rect 1180 484 1354 493
rect 1180 450 1196 484
rect 1230 450 1354 484
rect 1180 425 1354 450
rect 1388 485 1438 527
rect 1422 451 1438 485
rect 1542 485 1686 527
rect 1388 435 1438 451
rect 1472 459 1506 475
rect 1021 367 1133 401
rect 1021 339 1055 367
rect 755 305 771 339
rect 805 305 1055 339
rect 1194 357 1205 391
rect 1239 365 1286 391
rect 1194 333 1236 357
rect 649 251 987 271
rect 649 237 953 251
rect 581 163 602 197
rect 636 163 652 197
rect 581 153 652 163
rect 686 95 720 237
rect 761 187 857 203
rect 795 153 833 187
rect 891 169 919 203
rect 953 201 987 217
rect 867 153 919 169
rect 1021 167 1055 305
rect 203 69 237 85
rect 103 17 169 59
rect 309 55 325 89
rect 359 55 375 89
rect 409 61 458 95
rect 492 61 508 95
rect 549 61 565 95
rect 599 61 720 95
rect 895 93 961 109
rect 309 17 375 55
rect 895 59 911 93
rect 945 59 961 93
rect 895 17 961 59
rect 1003 89 1055 167
rect 1093 331 1236 333
rect 1270 331 1286 365
rect 1320 349 1354 425
rect 1542 451 1558 485
rect 1592 451 1636 485
rect 1670 451 1686 485
rect 1720 477 1801 493
rect 1952 485 1986 527
rect 1472 417 1506 425
rect 1754 443 1801 477
rect 1472 383 1632 417
rect 1093 299 1228 331
rect 1320 315 1514 349
rect 1548 315 1564 349
rect 1093 191 1135 299
rect 1320 297 1354 315
rect 1093 157 1101 191
rect 1093 141 1135 157
rect 1169 255 1239 265
rect 1169 239 1205 255
rect 1169 205 1197 239
rect 1231 205 1239 221
rect 1169 141 1239 205
rect 1273 263 1354 297
rect 1273 107 1307 263
rect 1421 250 1529 281
rect 1598 265 1632 383
rect 1720 409 1801 443
rect 1754 375 1801 409
rect 1720 341 1801 375
rect 1754 307 1801 341
rect 1720 291 1801 307
rect 1598 259 1687 265
rect 1455 241 1529 250
rect 1341 213 1385 229
rect 1375 179 1385 213
rect 1421 207 1437 216
rect 1471 207 1529 241
rect 1341 173 1385 179
rect 1481 187 1529 207
rect 1341 139 1447 173
rect 1117 93 1307 107
rect 1003 55 1023 89
rect 1057 55 1073 89
rect 1117 59 1133 93
rect 1167 59 1307 93
rect 1117 51 1307 59
rect 1341 89 1379 105
rect 1341 55 1345 89
rect 1413 93 1447 139
rect 1515 153 1529 187
rect 1481 127 1529 153
rect 1563 249 1687 259
rect 1563 215 1637 249
rect 1671 215 1687 249
rect 1563 199 1687 215
rect 1563 164 1628 199
rect 1735 165 1801 291
rect 1563 109 1627 164
rect 1413 75 1563 93
rect 1597 75 1627 109
rect 1413 59 1627 75
rect 1667 132 1701 154
rect 1341 17 1379 55
rect 1667 17 1701 98
rect 1735 131 1751 165
rect 1785 131 1801 165
rect 1735 97 1801 131
rect 1735 63 1751 97
rect 1785 63 1801 97
rect 1839 451 1855 485
rect 1889 451 1905 485
rect 1839 417 1905 451
rect 1839 383 1855 417
rect 1889 383 1905 417
rect 1839 265 1905 383
rect 2134 477 2185 493
rect 1952 417 1986 451
rect 1952 349 1986 383
rect 1952 299 1986 315
rect 2036 449 2087 465
rect 2070 415 2087 449
rect 2036 381 2087 415
rect 2070 347 2087 381
rect 2134 443 2151 477
rect 2134 409 2185 443
rect 2219 461 2285 527
rect 2219 427 2235 461
rect 2269 427 2285 461
rect 2319 477 2353 493
rect 2134 375 2151 409
rect 2319 409 2353 443
rect 2185 375 2284 393
rect 2134 359 2284 375
rect 2036 325 2087 347
rect 2036 289 2204 325
rect 2045 274 2204 289
rect 1839 249 2011 265
rect 1839 215 1977 249
rect 1839 199 2011 215
rect 2045 240 2076 274
rect 2114 249 2204 274
rect 2114 240 2148 249
rect 2045 215 2148 240
rect 2182 215 2204 249
rect 1839 119 1889 199
rect 2045 195 2204 215
rect 2238 264 2284 359
rect 2238 255 2250 264
rect 2272 221 2284 230
rect 2045 159 2087 195
rect 2238 161 2284 221
rect 2036 143 2087 159
rect 1839 85 1855 119
rect 1839 69 1889 85
rect 1952 113 1986 136
rect 1735 55 1801 63
rect 1952 17 1986 79
rect 2070 109 2087 143
rect 2036 53 2087 109
rect 2134 127 2284 161
rect 2134 119 2185 127
rect 2134 85 2151 119
rect 2319 119 2353 357
rect 2387 333 2452 490
rect 2486 485 2536 527
rect 2486 451 2502 485
rect 2486 435 2536 451
rect 2570 477 2620 493
rect 2570 443 2586 477
rect 2570 427 2620 443
rect 2663 483 2799 493
rect 2663 449 2679 483
rect 2713 449 2799 483
rect 2914 475 2980 527
rect 3107 485 3181 527
rect 2663 427 2799 449
rect 2570 401 2604 427
rect 2525 367 2604 401
rect 2638 391 2731 393
rect 2399 310 2491 333
rect 2399 276 2457 310
rect 2399 175 2491 276
rect 2399 141 2423 175
rect 2461 141 2491 175
rect 2399 123 2491 141
rect 2134 69 2185 85
rect 2219 59 2235 93
rect 2269 59 2285 93
rect 2525 95 2559 367
rect 2638 365 2697 391
rect 2672 357 2697 365
rect 2672 331 2731 357
rect 2638 315 2731 331
rect 2593 255 2663 277
rect 2593 221 2605 255
rect 2639 221 2663 255
rect 2593 203 2663 221
rect 2593 169 2616 203
rect 2650 169 2663 203
rect 2593 153 2663 169
rect 2697 197 2731 315
rect 2765 271 2799 427
rect 2833 459 2867 475
rect 2914 441 2930 475
rect 2964 441 2980 475
rect 3014 459 3048 475
rect 2833 407 2867 425
rect 3107 451 3127 485
rect 3161 451 3181 485
rect 3107 435 3181 451
rect 3215 477 3249 493
rect 3014 407 3048 425
rect 2833 373 3048 407
rect 3215 401 3249 443
rect 3296 484 3470 493
rect 3296 450 3312 484
rect 3346 450 3470 484
rect 3296 425 3470 450
rect 3504 485 3554 527
rect 3538 451 3554 485
rect 3658 485 3802 527
rect 3504 435 3554 451
rect 3588 459 3622 475
rect 3137 367 3249 401
rect 3137 339 3171 367
rect 2871 305 2887 339
rect 2921 305 3171 339
rect 3310 357 3321 391
rect 3355 365 3402 391
rect 3310 333 3352 357
rect 2765 251 3103 271
rect 2765 237 3069 251
rect 2697 163 2718 197
rect 2752 163 2768 197
rect 2697 153 2768 163
rect 2802 95 2836 237
rect 2877 187 2973 203
rect 2911 153 2949 187
rect 3007 169 3035 203
rect 3069 201 3103 217
rect 2983 153 3035 169
rect 3137 167 3171 305
rect 2319 69 2353 85
rect 2219 17 2285 59
rect 2425 55 2441 89
rect 2475 55 2491 89
rect 2525 61 2574 95
rect 2608 61 2624 95
rect 2665 61 2681 95
rect 2715 61 2836 95
rect 3011 93 3077 109
rect 2425 17 2491 55
rect 3011 59 3027 93
rect 3061 59 3077 93
rect 3011 17 3077 59
rect 3119 89 3171 167
rect 3209 331 3352 333
rect 3386 331 3402 365
rect 3436 349 3470 425
rect 3658 451 3674 485
rect 3708 451 3752 485
rect 3786 451 3802 485
rect 3836 477 3917 493
rect 4068 485 4102 527
rect 3588 417 3622 425
rect 3870 443 3917 477
rect 3588 383 3748 417
rect 3209 299 3344 331
rect 3436 315 3630 349
rect 3664 315 3680 349
rect 3209 191 3251 299
rect 3436 297 3470 315
rect 3209 157 3217 191
rect 3209 141 3251 157
rect 3285 255 3355 265
rect 3285 239 3321 255
rect 3285 205 3313 239
rect 3347 205 3355 221
rect 3285 141 3355 205
rect 3389 263 3470 297
rect 3389 107 3423 263
rect 3537 250 3645 281
rect 3714 265 3748 383
rect 3836 409 3917 443
rect 3870 375 3917 409
rect 3836 341 3917 375
rect 3870 307 3917 341
rect 3836 291 3917 307
rect 3714 259 3803 265
rect 3571 241 3645 250
rect 3457 213 3501 229
rect 3491 179 3501 213
rect 3537 207 3553 216
rect 3587 207 3645 241
rect 3457 173 3501 179
rect 3597 187 3645 207
rect 3457 139 3563 173
rect 3233 93 3423 107
rect 3119 55 3139 89
rect 3173 55 3189 89
rect 3233 59 3249 93
rect 3283 59 3423 93
rect 3233 51 3423 59
rect 3457 89 3495 105
rect 3457 55 3461 89
rect 3529 93 3563 139
rect 3631 153 3645 187
rect 3597 127 3645 153
rect 3679 249 3803 259
rect 3679 215 3753 249
rect 3787 215 3803 249
rect 3679 199 3803 215
rect 3679 164 3744 199
rect 3851 165 3917 291
rect 3679 109 3743 164
rect 3529 75 3679 93
rect 3713 75 3743 109
rect 3529 59 3743 75
rect 3783 132 3817 154
rect 3457 17 3495 55
rect 3783 17 3817 98
rect 3851 131 3867 165
rect 3901 131 3917 165
rect 3851 97 3917 131
rect 3851 63 3867 97
rect 3901 63 3917 97
rect 3955 451 3971 485
rect 4005 451 4021 485
rect 3955 417 4021 451
rect 3955 383 3971 417
rect 4005 383 4021 417
rect 3955 265 4021 383
rect 4250 477 4301 493
rect 4068 417 4102 451
rect 4068 349 4102 383
rect 4068 299 4102 315
rect 4152 449 4203 465
rect 4186 415 4203 449
rect 4152 381 4203 415
rect 4186 347 4203 381
rect 4250 443 4267 477
rect 4250 409 4301 443
rect 4335 461 4401 527
rect 4335 427 4351 461
rect 4385 427 4401 461
rect 4435 477 4469 493
rect 4250 375 4267 409
rect 4435 409 4469 443
rect 4301 375 4400 393
rect 4250 359 4400 375
rect 4152 325 4203 347
rect 4152 289 4320 325
rect 4161 274 4320 289
rect 3955 249 4127 265
rect 3955 215 4093 249
rect 3955 199 4127 215
rect 4161 240 4192 274
rect 4230 249 4320 274
rect 4230 240 4264 249
rect 4161 215 4264 240
rect 4298 215 4320 249
rect 3955 119 4005 199
rect 4161 195 4320 215
rect 4354 264 4400 359
rect 4354 255 4366 264
rect 4388 221 4400 230
rect 4161 159 4203 195
rect 4354 161 4400 221
rect 4152 143 4203 159
rect 3955 85 3971 119
rect 3955 69 4005 85
rect 4068 113 4102 136
rect 3851 55 3917 63
rect 4068 17 4102 79
rect 4186 109 4203 143
rect 4152 53 4203 109
rect 4250 127 4400 161
rect 4250 119 4301 127
rect 4250 85 4267 119
rect 4435 119 4469 357
rect 4503 333 4568 490
rect 4602 485 4652 527
rect 4602 451 4618 485
rect 4602 435 4652 451
rect 4686 477 4736 493
rect 4686 443 4702 477
rect 4686 427 4736 443
rect 4779 483 4915 493
rect 4779 449 4795 483
rect 4829 449 4915 483
rect 5030 475 5096 527
rect 5223 485 5297 527
rect 4779 427 4915 449
rect 4686 401 4720 427
rect 4641 367 4720 401
rect 4754 391 4847 393
rect 4515 310 4607 333
rect 4515 276 4573 310
rect 4515 175 4607 276
rect 4515 141 4539 175
rect 4577 141 4607 175
rect 4515 123 4607 141
rect 4250 69 4301 85
rect 4335 59 4351 93
rect 4385 59 4401 93
rect 4641 95 4675 367
rect 4754 365 4813 391
rect 4788 357 4813 365
rect 4788 331 4847 357
rect 4754 315 4847 331
rect 4709 255 4779 277
rect 4709 221 4721 255
rect 4755 221 4779 255
rect 4709 203 4779 221
rect 4709 169 4732 203
rect 4766 169 4779 203
rect 4709 153 4779 169
rect 4813 197 4847 315
rect 4881 271 4915 427
rect 4949 459 4983 475
rect 5030 441 5046 475
rect 5080 441 5096 475
rect 5130 459 5164 475
rect 4949 407 4983 425
rect 5223 451 5243 485
rect 5277 451 5297 485
rect 5223 435 5297 451
rect 5331 477 5365 493
rect 5130 407 5164 425
rect 4949 373 5164 407
rect 5331 401 5365 443
rect 5412 484 5586 493
rect 5412 450 5428 484
rect 5462 450 5586 484
rect 5412 425 5586 450
rect 5620 485 5670 527
rect 5654 451 5670 485
rect 5774 485 5918 527
rect 5620 435 5670 451
rect 5704 459 5738 475
rect 5253 367 5365 401
rect 5253 339 5287 367
rect 4987 305 5003 339
rect 5037 305 5287 339
rect 5426 357 5437 391
rect 5471 365 5518 391
rect 5426 333 5468 357
rect 4881 251 5219 271
rect 4881 237 5185 251
rect 4813 163 4834 197
rect 4868 163 4884 197
rect 4813 153 4884 163
rect 4918 95 4952 237
rect 4993 187 5089 203
rect 5027 153 5065 187
rect 5123 169 5151 203
rect 5185 201 5219 217
rect 5099 153 5151 169
rect 5253 167 5287 305
rect 4435 69 4469 85
rect 4335 17 4401 59
rect 4541 55 4557 89
rect 4591 55 4607 89
rect 4641 61 4690 95
rect 4724 61 4740 95
rect 4781 61 4797 95
rect 4831 61 4952 95
rect 5127 93 5193 109
rect 4541 17 4607 55
rect 5127 59 5143 93
rect 5177 59 5193 93
rect 5127 17 5193 59
rect 5235 89 5287 167
rect 5325 331 5468 333
rect 5502 331 5518 365
rect 5552 349 5586 425
rect 5774 451 5790 485
rect 5824 451 5868 485
rect 5902 451 5918 485
rect 5952 477 6033 493
rect 6184 485 6218 527
rect 5704 417 5738 425
rect 5986 443 6033 477
rect 5704 383 5864 417
rect 5325 299 5460 331
rect 5552 315 5746 349
rect 5780 315 5796 349
rect 5325 191 5367 299
rect 5552 297 5586 315
rect 5325 157 5333 191
rect 5325 141 5367 157
rect 5401 255 5471 265
rect 5401 239 5437 255
rect 5401 205 5429 239
rect 5463 205 5471 221
rect 5401 141 5471 205
rect 5505 263 5586 297
rect 5505 107 5539 263
rect 5653 250 5761 281
rect 5830 265 5864 383
rect 5952 409 6033 443
rect 5986 375 6033 409
rect 5952 341 6033 375
rect 5986 307 6033 341
rect 5952 291 6033 307
rect 5830 259 5919 265
rect 5687 241 5761 250
rect 5573 213 5617 229
rect 5607 179 5617 213
rect 5653 207 5669 216
rect 5703 207 5761 241
rect 5573 173 5617 179
rect 5713 187 5761 207
rect 5573 139 5679 173
rect 5349 93 5539 107
rect 5235 55 5255 89
rect 5289 55 5305 89
rect 5349 59 5365 93
rect 5399 59 5539 93
rect 5349 51 5539 59
rect 5573 89 5611 105
rect 5573 55 5577 89
rect 5645 93 5679 139
rect 5747 153 5761 187
rect 5713 127 5761 153
rect 5795 249 5919 259
rect 5795 215 5869 249
rect 5903 215 5919 249
rect 5795 199 5919 215
rect 5795 164 5860 199
rect 5967 165 6033 291
rect 5795 109 5859 164
rect 5645 75 5795 93
rect 5829 75 5859 109
rect 5645 59 5859 75
rect 5899 132 5933 154
rect 5573 17 5611 55
rect 5899 17 5933 98
rect 5967 131 5983 165
rect 6017 131 6033 165
rect 5967 97 6033 131
rect 5967 63 5983 97
rect 6017 63 6033 97
rect 6071 451 6087 485
rect 6121 451 6137 485
rect 6071 417 6137 451
rect 6071 383 6087 417
rect 6121 383 6137 417
rect 6071 265 6137 383
rect 6366 477 6417 493
rect 6184 417 6218 451
rect 6184 349 6218 383
rect 6184 299 6218 315
rect 6268 449 6319 465
rect 6302 415 6319 449
rect 6268 381 6319 415
rect 6302 347 6319 381
rect 6366 443 6383 477
rect 6366 409 6417 443
rect 6451 461 6517 527
rect 6451 427 6467 461
rect 6501 427 6517 461
rect 6551 477 6585 493
rect 6366 375 6383 409
rect 6551 409 6585 443
rect 6417 375 6516 393
rect 6366 359 6516 375
rect 6268 325 6319 347
rect 6268 289 6436 325
rect 6277 274 6436 289
rect 6071 249 6243 265
rect 6071 215 6209 249
rect 6071 199 6243 215
rect 6277 240 6308 274
rect 6346 249 6436 274
rect 6346 240 6380 249
rect 6277 215 6380 240
rect 6414 215 6436 249
rect 6071 119 6121 199
rect 6277 195 6436 215
rect 6470 264 6516 359
rect 6470 255 6482 264
rect 6504 221 6516 230
rect 6277 159 6319 195
rect 6470 161 6516 221
rect 6268 143 6319 159
rect 6071 85 6087 119
rect 6071 69 6121 85
rect 6184 113 6218 136
rect 5967 55 6033 63
rect 6184 17 6218 79
rect 6302 109 6319 143
rect 6268 53 6319 109
rect 6366 127 6516 161
rect 6366 119 6417 127
rect 6366 85 6383 119
rect 6551 119 6585 357
rect 6619 333 6684 490
rect 6718 485 6768 527
rect 6718 451 6734 485
rect 6718 435 6768 451
rect 6802 477 6852 493
rect 6802 443 6818 477
rect 6802 427 6852 443
rect 6895 483 7031 493
rect 6895 449 6911 483
rect 6945 449 7031 483
rect 7146 475 7212 527
rect 7339 485 7413 527
rect 6895 427 7031 449
rect 6802 401 6836 427
rect 6757 367 6836 401
rect 6870 391 6963 393
rect 6631 310 6723 333
rect 6631 276 6689 310
rect 6631 175 6723 276
rect 6631 141 6655 175
rect 6693 141 6723 175
rect 6631 123 6723 141
rect 6366 69 6417 85
rect 6451 59 6467 93
rect 6501 59 6517 93
rect 6757 95 6791 367
rect 6870 365 6929 391
rect 6904 357 6929 365
rect 6904 331 6963 357
rect 6870 315 6963 331
rect 6825 255 6895 277
rect 6825 221 6837 255
rect 6871 221 6895 255
rect 6825 203 6895 221
rect 6825 169 6848 203
rect 6882 169 6895 203
rect 6825 153 6895 169
rect 6929 197 6963 315
rect 6997 271 7031 427
rect 7065 459 7099 475
rect 7146 441 7162 475
rect 7196 441 7212 475
rect 7246 459 7280 475
rect 7065 407 7099 425
rect 7339 451 7359 485
rect 7393 451 7413 485
rect 7339 435 7413 451
rect 7447 477 7481 493
rect 7246 407 7280 425
rect 7065 373 7280 407
rect 7447 401 7481 443
rect 7528 484 7702 493
rect 7528 450 7544 484
rect 7578 450 7702 484
rect 7528 425 7702 450
rect 7736 485 7786 527
rect 7770 451 7786 485
rect 7890 485 8034 527
rect 7736 435 7786 451
rect 7820 459 7854 475
rect 7369 367 7481 401
rect 7369 339 7403 367
rect 7103 305 7119 339
rect 7153 305 7403 339
rect 7542 357 7553 391
rect 7587 365 7634 391
rect 7542 333 7584 357
rect 6997 251 7335 271
rect 6997 237 7301 251
rect 6929 163 6950 197
rect 6984 163 7000 197
rect 6929 153 7000 163
rect 7034 95 7068 237
rect 7109 187 7205 203
rect 7143 153 7181 187
rect 7239 169 7267 203
rect 7301 201 7335 217
rect 7215 153 7267 169
rect 7369 167 7403 305
rect 6551 69 6585 85
rect 6451 17 6517 59
rect 6657 55 6673 89
rect 6707 55 6723 89
rect 6757 61 6806 95
rect 6840 61 6856 95
rect 6897 61 6913 95
rect 6947 61 7068 95
rect 7243 93 7309 109
rect 6657 17 6723 55
rect 7243 59 7259 93
rect 7293 59 7309 93
rect 7243 17 7309 59
rect 7351 89 7403 167
rect 7441 331 7584 333
rect 7618 331 7634 365
rect 7668 349 7702 425
rect 7890 451 7906 485
rect 7940 451 7984 485
rect 8018 451 8034 485
rect 8068 477 8149 493
rect 8300 485 8334 527
rect 7820 417 7854 425
rect 8102 443 8149 477
rect 7820 383 7980 417
rect 7441 299 7576 331
rect 7668 315 7862 349
rect 7896 315 7912 349
rect 7441 191 7483 299
rect 7668 297 7702 315
rect 7441 157 7449 191
rect 7441 141 7483 157
rect 7517 255 7587 265
rect 7517 239 7553 255
rect 7517 205 7545 239
rect 7579 205 7587 221
rect 7517 141 7587 205
rect 7621 263 7702 297
rect 7621 107 7655 263
rect 7769 250 7877 281
rect 7946 265 7980 383
rect 8068 409 8149 443
rect 8102 375 8149 409
rect 8068 341 8149 375
rect 8102 307 8149 341
rect 8068 291 8149 307
rect 7946 259 8035 265
rect 7803 241 7877 250
rect 7689 213 7733 229
rect 7723 179 7733 213
rect 7769 207 7785 216
rect 7819 207 7877 241
rect 7689 173 7733 179
rect 7829 187 7877 207
rect 7689 139 7795 173
rect 7465 93 7655 107
rect 7351 55 7371 89
rect 7405 55 7421 89
rect 7465 59 7481 93
rect 7515 59 7655 93
rect 7465 51 7655 59
rect 7689 89 7727 105
rect 7689 55 7693 89
rect 7761 93 7795 139
rect 7863 153 7877 187
rect 7829 127 7877 153
rect 7911 249 8035 259
rect 7911 215 7985 249
rect 8019 215 8035 249
rect 7911 199 8035 215
rect 7911 164 7976 199
rect 8083 165 8149 291
rect 7911 109 7975 164
rect 7761 75 7911 93
rect 7945 75 7975 109
rect 7761 59 7975 75
rect 8015 132 8049 154
rect 7689 17 7727 55
rect 8015 17 8049 98
rect 8083 131 8099 165
rect 8133 131 8149 165
rect 8083 97 8149 131
rect 8083 63 8099 97
rect 8133 63 8149 97
rect 8187 451 8203 485
rect 8237 451 8253 485
rect 8187 417 8253 451
rect 8187 383 8203 417
rect 8237 383 8253 417
rect 8187 265 8253 383
rect 8482 477 8533 493
rect 8300 417 8334 451
rect 8300 349 8334 383
rect 8300 299 8334 315
rect 8384 449 8435 465
rect 8418 415 8435 449
rect 8384 381 8435 415
rect 8418 347 8435 381
rect 8482 443 8499 477
rect 8482 409 8533 443
rect 8567 461 8633 527
rect 8567 427 8583 461
rect 8617 427 8633 461
rect 8667 477 8701 493
rect 8482 375 8499 409
rect 8667 409 8701 443
rect 8533 375 8632 393
rect 8482 359 8632 375
rect 8384 325 8435 347
rect 8384 289 8552 325
rect 8393 274 8552 289
rect 8187 249 8359 265
rect 8187 215 8325 249
rect 8187 199 8359 215
rect 8393 240 8424 274
rect 8462 249 8552 274
rect 8462 240 8496 249
rect 8393 215 8496 240
rect 8530 215 8552 249
rect 8187 119 8237 199
rect 8393 195 8552 215
rect 8586 264 8632 359
rect 8586 255 8598 264
rect 8620 221 8632 230
rect 8393 159 8435 195
rect 8586 161 8632 221
rect 8384 143 8435 159
rect 8187 85 8203 119
rect 8187 69 8237 85
rect 8300 113 8334 136
rect 8083 55 8149 63
rect 8300 17 8334 79
rect 8418 109 8435 143
rect 8384 53 8435 109
rect 8482 127 8632 161
rect 8482 119 8533 127
rect 8482 85 8499 119
rect 8667 119 8701 357
rect 8735 333 8800 490
rect 8834 485 8884 527
rect 8834 451 8850 485
rect 8834 435 8884 451
rect 8918 477 8968 493
rect 8918 443 8934 477
rect 8918 427 8968 443
rect 9011 483 9147 493
rect 9011 449 9027 483
rect 9061 449 9147 483
rect 9262 475 9328 527
rect 9455 485 9529 527
rect 9011 427 9147 449
rect 8918 401 8952 427
rect 8873 367 8952 401
rect 8986 391 9079 393
rect 8747 310 8839 333
rect 8747 276 8805 310
rect 8747 175 8839 276
rect 8747 141 8771 175
rect 8809 141 8839 175
rect 8747 123 8839 141
rect 8482 69 8533 85
rect 8567 59 8583 93
rect 8617 59 8633 93
rect 8873 95 8907 367
rect 8986 365 9045 391
rect 9020 357 9045 365
rect 9020 331 9079 357
rect 8986 315 9079 331
rect 8941 255 9011 277
rect 8941 221 8953 255
rect 8987 221 9011 255
rect 8941 203 9011 221
rect 8941 169 8964 203
rect 8998 169 9011 203
rect 8941 153 9011 169
rect 9045 197 9079 315
rect 9113 271 9147 427
rect 9181 459 9215 475
rect 9262 441 9278 475
rect 9312 441 9328 475
rect 9362 459 9396 475
rect 9181 407 9215 425
rect 9455 451 9475 485
rect 9509 451 9529 485
rect 9455 435 9529 451
rect 9563 477 9597 493
rect 9362 407 9396 425
rect 9181 373 9396 407
rect 9563 401 9597 443
rect 9644 484 9818 493
rect 9644 450 9660 484
rect 9694 450 9818 484
rect 9644 425 9818 450
rect 9852 485 9902 527
rect 9886 451 9902 485
rect 10006 485 10150 527
rect 9852 435 9902 451
rect 9936 459 9970 475
rect 9485 367 9597 401
rect 9485 339 9519 367
rect 9219 305 9235 339
rect 9269 305 9519 339
rect 9658 357 9669 391
rect 9703 365 9750 391
rect 9658 333 9700 357
rect 9113 251 9451 271
rect 9113 237 9417 251
rect 9045 163 9066 197
rect 9100 163 9116 197
rect 9045 153 9116 163
rect 9150 95 9184 237
rect 9225 187 9321 203
rect 9259 153 9297 187
rect 9355 169 9383 203
rect 9417 201 9451 217
rect 9331 153 9383 169
rect 9485 167 9519 305
rect 8667 69 8701 85
rect 8567 17 8633 59
rect 8773 55 8789 89
rect 8823 55 8839 89
rect 8873 61 8922 95
rect 8956 61 8972 95
rect 9013 61 9029 95
rect 9063 61 9184 95
rect 9359 93 9425 109
rect 8773 17 8839 55
rect 9359 59 9375 93
rect 9409 59 9425 93
rect 9359 17 9425 59
rect 9467 89 9519 167
rect 9557 331 9700 333
rect 9734 331 9750 365
rect 9784 349 9818 425
rect 10006 451 10022 485
rect 10056 451 10100 485
rect 10134 451 10150 485
rect 10184 477 10265 493
rect 10416 485 10450 527
rect 9936 417 9970 425
rect 10218 443 10265 477
rect 9936 383 10096 417
rect 9557 299 9692 331
rect 9784 315 9978 349
rect 10012 315 10028 349
rect 9557 191 9599 299
rect 9784 297 9818 315
rect 9557 157 9565 191
rect 9557 141 9599 157
rect 9633 255 9703 265
rect 9633 239 9669 255
rect 9633 205 9661 239
rect 9695 205 9703 221
rect 9633 141 9703 205
rect 9737 263 9818 297
rect 9737 107 9771 263
rect 9885 250 9993 281
rect 10062 265 10096 383
rect 10184 409 10265 443
rect 10218 375 10265 409
rect 10184 341 10265 375
rect 10218 307 10265 341
rect 10184 291 10265 307
rect 10062 259 10151 265
rect 9919 241 9993 250
rect 9805 213 9849 229
rect 9839 179 9849 213
rect 9885 207 9901 216
rect 9935 207 9993 241
rect 9805 173 9849 179
rect 9945 187 9993 207
rect 9805 139 9911 173
rect 9581 93 9771 107
rect 9467 55 9487 89
rect 9521 55 9537 89
rect 9581 59 9597 93
rect 9631 59 9771 93
rect 9581 51 9771 59
rect 9805 89 9843 105
rect 9805 55 9809 89
rect 9877 93 9911 139
rect 9979 153 9993 187
rect 9945 127 9993 153
rect 10027 249 10151 259
rect 10027 215 10101 249
rect 10135 215 10151 249
rect 10027 199 10151 215
rect 10027 164 10092 199
rect 10199 165 10265 291
rect 10027 109 10091 164
rect 9877 75 10027 93
rect 10061 75 10091 109
rect 9877 59 10091 75
rect 10131 132 10165 154
rect 9805 17 9843 55
rect 10131 17 10165 98
rect 10199 131 10215 165
rect 10249 131 10265 165
rect 10199 97 10265 131
rect 10199 63 10215 97
rect 10249 63 10265 97
rect 10303 451 10319 485
rect 10353 451 10369 485
rect 10303 417 10369 451
rect 10303 383 10319 417
rect 10353 383 10369 417
rect 10303 265 10369 383
rect 10598 477 10649 493
rect 10416 417 10450 451
rect 10416 349 10450 383
rect 10416 299 10450 315
rect 10500 449 10551 465
rect 10534 415 10551 449
rect 10500 381 10551 415
rect 10534 347 10551 381
rect 10598 443 10615 477
rect 10598 409 10649 443
rect 10683 461 10749 527
rect 10683 427 10699 461
rect 10733 427 10749 461
rect 10783 477 10817 493
rect 10598 375 10615 409
rect 10783 409 10817 443
rect 10649 375 10748 393
rect 10598 359 10748 375
rect 10500 325 10551 347
rect 10500 289 10668 325
rect 10509 274 10668 289
rect 10303 249 10475 265
rect 10303 215 10441 249
rect 10303 199 10475 215
rect 10509 240 10540 274
rect 10578 249 10668 274
rect 10578 240 10612 249
rect 10509 215 10612 240
rect 10646 215 10668 249
rect 10303 119 10353 199
rect 10509 195 10668 215
rect 10702 264 10748 359
rect 10702 255 10714 264
rect 10736 221 10748 230
rect 10509 159 10551 195
rect 10702 161 10748 221
rect 10500 143 10551 159
rect 10303 85 10319 119
rect 10303 69 10353 85
rect 10416 113 10450 136
rect 10199 55 10265 63
rect 10416 17 10450 79
rect 10534 109 10551 143
rect 10500 53 10551 109
rect 10598 127 10748 161
rect 10598 119 10649 127
rect 10598 85 10615 119
rect 10783 119 10817 357
rect 10851 333 10916 490
rect 10950 485 11000 527
rect 10950 451 10966 485
rect 10950 435 11000 451
rect 11034 477 11084 493
rect 11034 443 11050 477
rect 11034 427 11084 443
rect 11127 483 11263 493
rect 11127 449 11143 483
rect 11177 449 11263 483
rect 11378 475 11444 527
rect 11571 485 11645 527
rect 11127 427 11263 449
rect 11034 401 11068 427
rect 10989 367 11068 401
rect 11102 391 11195 393
rect 10863 310 10955 333
rect 10863 276 10921 310
rect 10863 175 10955 276
rect 10863 141 10887 175
rect 10925 141 10955 175
rect 10863 123 10955 141
rect 10598 69 10649 85
rect 10683 59 10699 93
rect 10733 59 10749 93
rect 10989 95 11023 367
rect 11102 365 11161 391
rect 11136 357 11161 365
rect 11136 331 11195 357
rect 11102 315 11195 331
rect 11057 255 11127 277
rect 11057 221 11069 255
rect 11103 221 11127 255
rect 11057 203 11127 221
rect 11057 169 11080 203
rect 11114 169 11127 203
rect 11057 153 11127 169
rect 11161 197 11195 315
rect 11229 271 11263 427
rect 11297 459 11331 475
rect 11378 441 11394 475
rect 11428 441 11444 475
rect 11478 459 11512 475
rect 11297 407 11331 425
rect 11571 451 11591 485
rect 11625 451 11645 485
rect 11571 435 11645 451
rect 11679 477 11713 493
rect 11478 407 11512 425
rect 11297 373 11512 407
rect 11679 401 11713 443
rect 11760 484 11934 493
rect 11760 450 11776 484
rect 11810 450 11934 484
rect 11760 425 11934 450
rect 11968 485 12018 527
rect 12002 451 12018 485
rect 12122 485 12266 527
rect 11968 435 12018 451
rect 12052 459 12086 475
rect 11601 367 11713 401
rect 11601 339 11635 367
rect 11335 305 11351 339
rect 11385 305 11635 339
rect 11774 357 11785 391
rect 11819 365 11866 391
rect 11774 333 11816 357
rect 11229 251 11567 271
rect 11229 237 11533 251
rect 11161 163 11182 197
rect 11216 163 11232 197
rect 11161 153 11232 163
rect 11266 95 11300 237
rect 11341 187 11437 203
rect 11375 153 11413 187
rect 11471 169 11499 203
rect 11533 201 11567 217
rect 11447 153 11499 169
rect 11601 167 11635 305
rect 10783 69 10817 85
rect 10683 17 10749 59
rect 10889 55 10905 89
rect 10939 55 10955 89
rect 10989 61 11038 95
rect 11072 61 11088 95
rect 11129 61 11145 95
rect 11179 61 11300 95
rect 11475 93 11541 109
rect 10889 17 10955 55
rect 11475 59 11491 93
rect 11525 59 11541 93
rect 11475 17 11541 59
rect 11583 89 11635 167
rect 11673 331 11816 333
rect 11850 331 11866 365
rect 11900 349 11934 425
rect 12122 451 12138 485
rect 12172 451 12216 485
rect 12250 451 12266 485
rect 12300 477 12381 493
rect 12532 485 12566 527
rect 12052 417 12086 425
rect 12334 443 12381 477
rect 12052 383 12212 417
rect 11673 299 11808 331
rect 11900 315 12094 349
rect 12128 315 12144 349
rect 11673 191 11715 299
rect 11900 297 11934 315
rect 11673 157 11681 191
rect 11673 141 11715 157
rect 11749 255 11819 265
rect 11749 239 11785 255
rect 11749 205 11777 239
rect 11811 205 11819 221
rect 11749 141 11819 205
rect 11853 263 11934 297
rect 11853 107 11887 263
rect 12001 250 12109 281
rect 12178 265 12212 383
rect 12300 409 12381 443
rect 12334 375 12381 409
rect 12300 341 12381 375
rect 12334 307 12381 341
rect 12300 291 12381 307
rect 12178 259 12267 265
rect 12035 241 12109 250
rect 11921 213 11965 229
rect 11955 179 11965 213
rect 12001 207 12017 216
rect 12051 207 12109 241
rect 11921 173 11965 179
rect 12061 187 12109 207
rect 11921 139 12027 173
rect 11697 93 11887 107
rect 11583 55 11603 89
rect 11637 55 11653 89
rect 11697 59 11713 93
rect 11747 59 11887 93
rect 11697 51 11887 59
rect 11921 89 11959 105
rect 11921 55 11925 89
rect 11993 93 12027 139
rect 12095 153 12109 187
rect 12061 127 12109 153
rect 12143 249 12267 259
rect 12143 215 12217 249
rect 12251 215 12267 249
rect 12143 199 12267 215
rect 12143 164 12208 199
rect 12315 165 12381 291
rect 12143 109 12207 164
rect 11993 75 12143 93
rect 12177 75 12207 109
rect 11993 59 12207 75
rect 12247 132 12281 154
rect 11921 17 11959 55
rect 12247 17 12281 98
rect 12315 131 12331 165
rect 12365 131 12381 165
rect 12315 97 12381 131
rect 12315 63 12331 97
rect 12365 63 12381 97
rect 12419 451 12435 485
rect 12469 451 12485 485
rect 12419 417 12485 451
rect 12419 383 12435 417
rect 12469 383 12485 417
rect 12419 265 12485 383
rect 12714 477 12765 493
rect 12532 417 12566 451
rect 12532 349 12566 383
rect 12532 299 12566 315
rect 12616 449 12667 465
rect 12650 415 12667 449
rect 12616 381 12667 415
rect 12650 347 12667 381
rect 12714 443 12731 477
rect 12714 409 12765 443
rect 12799 461 12865 527
rect 12799 427 12815 461
rect 12849 427 12865 461
rect 12899 477 12933 493
rect 12714 375 12731 409
rect 12899 409 12933 443
rect 12765 375 12864 393
rect 12714 359 12864 375
rect 12616 325 12667 347
rect 12616 289 12784 325
rect 12625 274 12784 289
rect 12419 249 12591 265
rect 12419 215 12557 249
rect 12419 199 12591 215
rect 12625 240 12656 274
rect 12694 249 12784 274
rect 12694 240 12728 249
rect 12625 215 12728 240
rect 12762 215 12784 249
rect 12419 119 12469 199
rect 12625 195 12784 215
rect 12818 264 12864 359
rect 12818 255 12830 264
rect 12852 221 12864 230
rect 12625 159 12667 195
rect 12818 161 12864 221
rect 12616 143 12667 159
rect 12419 85 12435 119
rect 12419 69 12469 85
rect 12532 113 12566 136
rect 12315 55 12381 63
rect 12532 17 12566 79
rect 12650 109 12667 143
rect 12616 53 12667 109
rect 12714 127 12864 161
rect 12714 119 12765 127
rect 12714 85 12731 119
rect 12899 119 12933 357
rect 12967 333 13032 490
rect 13066 485 13116 527
rect 13066 451 13082 485
rect 13066 435 13116 451
rect 13150 477 13200 493
rect 13150 443 13166 477
rect 13150 427 13200 443
rect 13243 483 13379 493
rect 13243 449 13259 483
rect 13293 449 13379 483
rect 13494 475 13560 527
rect 13687 485 13761 527
rect 13243 427 13379 449
rect 13150 401 13184 427
rect 13105 367 13184 401
rect 13218 391 13311 393
rect 12979 310 13071 333
rect 12979 276 13037 310
rect 12979 175 13071 276
rect 12979 141 13003 175
rect 13041 141 13071 175
rect 12979 123 13071 141
rect 12714 69 12765 85
rect 12799 59 12815 93
rect 12849 59 12865 93
rect 13105 95 13139 367
rect 13218 365 13277 391
rect 13252 357 13277 365
rect 13252 331 13311 357
rect 13218 315 13311 331
rect 13173 255 13243 277
rect 13173 221 13185 255
rect 13219 221 13243 255
rect 13173 203 13243 221
rect 13173 169 13196 203
rect 13230 169 13243 203
rect 13173 153 13243 169
rect 13277 197 13311 315
rect 13345 271 13379 427
rect 13413 459 13447 475
rect 13494 441 13510 475
rect 13544 441 13560 475
rect 13594 459 13628 475
rect 13413 407 13447 425
rect 13687 451 13707 485
rect 13741 451 13761 485
rect 13687 435 13761 451
rect 13795 477 13829 493
rect 13594 407 13628 425
rect 13413 373 13628 407
rect 13795 401 13829 443
rect 13876 484 14050 493
rect 13876 450 13892 484
rect 13926 450 14050 484
rect 13876 425 14050 450
rect 14084 485 14134 527
rect 14118 451 14134 485
rect 14238 485 14382 527
rect 14084 435 14134 451
rect 14168 459 14202 475
rect 13717 367 13829 401
rect 13717 339 13751 367
rect 13451 305 13467 339
rect 13501 305 13751 339
rect 13890 357 13901 391
rect 13935 365 13982 391
rect 13890 333 13932 357
rect 13345 251 13683 271
rect 13345 237 13649 251
rect 13277 163 13298 197
rect 13332 163 13348 197
rect 13277 153 13348 163
rect 13382 95 13416 237
rect 13457 187 13553 203
rect 13491 153 13529 187
rect 13587 169 13615 203
rect 13649 201 13683 217
rect 13563 153 13615 169
rect 13717 167 13751 305
rect 12899 69 12933 85
rect 12799 17 12865 59
rect 13005 55 13021 89
rect 13055 55 13071 89
rect 13105 61 13154 95
rect 13188 61 13204 95
rect 13245 61 13261 95
rect 13295 61 13416 95
rect 13591 93 13657 109
rect 13005 17 13071 55
rect 13591 59 13607 93
rect 13641 59 13657 93
rect 13591 17 13657 59
rect 13699 89 13751 167
rect 13789 331 13932 333
rect 13966 331 13982 365
rect 14016 349 14050 425
rect 14238 451 14254 485
rect 14288 451 14332 485
rect 14366 451 14382 485
rect 14416 477 14497 493
rect 14648 485 14682 527
rect 14168 417 14202 425
rect 14450 443 14497 477
rect 14168 383 14328 417
rect 13789 299 13924 331
rect 14016 315 14210 349
rect 14244 315 14260 349
rect 13789 191 13831 299
rect 14016 297 14050 315
rect 13789 157 13797 191
rect 13789 141 13831 157
rect 13865 255 13935 265
rect 13865 239 13901 255
rect 13865 205 13893 239
rect 13927 205 13935 221
rect 13865 141 13935 205
rect 13969 263 14050 297
rect 13969 107 14003 263
rect 14117 250 14225 281
rect 14294 265 14328 383
rect 14416 409 14497 443
rect 14450 375 14497 409
rect 14416 341 14497 375
rect 14450 307 14497 341
rect 14416 291 14497 307
rect 14294 259 14383 265
rect 14151 241 14225 250
rect 14037 213 14081 229
rect 14071 179 14081 213
rect 14117 207 14133 216
rect 14167 207 14225 241
rect 14037 173 14081 179
rect 14177 187 14225 207
rect 14037 139 14143 173
rect 13813 93 14003 107
rect 13699 55 13719 89
rect 13753 55 13769 89
rect 13813 59 13829 93
rect 13863 59 14003 93
rect 13813 51 14003 59
rect 14037 89 14075 105
rect 14037 55 14041 89
rect 14109 93 14143 139
rect 14211 153 14225 187
rect 14177 127 14225 153
rect 14259 249 14383 259
rect 14259 215 14333 249
rect 14367 215 14383 249
rect 14259 199 14383 215
rect 14259 164 14324 199
rect 14431 165 14497 291
rect 14259 109 14323 164
rect 14109 75 14259 93
rect 14293 75 14323 109
rect 14109 59 14323 75
rect 14363 132 14397 154
rect 14037 17 14075 55
rect 14363 17 14397 98
rect 14431 131 14447 165
rect 14481 131 14497 165
rect 14431 97 14497 131
rect 14431 63 14447 97
rect 14481 63 14497 97
rect 14535 451 14551 485
rect 14585 451 14601 485
rect 14535 417 14601 451
rect 14535 383 14551 417
rect 14585 383 14601 417
rect 14535 265 14601 383
rect 14830 477 14881 493
rect 14648 417 14682 451
rect 14648 349 14682 383
rect 14648 299 14682 315
rect 14732 449 14783 465
rect 14766 415 14783 449
rect 14732 381 14783 415
rect 14766 347 14783 381
rect 14830 443 14847 477
rect 14830 409 14881 443
rect 14915 461 14981 527
rect 14915 427 14931 461
rect 14965 427 14981 461
rect 15015 477 15049 493
rect 14830 375 14847 409
rect 15015 409 15049 443
rect 14881 375 14980 393
rect 14830 359 14980 375
rect 14732 325 14783 347
rect 14732 289 14900 325
rect 14741 274 14900 289
rect 14535 249 14707 265
rect 14535 215 14673 249
rect 14535 199 14707 215
rect 14741 240 14772 274
rect 14810 249 14900 274
rect 14810 240 14844 249
rect 14741 215 14844 240
rect 14878 215 14900 249
rect 14535 119 14585 199
rect 14741 195 14900 215
rect 14934 264 14980 359
rect 14934 255 14946 264
rect 14968 221 14980 230
rect 14741 159 14783 195
rect 14934 161 14980 221
rect 14732 143 14783 159
rect 14535 85 14551 119
rect 14535 69 14585 85
rect 14648 113 14682 136
rect 14431 55 14497 63
rect 14648 17 14682 79
rect 14766 109 14783 143
rect 14732 53 14783 109
rect 14830 127 14980 161
rect 14830 119 14881 127
rect 14830 85 14847 119
rect 15015 119 15049 357
rect 15083 333 15148 490
rect 15182 485 15232 527
rect 15182 451 15198 485
rect 15182 435 15232 451
rect 15266 477 15316 493
rect 15266 443 15282 477
rect 15266 427 15316 443
rect 15359 483 15495 493
rect 15359 449 15375 483
rect 15409 449 15495 483
rect 15610 475 15676 527
rect 15803 485 15877 527
rect 15359 427 15495 449
rect 15266 401 15300 427
rect 15221 367 15300 401
rect 15334 391 15427 393
rect 15095 310 15187 333
rect 15095 276 15153 310
rect 15095 175 15187 276
rect 15095 141 15119 175
rect 15157 141 15187 175
rect 15095 123 15187 141
rect 14830 69 14881 85
rect 14915 59 14931 93
rect 14965 59 14981 93
rect 15221 95 15255 367
rect 15334 365 15393 391
rect 15368 357 15393 365
rect 15368 331 15427 357
rect 15334 315 15427 331
rect 15289 255 15359 277
rect 15289 221 15301 255
rect 15335 221 15359 255
rect 15289 203 15359 221
rect 15289 169 15312 203
rect 15346 169 15359 203
rect 15289 153 15359 169
rect 15393 197 15427 315
rect 15461 271 15495 427
rect 15529 459 15563 475
rect 15610 441 15626 475
rect 15660 441 15676 475
rect 15710 459 15744 475
rect 15529 407 15563 425
rect 15803 451 15823 485
rect 15857 451 15877 485
rect 15803 435 15877 451
rect 15911 477 15945 493
rect 15710 407 15744 425
rect 15529 373 15744 407
rect 15911 401 15945 443
rect 15992 484 16166 493
rect 15992 450 16008 484
rect 16042 450 16166 484
rect 15992 425 16166 450
rect 16200 485 16250 527
rect 16234 451 16250 485
rect 16354 485 16498 527
rect 16200 435 16250 451
rect 16284 459 16318 475
rect 15833 367 15945 401
rect 15833 339 15867 367
rect 15567 305 15583 339
rect 15617 305 15867 339
rect 16006 357 16017 391
rect 16051 365 16098 391
rect 16006 333 16048 357
rect 15461 251 15799 271
rect 15461 237 15765 251
rect 15393 163 15414 197
rect 15448 163 15464 197
rect 15393 153 15464 163
rect 15498 95 15532 237
rect 15573 187 15669 203
rect 15607 153 15645 187
rect 15703 169 15731 203
rect 15765 201 15799 217
rect 15679 153 15731 169
rect 15833 167 15867 305
rect 15015 69 15049 85
rect 14915 17 14981 59
rect 15121 55 15137 89
rect 15171 55 15187 89
rect 15221 61 15270 95
rect 15304 61 15320 95
rect 15361 61 15377 95
rect 15411 61 15532 95
rect 15707 93 15773 109
rect 15121 17 15187 55
rect 15707 59 15723 93
rect 15757 59 15773 93
rect 15707 17 15773 59
rect 15815 89 15867 167
rect 15905 331 16048 333
rect 16082 331 16098 365
rect 16132 349 16166 425
rect 16354 451 16370 485
rect 16404 451 16448 485
rect 16482 451 16498 485
rect 16532 477 16613 493
rect 16764 485 16798 527
rect 16284 417 16318 425
rect 16566 443 16613 477
rect 16284 383 16444 417
rect 15905 299 16040 331
rect 16132 315 16326 349
rect 16360 315 16376 349
rect 15905 191 15947 299
rect 16132 297 16166 315
rect 15905 157 15913 191
rect 15905 141 15947 157
rect 15981 255 16051 265
rect 15981 239 16017 255
rect 15981 205 16009 239
rect 16043 205 16051 221
rect 15981 141 16051 205
rect 16085 263 16166 297
rect 16085 107 16119 263
rect 16233 250 16341 281
rect 16410 265 16444 383
rect 16532 409 16613 443
rect 16566 375 16613 409
rect 16532 341 16613 375
rect 16566 307 16613 341
rect 16532 291 16613 307
rect 16410 259 16499 265
rect 16267 241 16341 250
rect 16153 213 16197 229
rect 16187 179 16197 213
rect 16233 207 16249 216
rect 16283 207 16341 241
rect 16153 173 16197 179
rect 16293 187 16341 207
rect 16153 139 16259 173
rect 15929 93 16119 107
rect 15815 55 15835 89
rect 15869 55 15885 89
rect 15929 59 15945 93
rect 15979 59 16119 93
rect 15929 51 16119 59
rect 16153 89 16191 105
rect 16153 55 16157 89
rect 16225 93 16259 139
rect 16327 153 16341 187
rect 16293 127 16341 153
rect 16375 249 16499 259
rect 16375 215 16449 249
rect 16483 215 16499 249
rect 16375 199 16499 215
rect 16375 164 16440 199
rect 16547 165 16613 291
rect 16375 109 16439 164
rect 16225 75 16375 93
rect 16409 75 16439 109
rect 16225 59 16439 75
rect 16479 132 16513 154
rect 16153 17 16191 55
rect 16479 17 16513 98
rect 16547 131 16563 165
rect 16597 131 16613 165
rect 16547 97 16613 131
rect 16547 63 16563 97
rect 16597 63 16613 97
rect 16651 451 16667 485
rect 16701 451 16717 485
rect 16651 417 16717 451
rect 16651 383 16667 417
rect 16701 383 16717 417
rect 16651 265 16717 383
rect 16946 477 16997 493
rect 16764 417 16798 451
rect 16764 349 16798 383
rect 16764 299 16798 315
rect 16848 449 16899 465
rect 16882 415 16899 449
rect 16848 381 16899 415
rect 16882 347 16899 381
rect 16946 443 16963 477
rect 16946 409 16997 443
rect 17031 461 17097 527
rect 17031 427 17047 461
rect 17081 427 17097 461
rect 17131 477 17165 493
rect 16946 375 16963 409
rect 17131 409 17165 443
rect 16997 375 17096 393
rect 16946 359 17096 375
rect 16848 325 16899 347
rect 16848 289 17016 325
rect 16857 274 17016 289
rect 16651 249 16823 265
rect 16651 215 16789 249
rect 16651 199 16823 215
rect 16857 240 16888 274
rect 16926 249 17016 274
rect 16926 240 16960 249
rect 16857 215 16960 240
rect 16994 215 17016 249
rect 16651 119 16701 199
rect 16857 195 17016 215
rect 17050 264 17096 359
rect 17050 255 17062 264
rect 17084 221 17096 230
rect 16857 159 16899 195
rect 17050 161 17096 221
rect 16848 143 16899 159
rect 16651 85 16667 119
rect 16651 69 16701 85
rect 16764 113 16798 136
rect 16547 55 16613 63
rect 16764 17 16798 79
rect 16882 109 16899 143
rect 16848 53 16899 109
rect 16946 127 17096 161
rect 16946 119 16997 127
rect 16946 85 16963 119
rect 17131 119 17165 357
rect 17199 333 17264 490
rect 17298 485 17348 527
rect 17298 451 17314 485
rect 17298 435 17348 451
rect 17382 477 17432 493
rect 17382 443 17398 477
rect 17382 427 17432 443
rect 17475 483 17611 493
rect 17475 449 17491 483
rect 17525 449 17611 483
rect 17726 475 17792 527
rect 17919 485 17993 527
rect 17475 427 17611 449
rect 17382 401 17416 427
rect 17337 367 17416 401
rect 17450 391 17543 393
rect 17211 310 17303 333
rect 17211 276 17269 310
rect 17211 175 17303 276
rect 17211 141 17235 175
rect 17273 141 17303 175
rect 17211 123 17303 141
rect 16946 69 16997 85
rect 17031 59 17047 93
rect 17081 59 17097 93
rect 17337 95 17371 367
rect 17450 365 17509 391
rect 17484 357 17509 365
rect 17484 331 17543 357
rect 17450 315 17543 331
rect 17405 255 17475 277
rect 17405 221 17417 255
rect 17451 221 17475 255
rect 17405 203 17475 221
rect 17405 169 17428 203
rect 17462 169 17475 203
rect 17405 153 17475 169
rect 17509 197 17543 315
rect 17577 271 17611 427
rect 17645 459 17679 475
rect 17726 441 17742 475
rect 17776 441 17792 475
rect 17826 459 17860 475
rect 17645 407 17679 425
rect 17919 451 17939 485
rect 17973 451 17993 485
rect 17919 435 17993 451
rect 18027 477 18061 493
rect 17826 407 17860 425
rect 17645 373 17860 407
rect 18027 401 18061 443
rect 18108 484 18282 493
rect 18108 450 18124 484
rect 18158 450 18282 484
rect 18108 425 18282 450
rect 18316 485 18366 527
rect 18350 451 18366 485
rect 18470 485 18614 527
rect 18316 435 18366 451
rect 18400 459 18434 475
rect 17949 367 18061 401
rect 17949 339 17983 367
rect 17683 305 17699 339
rect 17733 305 17983 339
rect 18122 357 18133 391
rect 18167 365 18214 391
rect 18122 333 18164 357
rect 17577 251 17915 271
rect 17577 237 17881 251
rect 17509 163 17530 197
rect 17564 163 17580 197
rect 17509 153 17580 163
rect 17614 95 17648 237
rect 17689 187 17785 203
rect 17723 153 17761 187
rect 17819 169 17847 203
rect 17881 201 17915 217
rect 17795 153 17847 169
rect 17949 167 17983 305
rect 17131 69 17165 85
rect 17031 17 17097 59
rect 17237 55 17253 89
rect 17287 55 17303 89
rect 17337 61 17386 95
rect 17420 61 17436 95
rect 17477 61 17493 95
rect 17527 61 17648 95
rect 17823 93 17889 109
rect 17237 17 17303 55
rect 17823 59 17839 93
rect 17873 59 17889 93
rect 17823 17 17889 59
rect 17931 89 17983 167
rect 18021 331 18164 333
rect 18198 331 18214 365
rect 18248 349 18282 425
rect 18470 451 18486 485
rect 18520 451 18564 485
rect 18598 451 18614 485
rect 18648 477 18729 493
rect 18880 485 18914 527
rect 18400 417 18434 425
rect 18682 443 18729 477
rect 18400 383 18560 417
rect 18021 299 18156 331
rect 18248 315 18442 349
rect 18476 315 18492 349
rect 18021 191 18063 299
rect 18248 297 18282 315
rect 18021 157 18029 191
rect 18021 141 18063 157
rect 18097 255 18167 265
rect 18097 239 18133 255
rect 18097 205 18125 239
rect 18159 205 18167 221
rect 18097 141 18167 205
rect 18201 263 18282 297
rect 18201 107 18235 263
rect 18349 250 18457 281
rect 18526 265 18560 383
rect 18648 409 18729 443
rect 18682 375 18729 409
rect 18648 341 18729 375
rect 18682 307 18729 341
rect 18648 291 18729 307
rect 18526 259 18615 265
rect 18383 241 18457 250
rect 18269 213 18313 229
rect 18303 179 18313 213
rect 18349 207 18365 216
rect 18399 207 18457 241
rect 18269 173 18313 179
rect 18409 187 18457 207
rect 18269 139 18375 173
rect 18045 93 18235 107
rect 17931 55 17951 89
rect 17985 55 18001 89
rect 18045 59 18061 93
rect 18095 59 18235 93
rect 18045 51 18235 59
rect 18269 89 18307 105
rect 18269 55 18273 89
rect 18341 93 18375 139
rect 18443 153 18457 187
rect 18409 127 18457 153
rect 18491 249 18615 259
rect 18491 215 18565 249
rect 18599 215 18615 249
rect 18491 199 18615 215
rect 18491 164 18556 199
rect 18663 165 18729 291
rect 18491 109 18555 164
rect 18341 75 18491 93
rect 18525 75 18555 109
rect 18341 59 18555 75
rect 18595 132 18629 154
rect 18269 17 18307 55
rect 18595 17 18629 98
rect 18663 131 18679 165
rect 18713 131 18729 165
rect 18663 97 18729 131
rect 18663 63 18679 97
rect 18713 63 18729 97
rect 18767 451 18783 485
rect 18817 451 18833 485
rect 18767 417 18833 451
rect 18767 383 18783 417
rect 18817 383 18833 417
rect 18767 265 18833 383
rect 19062 477 19113 493
rect 18880 417 18914 451
rect 18880 349 18914 383
rect 18880 299 18914 315
rect 18964 449 19015 465
rect 18998 415 19015 449
rect 18964 381 19015 415
rect 18998 347 19015 381
rect 19062 443 19079 477
rect 19062 409 19113 443
rect 19147 461 19213 527
rect 19147 427 19163 461
rect 19197 427 19213 461
rect 19247 477 19281 493
rect 19062 375 19079 409
rect 19247 409 19281 443
rect 19113 375 19212 393
rect 19062 359 19212 375
rect 18964 325 19015 347
rect 18964 289 19132 325
rect 18973 274 19132 289
rect 18767 249 18939 265
rect 18767 215 18905 249
rect 18767 199 18939 215
rect 18973 240 19004 274
rect 19042 249 19132 274
rect 19042 240 19076 249
rect 18973 215 19076 240
rect 19110 215 19132 249
rect 18767 119 18817 199
rect 18973 195 19132 215
rect 19166 264 19212 359
rect 19166 255 19178 264
rect 19200 221 19212 230
rect 18973 159 19015 195
rect 19166 161 19212 221
rect 18964 143 19015 159
rect 18767 85 18783 119
rect 18767 69 18817 85
rect 18880 113 18914 136
rect 18663 55 18729 63
rect 18880 17 18914 79
rect 18998 109 19015 143
rect 18964 53 19015 109
rect 19062 127 19212 161
rect 19062 119 19113 127
rect 19062 85 19079 119
rect 19247 119 19281 357
rect 19315 333 19380 490
rect 19414 485 19464 527
rect 19414 451 19430 485
rect 19414 435 19464 451
rect 19498 477 19548 493
rect 19498 443 19514 477
rect 19498 427 19548 443
rect 19591 483 19727 493
rect 19591 449 19607 483
rect 19641 449 19727 483
rect 19842 475 19908 527
rect 20035 485 20109 527
rect 19591 427 19727 449
rect 19498 401 19532 427
rect 19453 367 19532 401
rect 19566 391 19659 393
rect 19327 310 19419 333
rect 19327 276 19385 310
rect 19327 175 19419 276
rect 19327 141 19351 175
rect 19389 141 19419 175
rect 19327 123 19419 141
rect 19062 69 19113 85
rect 19147 59 19163 93
rect 19197 59 19213 93
rect 19453 95 19487 367
rect 19566 365 19625 391
rect 19600 357 19625 365
rect 19600 331 19659 357
rect 19566 315 19659 331
rect 19521 255 19591 277
rect 19521 221 19533 255
rect 19567 221 19591 255
rect 19521 203 19591 221
rect 19521 169 19544 203
rect 19578 169 19591 203
rect 19521 153 19591 169
rect 19625 197 19659 315
rect 19693 271 19727 427
rect 19761 459 19795 475
rect 19842 441 19858 475
rect 19892 441 19908 475
rect 19942 459 19976 475
rect 19761 407 19795 425
rect 20035 451 20055 485
rect 20089 451 20109 485
rect 20035 435 20109 451
rect 20143 477 20177 493
rect 19942 407 19976 425
rect 19761 373 19976 407
rect 20143 401 20177 443
rect 20224 484 20398 493
rect 20224 450 20240 484
rect 20274 450 20398 484
rect 20224 425 20398 450
rect 20432 485 20482 527
rect 20466 451 20482 485
rect 20586 485 20730 527
rect 20432 435 20482 451
rect 20516 459 20550 475
rect 20065 367 20177 401
rect 20065 339 20099 367
rect 19799 305 19815 339
rect 19849 305 20099 339
rect 20238 357 20249 391
rect 20283 365 20330 391
rect 20238 333 20280 357
rect 19693 251 20031 271
rect 19693 237 19997 251
rect 19625 163 19646 197
rect 19680 163 19696 197
rect 19625 153 19696 163
rect 19730 95 19764 237
rect 19805 187 19901 203
rect 19839 153 19877 187
rect 19935 169 19963 203
rect 19997 201 20031 217
rect 19911 153 19963 169
rect 20065 167 20099 305
rect 19247 69 19281 85
rect 19147 17 19213 59
rect 19353 55 19369 89
rect 19403 55 19419 89
rect 19453 61 19502 95
rect 19536 61 19552 95
rect 19593 61 19609 95
rect 19643 61 19764 95
rect 19939 93 20005 109
rect 19353 17 19419 55
rect 19939 59 19955 93
rect 19989 59 20005 93
rect 19939 17 20005 59
rect 20047 89 20099 167
rect 20137 331 20280 333
rect 20314 331 20330 365
rect 20364 349 20398 425
rect 20586 451 20602 485
rect 20636 451 20680 485
rect 20714 451 20730 485
rect 20764 477 20845 493
rect 20996 485 21030 527
rect 20516 417 20550 425
rect 20798 443 20845 477
rect 20516 383 20676 417
rect 20137 299 20272 331
rect 20364 315 20558 349
rect 20592 315 20608 349
rect 20137 191 20179 299
rect 20364 297 20398 315
rect 20137 157 20145 191
rect 20137 141 20179 157
rect 20213 255 20283 265
rect 20213 239 20249 255
rect 20213 205 20241 239
rect 20275 205 20283 221
rect 20213 141 20283 205
rect 20317 263 20398 297
rect 20317 107 20351 263
rect 20465 250 20573 281
rect 20642 265 20676 383
rect 20764 409 20845 443
rect 20798 375 20845 409
rect 20764 341 20845 375
rect 20798 307 20845 341
rect 20764 291 20845 307
rect 20642 259 20731 265
rect 20499 241 20573 250
rect 20385 213 20429 229
rect 20419 179 20429 213
rect 20465 207 20481 216
rect 20515 207 20573 241
rect 20385 173 20429 179
rect 20525 187 20573 207
rect 20385 139 20491 173
rect 20161 93 20351 107
rect 20047 55 20067 89
rect 20101 55 20117 89
rect 20161 59 20177 93
rect 20211 59 20351 93
rect 20161 51 20351 59
rect 20385 89 20423 105
rect 20385 55 20389 89
rect 20457 93 20491 139
rect 20559 153 20573 187
rect 20525 127 20573 153
rect 20607 249 20731 259
rect 20607 215 20681 249
rect 20715 215 20731 249
rect 20607 199 20731 215
rect 20607 164 20672 199
rect 20779 165 20845 291
rect 20607 109 20671 164
rect 20457 75 20607 93
rect 20641 75 20671 109
rect 20457 59 20671 75
rect 20711 132 20745 154
rect 20385 17 20423 55
rect 20711 17 20745 98
rect 20779 131 20795 165
rect 20829 131 20845 165
rect 20779 97 20845 131
rect 20779 63 20795 97
rect 20829 63 20845 97
rect 20883 451 20899 485
rect 20933 451 20949 485
rect 20883 417 20949 451
rect 20883 383 20899 417
rect 20933 383 20949 417
rect 20883 265 20949 383
rect 21178 477 21229 493
rect 20996 417 21030 451
rect 20996 349 21030 383
rect 20996 299 21030 315
rect 21080 449 21131 465
rect 21114 415 21131 449
rect 21080 381 21131 415
rect 21114 347 21131 381
rect 21178 443 21195 477
rect 21178 409 21229 443
rect 21263 461 21329 527
rect 21263 427 21279 461
rect 21313 427 21329 461
rect 21363 477 21397 493
rect 21178 375 21195 409
rect 21363 409 21397 443
rect 21229 375 21328 393
rect 21178 359 21328 375
rect 21080 325 21131 347
rect 21080 289 21248 325
rect 21089 274 21248 289
rect 20883 249 21055 265
rect 20883 215 21021 249
rect 20883 199 21055 215
rect 21089 240 21120 274
rect 21158 249 21248 274
rect 21158 240 21192 249
rect 21089 215 21192 240
rect 21226 215 21248 249
rect 20883 119 20933 199
rect 21089 195 21248 215
rect 21282 264 21328 359
rect 21282 255 21294 264
rect 21316 221 21328 230
rect 21089 159 21131 195
rect 21282 161 21328 221
rect 21080 143 21131 159
rect 20883 85 20899 119
rect 20883 69 20933 85
rect 20996 113 21030 136
rect 20779 55 20845 63
rect 20996 17 21030 79
rect 21114 109 21131 143
rect 21080 53 21131 109
rect 21178 127 21328 161
rect 21178 119 21229 127
rect 21178 85 21195 119
rect 21363 119 21397 357
rect 21431 333 21496 490
rect 21530 485 21580 527
rect 21530 451 21546 485
rect 21530 435 21580 451
rect 21614 477 21664 493
rect 21614 443 21630 477
rect 21614 427 21664 443
rect 21707 483 21843 493
rect 21707 449 21723 483
rect 21757 449 21843 483
rect 21958 475 22024 527
rect 22151 485 22225 527
rect 21707 427 21843 449
rect 21614 401 21648 427
rect 21569 367 21648 401
rect 21682 391 21775 393
rect 21443 310 21535 333
rect 21443 276 21501 310
rect 21443 175 21535 276
rect 21443 141 21467 175
rect 21505 141 21535 175
rect 21443 123 21535 141
rect 21178 69 21229 85
rect 21263 59 21279 93
rect 21313 59 21329 93
rect 21569 95 21603 367
rect 21682 365 21741 391
rect 21716 357 21741 365
rect 21716 331 21775 357
rect 21682 315 21775 331
rect 21637 255 21707 277
rect 21637 221 21649 255
rect 21683 221 21707 255
rect 21637 203 21707 221
rect 21637 169 21660 203
rect 21694 169 21707 203
rect 21637 153 21707 169
rect 21741 197 21775 315
rect 21809 271 21843 427
rect 21877 459 21911 475
rect 21958 441 21974 475
rect 22008 441 22024 475
rect 22058 459 22092 475
rect 21877 407 21911 425
rect 22151 451 22171 485
rect 22205 451 22225 485
rect 22151 435 22225 451
rect 22259 477 22293 493
rect 22058 407 22092 425
rect 21877 373 22092 407
rect 22259 401 22293 443
rect 22340 484 22514 493
rect 22340 450 22356 484
rect 22390 450 22514 484
rect 22340 425 22514 450
rect 22548 485 22598 527
rect 22582 451 22598 485
rect 22702 485 22846 527
rect 22548 435 22598 451
rect 22632 459 22666 475
rect 22181 367 22293 401
rect 22181 339 22215 367
rect 21915 305 21931 339
rect 21965 305 22215 339
rect 22354 357 22365 391
rect 22399 365 22446 391
rect 22354 333 22396 357
rect 21809 251 22147 271
rect 21809 237 22113 251
rect 21741 163 21762 197
rect 21796 163 21812 197
rect 21741 153 21812 163
rect 21846 95 21880 237
rect 21921 187 22017 203
rect 21955 153 21993 187
rect 22051 169 22079 203
rect 22113 201 22147 217
rect 22027 153 22079 169
rect 22181 167 22215 305
rect 21363 69 21397 85
rect 21263 17 21329 59
rect 21469 55 21485 89
rect 21519 55 21535 89
rect 21569 61 21618 95
rect 21652 61 21668 95
rect 21709 61 21725 95
rect 21759 61 21880 95
rect 22055 93 22121 109
rect 21469 17 21535 55
rect 22055 59 22071 93
rect 22105 59 22121 93
rect 22055 17 22121 59
rect 22163 89 22215 167
rect 22253 331 22396 333
rect 22430 331 22446 365
rect 22480 349 22514 425
rect 22702 451 22718 485
rect 22752 451 22796 485
rect 22830 451 22846 485
rect 22880 477 22961 493
rect 23112 485 23146 527
rect 22632 417 22666 425
rect 22914 443 22961 477
rect 22632 383 22792 417
rect 22253 299 22388 331
rect 22480 315 22674 349
rect 22708 315 22724 349
rect 22253 191 22295 299
rect 22480 297 22514 315
rect 22253 157 22261 191
rect 22253 141 22295 157
rect 22329 255 22399 265
rect 22329 239 22365 255
rect 22329 205 22357 239
rect 22391 205 22399 221
rect 22329 141 22399 205
rect 22433 263 22514 297
rect 22433 107 22467 263
rect 22581 250 22689 281
rect 22758 265 22792 383
rect 22880 409 22961 443
rect 22914 375 22961 409
rect 22880 341 22961 375
rect 22914 307 22961 341
rect 22880 291 22961 307
rect 22758 259 22847 265
rect 22615 241 22689 250
rect 22501 213 22545 229
rect 22535 179 22545 213
rect 22581 207 22597 216
rect 22631 207 22689 241
rect 22501 173 22545 179
rect 22641 187 22689 207
rect 22501 139 22607 173
rect 22277 93 22467 107
rect 22163 55 22183 89
rect 22217 55 22233 89
rect 22277 59 22293 93
rect 22327 59 22467 93
rect 22277 51 22467 59
rect 22501 89 22539 105
rect 22501 55 22505 89
rect 22573 93 22607 139
rect 22675 153 22689 187
rect 22641 127 22689 153
rect 22723 249 22847 259
rect 22723 215 22797 249
rect 22831 215 22847 249
rect 22723 199 22847 215
rect 22723 164 22788 199
rect 22895 165 22961 291
rect 22723 109 22787 164
rect 22573 75 22723 93
rect 22757 75 22787 109
rect 22573 59 22787 75
rect 22827 132 22861 154
rect 22501 17 22539 55
rect 22827 17 22861 98
rect 22895 131 22911 165
rect 22945 131 22961 165
rect 22895 97 22961 131
rect 22895 63 22911 97
rect 22945 63 22961 97
rect 22999 451 23015 485
rect 23049 451 23065 485
rect 22999 417 23065 451
rect 22999 383 23015 417
rect 23049 383 23065 417
rect 22999 265 23065 383
rect 23294 477 23345 493
rect 23112 417 23146 451
rect 23112 349 23146 383
rect 23112 299 23146 315
rect 23196 449 23247 465
rect 23230 415 23247 449
rect 23196 381 23247 415
rect 23230 347 23247 381
rect 23294 443 23311 477
rect 23294 409 23345 443
rect 23379 461 23445 527
rect 23379 427 23395 461
rect 23429 427 23445 461
rect 23479 477 23513 493
rect 23294 375 23311 409
rect 23479 409 23513 443
rect 23345 375 23444 393
rect 23294 359 23444 375
rect 23196 325 23247 347
rect 23196 289 23364 325
rect 23205 274 23364 289
rect 22999 249 23171 265
rect 22999 215 23137 249
rect 22999 199 23171 215
rect 23205 240 23236 274
rect 23274 249 23364 274
rect 23274 240 23308 249
rect 23205 215 23308 240
rect 23342 215 23364 249
rect 22999 119 23049 199
rect 23205 195 23364 215
rect 23398 264 23444 359
rect 23398 255 23410 264
rect 23432 221 23444 230
rect 23205 159 23247 195
rect 23398 161 23444 221
rect 23196 143 23247 159
rect 22999 85 23015 119
rect 22999 69 23049 85
rect 23112 113 23146 136
rect 22895 55 22961 63
rect 23112 17 23146 79
rect 23230 109 23247 143
rect 23196 53 23247 109
rect 23294 127 23444 161
rect 23294 119 23345 127
rect 23294 85 23311 119
rect 23479 119 23513 357
rect 23547 333 23612 490
rect 23646 485 23696 527
rect 23646 451 23662 485
rect 23646 435 23696 451
rect 23730 477 23780 493
rect 23730 443 23746 477
rect 23730 427 23780 443
rect 23823 483 23959 493
rect 23823 449 23839 483
rect 23873 449 23959 483
rect 24074 475 24140 527
rect 24267 485 24341 527
rect 23823 427 23959 449
rect 23730 401 23764 427
rect 23685 367 23764 401
rect 23798 391 23891 393
rect 23559 310 23651 333
rect 23559 276 23617 310
rect 23559 175 23651 276
rect 23559 141 23583 175
rect 23621 141 23651 175
rect 23559 123 23651 141
rect 23294 69 23345 85
rect 23379 59 23395 93
rect 23429 59 23445 93
rect 23685 95 23719 367
rect 23798 365 23857 391
rect 23832 357 23857 365
rect 23832 331 23891 357
rect 23798 315 23891 331
rect 23753 255 23823 277
rect 23753 221 23765 255
rect 23799 221 23823 255
rect 23753 203 23823 221
rect 23753 169 23776 203
rect 23810 169 23823 203
rect 23753 153 23823 169
rect 23857 197 23891 315
rect 23925 271 23959 427
rect 23993 459 24027 475
rect 24074 441 24090 475
rect 24124 441 24140 475
rect 24174 459 24208 475
rect 23993 407 24027 425
rect 24267 451 24287 485
rect 24321 451 24341 485
rect 24267 435 24341 451
rect 24375 477 24409 493
rect 24174 407 24208 425
rect 23993 373 24208 407
rect 24375 401 24409 443
rect 24456 484 24630 493
rect 24456 450 24472 484
rect 24506 450 24630 484
rect 24456 425 24630 450
rect 24664 485 24714 527
rect 24698 451 24714 485
rect 24818 485 24962 527
rect 24664 435 24714 451
rect 24748 459 24782 475
rect 24297 367 24409 401
rect 24297 339 24331 367
rect 24031 305 24047 339
rect 24081 305 24331 339
rect 24470 357 24481 391
rect 24515 365 24562 391
rect 24470 333 24512 357
rect 23925 251 24263 271
rect 23925 237 24229 251
rect 23857 163 23878 197
rect 23912 163 23928 197
rect 23857 153 23928 163
rect 23962 95 23996 237
rect 24037 187 24133 203
rect 24071 153 24109 187
rect 24167 169 24195 203
rect 24229 201 24263 217
rect 24143 153 24195 169
rect 24297 167 24331 305
rect 23479 69 23513 85
rect 23379 17 23445 59
rect 23585 55 23601 89
rect 23635 55 23651 89
rect 23685 61 23734 95
rect 23768 61 23784 95
rect 23825 61 23841 95
rect 23875 61 23996 95
rect 24171 93 24237 109
rect 23585 17 23651 55
rect 24171 59 24187 93
rect 24221 59 24237 93
rect 24171 17 24237 59
rect 24279 89 24331 167
rect 24369 331 24512 333
rect 24546 331 24562 365
rect 24596 349 24630 425
rect 24818 451 24834 485
rect 24868 451 24912 485
rect 24946 451 24962 485
rect 24996 477 25077 493
rect 25228 485 25262 527
rect 24748 417 24782 425
rect 25030 443 25077 477
rect 24748 383 24908 417
rect 24369 299 24504 331
rect 24596 315 24790 349
rect 24824 315 24840 349
rect 24369 191 24411 299
rect 24596 297 24630 315
rect 24369 157 24377 191
rect 24369 141 24411 157
rect 24445 255 24515 265
rect 24445 239 24481 255
rect 24445 205 24473 239
rect 24507 205 24515 221
rect 24445 141 24515 205
rect 24549 263 24630 297
rect 24549 107 24583 263
rect 24697 250 24805 281
rect 24874 265 24908 383
rect 24996 409 25077 443
rect 25030 375 25077 409
rect 24996 341 25077 375
rect 25030 307 25077 341
rect 24996 291 25077 307
rect 24874 259 24963 265
rect 24731 241 24805 250
rect 24617 213 24661 229
rect 24651 179 24661 213
rect 24697 207 24713 216
rect 24747 207 24805 241
rect 24617 173 24661 179
rect 24757 187 24805 207
rect 24617 139 24723 173
rect 24393 93 24583 107
rect 24279 55 24299 89
rect 24333 55 24349 89
rect 24393 59 24409 93
rect 24443 59 24583 93
rect 24393 51 24583 59
rect 24617 89 24655 105
rect 24617 55 24621 89
rect 24689 93 24723 139
rect 24791 153 24805 187
rect 24757 127 24805 153
rect 24839 249 24963 259
rect 24839 215 24913 249
rect 24947 215 24963 249
rect 24839 199 24963 215
rect 24839 164 24904 199
rect 25011 165 25077 291
rect 24839 109 24903 164
rect 24689 75 24839 93
rect 24873 75 24903 109
rect 24689 59 24903 75
rect 24943 132 24977 154
rect 24617 17 24655 55
rect 24943 17 24977 98
rect 25011 131 25027 165
rect 25061 131 25077 165
rect 25011 97 25077 131
rect 25011 63 25027 97
rect 25061 63 25077 97
rect 25115 451 25131 485
rect 25165 451 25181 485
rect 25115 417 25181 451
rect 25115 383 25131 417
rect 25165 383 25181 417
rect 25115 265 25181 383
rect 25410 477 25461 493
rect 25228 417 25262 451
rect 25228 349 25262 383
rect 25228 299 25262 315
rect 25312 449 25363 465
rect 25346 415 25363 449
rect 25312 381 25363 415
rect 25346 347 25363 381
rect 25410 443 25427 477
rect 25410 409 25461 443
rect 25495 461 25561 527
rect 25495 427 25511 461
rect 25545 427 25561 461
rect 25595 477 25629 493
rect 25410 375 25427 409
rect 25595 409 25629 443
rect 25461 375 25560 393
rect 25410 359 25560 375
rect 25312 325 25363 347
rect 25312 289 25480 325
rect 25321 274 25480 289
rect 25115 249 25287 265
rect 25115 215 25253 249
rect 25115 199 25287 215
rect 25321 240 25352 274
rect 25390 249 25480 274
rect 25390 240 25424 249
rect 25321 215 25424 240
rect 25458 215 25480 249
rect 25115 119 25165 199
rect 25321 195 25480 215
rect 25514 264 25560 359
rect 25514 255 25526 264
rect 25548 221 25560 230
rect 25321 159 25363 195
rect 25514 161 25560 221
rect 25312 143 25363 159
rect 25115 85 25131 119
rect 25115 69 25165 85
rect 25228 113 25262 136
rect 25011 55 25077 63
rect 25228 17 25262 79
rect 25346 109 25363 143
rect 25312 53 25363 109
rect 25410 127 25560 161
rect 25410 119 25461 127
rect 25410 85 25427 119
rect 25595 119 25629 357
rect 25663 333 25728 490
rect 25762 485 25812 527
rect 25762 451 25778 485
rect 25762 435 25812 451
rect 25846 477 25896 493
rect 25846 443 25862 477
rect 25846 427 25896 443
rect 25939 483 26075 493
rect 25939 449 25955 483
rect 25989 449 26075 483
rect 26190 475 26256 527
rect 26383 485 26457 527
rect 25939 427 26075 449
rect 25846 401 25880 427
rect 25801 367 25880 401
rect 25914 391 26007 393
rect 25675 310 25767 333
rect 25675 276 25733 310
rect 25675 175 25767 276
rect 25675 141 25699 175
rect 25737 141 25767 175
rect 25675 123 25767 141
rect 25410 69 25461 85
rect 25495 59 25511 93
rect 25545 59 25561 93
rect 25801 95 25835 367
rect 25914 365 25973 391
rect 25948 357 25973 365
rect 25948 331 26007 357
rect 25914 315 26007 331
rect 25869 255 25939 277
rect 25869 221 25881 255
rect 25915 221 25939 255
rect 25869 203 25939 221
rect 25869 169 25892 203
rect 25926 169 25939 203
rect 25869 153 25939 169
rect 25973 197 26007 315
rect 26041 271 26075 427
rect 26109 459 26143 475
rect 26190 441 26206 475
rect 26240 441 26256 475
rect 26290 459 26324 475
rect 26109 407 26143 425
rect 26383 451 26403 485
rect 26437 451 26457 485
rect 26383 435 26457 451
rect 26491 477 26525 493
rect 26290 407 26324 425
rect 26109 373 26324 407
rect 26491 401 26525 443
rect 26572 484 26746 493
rect 26572 450 26588 484
rect 26622 450 26746 484
rect 26572 425 26746 450
rect 26780 485 26830 527
rect 26814 451 26830 485
rect 26934 485 27078 527
rect 26780 435 26830 451
rect 26864 459 26898 475
rect 26413 367 26525 401
rect 26413 339 26447 367
rect 26147 305 26163 339
rect 26197 305 26447 339
rect 26586 357 26597 391
rect 26631 365 26678 391
rect 26586 333 26628 357
rect 26041 251 26379 271
rect 26041 237 26345 251
rect 25973 163 25994 197
rect 26028 163 26044 197
rect 25973 153 26044 163
rect 26078 95 26112 237
rect 26153 187 26249 203
rect 26187 153 26225 187
rect 26283 169 26311 203
rect 26345 201 26379 217
rect 26259 153 26311 169
rect 26413 167 26447 305
rect 25595 69 25629 85
rect 25495 17 25561 59
rect 25701 55 25717 89
rect 25751 55 25767 89
rect 25801 61 25850 95
rect 25884 61 25900 95
rect 25941 61 25957 95
rect 25991 61 26112 95
rect 26287 93 26353 109
rect 25701 17 25767 55
rect 26287 59 26303 93
rect 26337 59 26353 93
rect 26287 17 26353 59
rect 26395 89 26447 167
rect 26485 331 26628 333
rect 26662 331 26678 365
rect 26712 349 26746 425
rect 26934 451 26950 485
rect 26984 451 27028 485
rect 27062 451 27078 485
rect 27112 477 27193 493
rect 27344 485 27378 527
rect 26864 417 26898 425
rect 27146 443 27193 477
rect 26864 383 27024 417
rect 26485 299 26620 331
rect 26712 315 26906 349
rect 26940 315 26956 349
rect 26485 191 26527 299
rect 26712 297 26746 315
rect 26485 157 26493 191
rect 26485 141 26527 157
rect 26561 255 26631 265
rect 26561 239 26597 255
rect 26561 205 26589 239
rect 26623 205 26631 221
rect 26561 141 26631 205
rect 26665 263 26746 297
rect 26665 107 26699 263
rect 26813 250 26921 281
rect 26990 265 27024 383
rect 27112 409 27193 443
rect 27146 375 27193 409
rect 27112 341 27193 375
rect 27146 307 27193 341
rect 27112 291 27193 307
rect 26990 259 27079 265
rect 26847 241 26921 250
rect 26733 213 26777 229
rect 26767 179 26777 213
rect 26813 207 26829 216
rect 26863 207 26921 241
rect 26733 173 26777 179
rect 26873 187 26921 207
rect 26733 139 26839 173
rect 26509 93 26699 107
rect 26395 55 26415 89
rect 26449 55 26465 89
rect 26509 59 26525 93
rect 26559 59 26699 93
rect 26509 51 26699 59
rect 26733 89 26771 105
rect 26733 55 26737 89
rect 26805 93 26839 139
rect 26907 153 26921 187
rect 26873 127 26921 153
rect 26955 249 27079 259
rect 26955 215 27029 249
rect 27063 215 27079 249
rect 26955 199 27079 215
rect 26955 164 27020 199
rect 27127 165 27193 291
rect 26955 109 27019 164
rect 26805 75 26955 93
rect 26989 75 27019 109
rect 26805 59 27019 75
rect 27059 132 27093 154
rect 26733 17 26771 55
rect 27059 17 27093 98
rect 27127 131 27143 165
rect 27177 131 27193 165
rect 27127 97 27193 131
rect 27127 63 27143 97
rect 27177 63 27193 97
rect 27231 451 27247 485
rect 27281 451 27297 485
rect 27231 417 27297 451
rect 27231 383 27247 417
rect 27281 383 27297 417
rect 27231 265 27297 383
rect 27526 477 27577 493
rect 27344 417 27378 451
rect 27344 349 27378 383
rect 27344 299 27378 315
rect 27428 449 27479 465
rect 27462 415 27479 449
rect 27428 381 27479 415
rect 27462 347 27479 381
rect 27526 443 27543 477
rect 27526 409 27577 443
rect 27611 461 27677 527
rect 27611 427 27627 461
rect 27661 427 27677 461
rect 27711 477 27745 493
rect 27526 375 27543 409
rect 27711 409 27745 443
rect 27577 375 27676 393
rect 27526 359 27676 375
rect 27428 325 27479 347
rect 27428 289 27596 325
rect 27437 274 27596 289
rect 27231 249 27403 265
rect 27231 215 27369 249
rect 27231 199 27403 215
rect 27437 240 27468 274
rect 27506 249 27596 274
rect 27506 240 27540 249
rect 27437 215 27540 240
rect 27574 215 27596 249
rect 27231 119 27281 199
rect 27437 195 27596 215
rect 27630 264 27676 359
rect 27630 255 27642 264
rect 27664 221 27676 230
rect 27437 159 27479 195
rect 27630 161 27676 221
rect 27428 143 27479 159
rect 27231 85 27247 119
rect 27231 69 27281 85
rect 27344 113 27378 136
rect 27127 55 27193 63
rect 27344 17 27378 79
rect 27462 109 27479 143
rect 27428 53 27479 109
rect 27526 127 27676 161
rect 27526 119 27577 127
rect 27526 85 27543 119
rect 27711 119 27745 357
rect 27779 333 27844 490
rect 27878 485 27928 527
rect 27878 451 27894 485
rect 27878 435 27928 451
rect 27962 477 28012 493
rect 27962 443 27978 477
rect 27962 427 28012 443
rect 28055 483 28191 493
rect 28055 449 28071 483
rect 28105 449 28191 483
rect 28306 475 28372 527
rect 28499 485 28573 527
rect 28055 427 28191 449
rect 27962 401 27996 427
rect 27917 367 27996 401
rect 28030 391 28123 393
rect 27791 310 27883 333
rect 27791 276 27849 310
rect 27791 175 27883 276
rect 27791 141 27815 175
rect 27853 141 27883 175
rect 27791 123 27883 141
rect 27526 69 27577 85
rect 27611 59 27627 93
rect 27661 59 27677 93
rect 27917 95 27951 367
rect 28030 365 28089 391
rect 28064 357 28089 365
rect 28064 331 28123 357
rect 28030 315 28123 331
rect 27985 255 28055 277
rect 27985 221 27997 255
rect 28031 221 28055 255
rect 27985 203 28055 221
rect 27985 169 28008 203
rect 28042 169 28055 203
rect 27985 153 28055 169
rect 28089 197 28123 315
rect 28157 271 28191 427
rect 28225 459 28259 475
rect 28306 441 28322 475
rect 28356 441 28372 475
rect 28406 459 28440 475
rect 28225 407 28259 425
rect 28499 451 28519 485
rect 28553 451 28573 485
rect 28499 435 28573 451
rect 28607 477 28641 493
rect 28406 407 28440 425
rect 28225 373 28440 407
rect 28607 401 28641 443
rect 28688 484 28862 493
rect 28688 450 28704 484
rect 28738 450 28862 484
rect 28688 425 28862 450
rect 28896 485 28946 527
rect 28930 451 28946 485
rect 29050 485 29194 527
rect 28896 435 28946 451
rect 28980 459 29014 475
rect 28529 367 28641 401
rect 28529 339 28563 367
rect 28263 305 28279 339
rect 28313 305 28563 339
rect 28702 357 28713 391
rect 28747 365 28794 391
rect 28702 333 28744 357
rect 28157 251 28495 271
rect 28157 237 28461 251
rect 28089 163 28110 197
rect 28144 163 28160 197
rect 28089 153 28160 163
rect 28194 95 28228 237
rect 28269 187 28365 203
rect 28303 153 28341 187
rect 28399 169 28427 203
rect 28461 201 28495 217
rect 28375 153 28427 169
rect 28529 167 28563 305
rect 27711 69 27745 85
rect 27611 17 27677 59
rect 27817 55 27833 89
rect 27867 55 27883 89
rect 27917 61 27966 95
rect 28000 61 28016 95
rect 28057 61 28073 95
rect 28107 61 28228 95
rect 28403 93 28469 109
rect 27817 17 27883 55
rect 28403 59 28419 93
rect 28453 59 28469 93
rect 28403 17 28469 59
rect 28511 89 28563 167
rect 28601 331 28744 333
rect 28778 331 28794 365
rect 28828 349 28862 425
rect 29050 451 29066 485
rect 29100 451 29144 485
rect 29178 451 29194 485
rect 29228 477 29309 493
rect 29460 485 29494 527
rect 28980 417 29014 425
rect 29262 443 29309 477
rect 28980 383 29140 417
rect 28601 299 28736 331
rect 28828 315 29022 349
rect 29056 315 29072 349
rect 28601 191 28643 299
rect 28828 297 28862 315
rect 28601 157 28609 191
rect 28601 141 28643 157
rect 28677 255 28747 265
rect 28677 239 28713 255
rect 28677 205 28705 239
rect 28739 205 28747 221
rect 28677 141 28747 205
rect 28781 263 28862 297
rect 28781 107 28815 263
rect 28929 250 29037 281
rect 29106 265 29140 383
rect 29228 409 29309 443
rect 29262 375 29309 409
rect 29228 341 29309 375
rect 29262 307 29309 341
rect 29228 291 29309 307
rect 29106 259 29195 265
rect 28963 241 29037 250
rect 28849 213 28893 229
rect 28883 179 28893 213
rect 28929 207 28945 216
rect 28979 207 29037 241
rect 28849 173 28893 179
rect 28989 187 29037 207
rect 28849 139 28955 173
rect 28625 93 28815 107
rect 28511 55 28531 89
rect 28565 55 28581 89
rect 28625 59 28641 93
rect 28675 59 28815 93
rect 28625 51 28815 59
rect 28849 89 28887 105
rect 28849 55 28853 89
rect 28921 93 28955 139
rect 29023 153 29037 187
rect 28989 127 29037 153
rect 29071 249 29195 259
rect 29071 215 29145 249
rect 29179 215 29195 249
rect 29071 199 29195 215
rect 29071 164 29136 199
rect 29243 165 29309 291
rect 29071 109 29135 164
rect 28921 75 29071 93
rect 29105 75 29135 109
rect 28921 59 29135 75
rect 29175 132 29209 154
rect 28849 17 28887 55
rect 29175 17 29209 98
rect 29243 131 29259 165
rect 29293 131 29309 165
rect 29243 97 29309 131
rect 29243 63 29259 97
rect 29293 63 29309 97
rect 29347 451 29363 485
rect 29397 451 29413 485
rect 29347 417 29413 451
rect 29347 383 29363 417
rect 29397 383 29413 417
rect 29347 265 29413 383
rect 29642 477 29693 493
rect 29460 417 29494 451
rect 29460 349 29494 383
rect 29460 299 29494 315
rect 29544 449 29595 465
rect 29578 415 29595 449
rect 29544 381 29595 415
rect 29578 347 29595 381
rect 29642 443 29659 477
rect 29642 409 29693 443
rect 29727 461 29793 527
rect 29727 427 29743 461
rect 29777 427 29793 461
rect 29827 477 29861 493
rect 29642 375 29659 409
rect 29827 409 29861 443
rect 29693 375 29792 393
rect 29642 359 29792 375
rect 29544 325 29595 347
rect 29544 289 29712 325
rect 29553 274 29712 289
rect 29347 249 29519 265
rect 29347 215 29485 249
rect 29347 199 29519 215
rect 29553 240 29584 274
rect 29622 249 29712 274
rect 29622 240 29656 249
rect 29553 215 29656 240
rect 29690 215 29712 249
rect 29347 119 29397 199
rect 29553 195 29712 215
rect 29746 264 29792 359
rect 29746 255 29758 264
rect 29780 221 29792 230
rect 29553 159 29595 195
rect 29746 161 29792 221
rect 29544 143 29595 159
rect 29347 85 29363 119
rect 29347 69 29397 85
rect 29460 113 29494 136
rect 29243 55 29309 63
rect 29460 17 29494 79
rect 29578 109 29595 143
rect 29544 53 29595 109
rect 29642 127 29792 161
rect 29642 119 29693 127
rect 29642 85 29659 119
rect 29827 119 29861 357
rect 29895 333 29960 490
rect 29994 485 30044 527
rect 29994 451 30010 485
rect 29994 435 30044 451
rect 30078 477 30128 493
rect 30078 443 30094 477
rect 30078 427 30128 443
rect 30171 483 30307 493
rect 30171 449 30187 483
rect 30221 449 30307 483
rect 30422 475 30488 527
rect 30615 485 30689 527
rect 30171 427 30307 449
rect 30078 401 30112 427
rect 30033 367 30112 401
rect 30146 391 30239 393
rect 29907 310 29999 333
rect 29907 276 29965 310
rect 29907 175 29999 276
rect 29907 141 29931 175
rect 29969 141 29999 175
rect 29907 123 29999 141
rect 29642 69 29693 85
rect 29727 59 29743 93
rect 29777 59 29793 93
rect 30033 95 30067 367
rect 30146 365 30205 391
rect 30180 357 30205 365
rect 30180 331 30239 357
rect 30146 315 30239 331
rect 30101 255 30171 277
rect 30101 221 30113 255
rect 30147 221 30171 255
rect 30101 203 30171 221
rect 30101 169 30124 203
rect 30158 169 30171 203
rect 30101 153 30171 169
rect 30205 197 30239 315
rect 30273 271 30307 427
rect 30341 459 30375 475
rect 30422 441 30438 475
rect 30472 441 30488 475
rect 30522 459 30556 475
rect 30341 407 30375 425
rect 30615 451 30635 485
rect 30669 451 30689 485
rect 30615 435 30689 451
rect 30723 477 30757 493
rect 30522 407 30556 425
rect 30341 373 30556 407
rect 30723 401 30757 443
rect 30804 484 30978 493
rect 30804 450 30820 484
rect 30854 450 30978 484
rect 30804 425 30978 450
rect 31012 485 31062 527
rect 31046 451 31062 485
rect 31166 485 31310 527
rect 31012 435 31062 451
rect 31096 459 31130 475
rect 30645 367 30757 401
rect 30645 339 30679 367
rect 30379 305 30395 339
rect 30429 305 30679 339
rect 30818 357 30829 391
rect 30863 365 30910 391
rect 30818 333 30860 357
rect 30273 251 30611 271
rect 30273 237 30577 251
rect 30205 163 30226 197
rect 30260 163 30276 197
rect 30205 153 30276 163
rect 30310 95 30344 237
rect 30385 187 30481 203
rect 30419 153 30457 187
rect 30515 169 30543 203
rect 30577 201 30611 217
rect 30491 153 30543 169
rect 30645 167 30679 305
rect 29827 69 29861 85
rect 29727 17 29793 59
rect 29933 55 29949 89
rect 29983 55 29999 89
rect 30033 61 30082 95
rect 30116 61 30132 95
rect 30173 61 30189 95
rect 30223 61 30344 95
rect 30519 93 30585 109
rect 29933 17 29999 55
rect 30519 59 30535 93
rect 30569 59 30585 93
rect 30519 17 30585 59
rect 30627 89 30679 167
rect 30717 331 30860 333
rect 30894 331 30910 365
rect 30944 349 30978 425
rect 31166 451 31182 485
rect 31216 451 31260 485
rect 31294 451 31310 485
rect 31344 477 31425 493
rect 31576 485 31610 527
rect 31096 417 31130 425
rect 31378 443 31425 477
rect 31096 383 31256 417
rect 30717 299 30852 331
rect 30944 315 31138 349
rect 31172 315 31188 349
rect 30717 191 30759 299
rect 30944 297 30978 315
rect 30717 157 30725 191
rect 30717 141 30759 157
rect 30793 255 30863 265
rect 30793 239 30829 255
rect 30793 205 30821 239
rect 30855 205 30863 221
rect 30793 141 30863 205
rect 30897 263 30978 297
rect 30897 107 30931 263
rect 31045 250 31153 281
rect 31222 265 31256 383
rect 31344 409 31425 443
rect 31378 375 31425 409
rect 31344 341 31425 375
rect 31378 307 31425 341
rect 31344 291 31425 307
rect 31222 259 31311 265
rect 31079 241 31153 250
rect 30965 213 31009 229
rect 30999 179 31009 213
rect 31045 207 31061 216
rect 31095 207 31153 241
rect 30965 173 31009 179
rect 31105 187 31153 207
rect 30965 139 31071 173
rect 30741 93 30931 107
rect 30627 55 30647 89
rect 30681 55 30697 89
rect 30741 59 30757 93
rect 30791 59 30931 93
rect 30741 51 30931 59
rect 30965 89 31003 105
rect 30965 55 30969 89
rect 31037 93 31071 139
rect 31139 153 31153 187
rect 31105 127 31153 153
rect 31187 249 31311 259
rect 31187 215 31261 249
rect 31295 215 31311 249
rect 31187 199 31311 215
rect 31187 164 31252 199
rect 31359 165 31425 291
rect 31187 109 31251 164
rect 31037 75 31187 93
rect 31221 75 31251 109
rect 31037 59 31251 75
rect 31291 132 31325 154
rect 30965 17 31003 55
rect 31291 17 31325 98
rect 31359 131 31375 165
rect 31409 131 31425 165
rect 31359 97 31425 131
rect 31359 63 31375 97
rect 31409 63 31425 97
rect 31463 451 31479 485
rect 31513 451 31529 485
rect 31463 417 31529 451
rect 31463 383 31479 417
rect 31513 383 31529 417
rect 31463 265 31529 383
rect 31758 477 31809 493
rect 31576 417 31610 451
rect 31576 349 31610 383
rect 31576 299 31610 315
rect 31660 449 31711 465
rect 31694 415 31711 449
rect 31660 381 31711 415
rect 31694 347 31711 381
rect 31758 443 31775 477
rect 31758 409 31809 443
rect 31843 461 31909 527
rect 31843 427 31859 461
rect 31893 427 31909 461
rect 31943 477 31977 493
rect 31758 375 31775 409
rect 31943 409 31977 443
rect 31809 375 31908 393
rect 31758 359 31908 375
rect 31660 325 31711 347
rect 31660 289 31828 325
rect 31669 274 31828 289
rect 31463 249 31635 265
rect 31463 215 31601 249
rect 31463 199 31635 215
rect 31669 240 31700 274
rect 31738 249 31828 274
rect 31738 240 31772 249
rect 31669 215 31772 240
rect 31806 215 31828 249
rect 31463 119 31513 199
rect 31669 195 31828 215
rect 31862 264 31908 359
rect 31862 255 31874 264
rect 31896 221 31908 230
rect 31669 159 31711 195
rect 31862 161 31908 221
rect 31660 143 31711 159
rect 31463 85 31479 119
rect 31463 69 31513 85
rect 31576 113 31610 136
rect 31359 55 31425 63
rect 31576 17 31610 79
rect 31694 109 31711 143
rect 31660 53 31711 109
rect 31758 127 31908 161
rect 31758 119 31809 127
rect 31758 85 31775 119
rect 31943 119 31977 357
rect 32011 333 32076 490
rect 32110 485 32160 527
rect 32110 451 32126 485
rect 32110 435 32160 451
rect 32194 477 32244 493
rect 32194 443 32210 477
rect 32194 427 32244 443
rect 32287 483 32423 493
rect 32287 449 32303 483
rect 32337 449 32423 483
rect 32538 475 32604 527
rect 32731 485 32805 527
rect 32287 427 32423 449
rect 32194 401 32228 427
rect 32149 367 32228 401
rect 32262 391 32355 393
rect 32023 310 32115 333
rect 32023 276 32081 310
rect 32023 175 32115 276
rect 32023 141 32047 175
rect 32085 141 32115 175
rect 32023 123 32115 141
rect 31758 69 31809 85
rect 31843 59 31859 93
rect 31893 59 31909 93
rect 32149 95 32183 367
rect 32262 365 32321 391
rect 32296 357 32321 365
rect 32296 331 32355 357
rect 32262 315 32355 331
rect 32217 255 32287 277
rect 32217 221 32229 255
rect 32263 221 32287 255
rect 32217 203 32287 221
rect 32217 169 32240 203
rect 32274 169 32287 203
rect 32217 153 32287 169
rect 32321 197 32355 315
rect 32389 271 32423 427
rect 32457 459 32491 475
rect 32538 441 32554 475
rect 32588 441 32604 475
rect 32638 459 32672 475
rect 32457 407 32491 425
rect 32731 451 32751 485
rect 32785 451 32805 485
rect 32731 435 32805 451
rect 32839 477 32873 493
rect 32638 407 32672 425
rect 32457 373 32672 407
rect 32839 401 32873 443
rect 32920 484 33094 493
rect 32920 450 32936 484
rect 32970 450 33094 484
rect 32920 425 33094 450
rect 33128 485 33178 527
rect 33162 451 33178 485
rect 33282 485 33426 527
rect 33128 435 33178 451
rect 33212 459 33246 475
rect 32761 367 32873 401
rect 32761 339 32795 367
rect 32495 305 32511 339
rect 32545 305 32795 339
rect 32934 357 32945 391
rect 32979 365 33026 391
rect 32934 333 32976 357
rect 32389 251 32727 271
rect 32389 237 32693 251
rect 32321 163 32342 197
rect 32376 163 32392 197
rect 32321 153 32392 163
rect 32426 95 32460 237
rect 32501 187 32597 203
rect 32535 153 32573 187
rect 32631 169 32659 203
rect 32693 201 32727 217
rect 32607 153 32659 169
rect 32761 167 32795 305
rect 31943 69 31977 85
rect 31843 17 31909 59
rect 32049 55 32065 89
rect 32099 55 32115 89
rect 32149 61 32198 95
rect 32232 61 32248 95
rect 32289 61 32305 95
rect 32339 61 32460 95
rect 32635 93 32701 109
rect 32049 17 32115 55
rect 32635 59 32651 93
rect 32685 59 32701 93
rect 32635 17 32701 59
rect 32743 89 32795 167
rect 32833 331 32976 333
rect 33010 331 33026 365
rect 33060 349 33094 425
rect 33282 451 33298 485
rect 33332 451 33376 485
rect 33410 451 33426 485
rect 33460 477 33541 493
rect 33692 485 33726 527
rect 33212 417 33246 425
rect 33494 443 33541 477
rect 33212 383 33372 417
rect 32833 299 32968 331
rect 33060 315 33254 349
rect 33288 315 33304 349
rect 32833 191 32875 299
rect 33060 297 33094 315
rect 32833 157 32841 191
rect 32833 141 32875 157
rect 32909 255 32979 265
rect 32909 239 32945 255
rect 32909 205 32937 239
rect 32971 205 32979 221
rect 32909 141 32979 205
rect 33013 263 33094 297
rect 33013 107 33047 263
rect 33161 250 33269 281
rect 33338 265 33372 383
rect 33460 409 33541 443
rect 33494 375 33541 409
rect 33460 341 33541 375
rect 33494 307 33541 341
rect 33460 291 33541 307
rect 33338 259 33427 265
rect 33195 241 33269 250
rect 33081 213 33125 229
rect 33115 179 33125 213
rect 33161 207 33177 216
rect 33211 207 33269 241
rect 33081 173 33125 179
rect 33221 187 33269 207
rect 33081 139 33187 173
rect 32857 93 33047 107
rect 32743 55 32763 89
rect 32797 55 32813 89
rect 32857 59 32873 93
rect 32907 59 33047 93
rect 32857 51 33047 59
rect 33081 89 33119 105
rect 33081 55 33085 89
rect 33153 93 33187 139
rect 33255 153 33269 187
rect 33221 127 33269 153
rect 33303 249 33427 259
rect 33303 215 33377 249
rect 33411 215 33427 249
rect 33303 199 33427 215
rect 33303 164 33368 199
rect 33475 165 33541 291
rect 33303 109 33367 164
rect 33153 75 33303 93
rect 33337 75 33367 109
rect 33153 59 33367 75
rect 33407 132 33441 154
rect 33081 17 33119 55
rect 33407 17 33441 98
rect 33475 131 33491 165
rect 33525 131 33541 165
rect 33475 97 33541 131
rect 33475 63 33491 97
rect 33525 63 33541 97
rect 33579 451 33595 485
rect 33629 451 33645 485
rect 33579 417 33645 451
rect 33579 383 33595 417
rect 33629 383 33645 417
rect 33579 265 33645 383
rect 33874 477 33925 493
rect 33692 417 33726 451
rect 33692 349 33726 383
rect 33692 299 33726 315
rect 33776 449 33827 465
rect 33810 415 33827 449
rect 33776 381 33827 415
rect 33810 347 33827 381
rect 33874 443 33891 477
rect 33874 409 33925 443
rect 33959 461 34025 527
rect 33959 427 33975 461
rect 34009 427 34025 461
rect 34059 477 34093 493
rect 33874 375 33891 409
rect 34059 409 34093 443
rect 33925 375 34024 393
rect 33874 359 34024 375
rect 33776 325 33827 347
rect 33776 289 33944 325
rect 33785 274 33944 289
rect 33579 249 33751 265
rect 33579 215 33717 249
rect 33579 199 33751 215
rect 33785 240 33816 274
rect 33854 249 33944 274
rect 33854 240 33888 249
rect 33785 215 33888 240
rect 33922 215 33944 249
rect 33579 119 33629 199
rect 33785 195 33944 215
rect 33978 264 34024 359
rect 33978 255 33990 264
rect 34012 221 34024 230
rect 33785 159 33827 195
rect 33978 161 34024 221
rect 33776 143 33827 159
rect 33579 85 33595 119
rect 33579 69 33629 85
rect 33692 113 33726 136
rect 33475 55 33541 63
rect 33692 17 33726 79
rect 33810 109 33827 143
rect 33776 53 33827 109
rect 33874 127 34024 161
rect 33874 119 33925 127
rect 33874 85 33891 119
rect 34059 119 34093 357
rect 34127 333 34192 490
rect 34226 485 34276 527
rect 34226 451 34242 485
rect 34226 435 34276 451
rect 34310 477 34360 493
rect 34310 443 34326 477
rect 34310 427 34360 443
rect 34403 483 34539 493
rect 34403 449 34419 483
rect 34453 449 34539 483
rect 34654 475 34720 527
rect 34847 485 34921 527
rect 34403 427 34539 449
rect 34310 401 34344 427
rect 34265 367 34344 401
rect 34378 391 34471 393
rect 34139 310 34231 333
rect 34139 276 34197 310
rect 34139 175 34231 276
rect 34139 141 34163 175
rect 34201 141 34231 175
rect 34139 123 34231 141
rect 33874 69 33925 85
rect 33959 59 33975 93
rect 34009 59 34025 93
rect 34265 95 34299 367
rect 34378 365 34437 391
rect 34412 357 34437 365
rect 34412 331 34471 357
rect 34378 315 34471 331
rect 34333 255 34403 277
rect 34333 221 34345 255
rect 34379 221 34403 255
rect 34333 203 34403 221
rect 34333 169 34356 203
rect 34390 169 34403 203
rect 34333 153 34403 169
rect 34437 197 34471 315
rect 34505 271 34539 427
rect 34573 459 34607 475
rect 34654 441 34670 475
rect 34704 441 34720 475
rect 34754 459 34788 475
rect 34573 407 34607 425
rect 34847 451 34867 485
rect 34901 451 34921 485
rect 34847 435 34921 451
rect 34955 477 34989 493
rect 34754 407 34788 425
rect 34573 373 34788 407
rect 34955 401 34989 443
rect 35036 484 35210 493
rect 35036 450 35052 484
rect 35086 450 35210 484
rect 35036 425 35210 450
rect 35244 485 35294 527
rect 35278 451 35294 485
rect 35398 485 35542 527
rect 35244 435 35294 451
rect 35328 459 35362 475
rect 34877 367 34989 401
rect 34877 339 34911 367
rect 34611 305 34627 339
rect 34661 305 34911 339
rect 35050 357 35061 391
rect 35095 365 35142 391
rect 35050 333 35092 357
rect 34505 251 34843 271
rect 34505 237 34809 251
rect 34437 163 34458 197
rect 34492 163 34508 197
rect 34437 153 34508 163
rect 34542 95 34576 237
rect 34617 187 34713 203
rect 34651 153 34689 187
rect 34747 169 34775 203
rect 34809 201 34843 217
rect 34723 153 34775 169
rect 34877 167 34911 305
rect 34059 69 34093 85
rect 33959 17 34025 59
rect 34165 55 34181 89
rect 34215 55 34231 89
rect 34265 61 34314 95
rect 34348 61 34364 95
rect 34405 61 34421 95
rect 34455 61 34576 95
rect 34751 93 34817 109
rect 34165 17 34231 55
rect 34751 59 34767 93
rect 34801 59 34817 93
rect 34751 17 34817 59
rect 34859 89 34911 167
rect 34949 331 35092 333
rect 35126 331 35142 365
rect 35176 349 35210 425
rect 35398 451 35414 485
rect 35448 451 35492 485
rect 35526 451 35542 485
rect 35576 477 35657 493
rect 35808 485 35842 527
rect 35328 417 35362 425
rect 35610 443 35657 477
rect 35328 383 35488 417
rect 34949 299 35084 331
rect 35176 315 35370 349
rect 35404 315 35420 349
rect 34949 191 34991 299
rect 35176 297 35210 315
rect 34949 157 34957 191
rect 34949 141 34991 157
rect 35025 255 35095 265
rect 35025 239 35061 255
rect 35025 205 35053 239
rect 35087 205 35095 221
rect 35025 141 35095 205
rect 35129 263 35210 297
rect 35129 107 35163 263
rect 35277 250 35385 281
rect 35454 265 35488 383
rect 35576 409 35657 443
rect 35610 375 35657 409
rect 35576 341 35657 375
rect 35610 307 35657 341
rect 35576 291 35657 307
rect 35454 259 35543 265
rect 35311 241 35385 250
rect 35197 213 35241 229
rect 35231 179 35241 213
rect 35277 207 35293 216
rect 35327 207 35385 241
rect 35197 173 35241 179
rect 35337 187 35385 207
rect 35197 139 35303 173
rect 34973 93 35163 107
rect 34859 55 34879 89
rect 34913 55 34929 89
rect 34973 59 34989 93
rect 35023 59 35163 93
rect 34973 51 35163 59
rect 35197 89 35235 105
rect 35197 55 35201 89
rect 35269 93 35303 139
rect 35371 153 35385 187
rect 35337 127 35385 153
rect 35419 249 35543 259
rect 35419 215 35493 249
rect 35527 215 35543 249
rect 35419 199 35543 215
rect 35419 164 35484 199
rect 35591 165 35657 291
rect 35419 109 35483 164
rect 35269 75 35419 93
rect 35453 75 35483 109
rect 35269 59 35483 75
rect 35523 132 35557 154
rect 35197 17 35235 55
rect 35523 17 35557 98
rect 35591 131 35607 165
rect 35641 131 35657 165
rect 35591 97 35657 131
rect 35591 63 35607 97
rect 35641 63 35657 97
rect 35695 451 35711 485
rect 35745 451 35761 485
rect 35695 417 35761 451
rect 35695 383 35711 417
rect 35745 383 35761 417
rect 35695 265 35761 383
rect 35990 477 36041 493
rect 35808 417 35842 451
rect 35808 349 35842 383
rect 35808 299 35842 315
rect 35892 449 35943 465
rect 35926 415 35943 449
rect 35892 381 35943 415
rect 35926 347 35943 381
rect 35990 443 36007 477
rect 35990 409 36041 443
rect 36075 461 36141 527
rect 36075 427 36091 461
rect 36125 427 36141 461
rect 36175 477 36209 493
rect 35990 375 36007 409
rect 36175 409 36209 443
rect 36041 375 36140 393
rect 35990 359 36140 375
rect 35892 325 35943 347
rect 35892 289 36060 325
rect 35901 274 36060 289
rect 35695 249 35867 265
rect 35695 215 35833 249
rect 35695 199 35867 215
rect 35901 240 35932 274
rect 35970 249 36060 274
rect 35970 240 36004 249
rect 35901 215 36004 240
rect 36038 215 36060 249
rect 35695 119 35745 199
rect 35901 195 36060 215
rect 36094 264 36140 359
rect 36094 255 36106 264
rect 36128 221 36140 230
rect 35901 159 35943 195
rect 36094 161 36140 221
rect 35892 143 35943 159
rect 35695 85 35711 119
rect 35695 69 35745 85
rect 35808 113 35842 136
rect 35591 55 35657 63
rect 35808 17 35842 79
rect 35926 109 35943 143
rect 35892 53 35943 109
rect 35990 127 36140 161
rect 35990 119 36041 127
rect 35990 85 36007 119
rect 36175 119 36209 357
rect 36243 333 36308 490
rect 36342 485 36392 527
rect 36342 451 36358 485
rect 36342 435 36392 451
rect 36426 477 36476 493
rect 36426 443 36442 477
rect 36426 427 36476 443
rect 36519 483 36655 493
rect 36519 449 36535 483
rect 36569 449 36655 483
rect 36770 475 36836 527
rect 36963 485 37037 527
rect 36519 427 36655 449
rect 36426 401 36460 427
rect 36381 367 36460 401
rect 36494 391 36587 393
rect 36255 310 36347 333
rect 36255 276 36313 310
rect 36255 175 36347 276
rect 36255 141 36279 175
rect 36317 141 36347 175
rect 36255 123 36347 141
rect 35990 69 36041 85
rect 36075 59 36091 93
rect 36125 59 36141 93
rect 36381 95 36415 367
rect 36494 365 36553 391
rect 36528 357 36553 365
rect 36528 331 36587 357
rect 36494 315 36587 331
rect 36449 255 36519 277
rect 36449 221 36461 255
rect 36495 221 36519 255
rect 36449 203 36519 221
rect 36449 169 36472 203
rect 36506 169 36519 203
rect 36449 153 36519 169
rect 36553 197 36587 315
rect 36621 271 36655 427
rect 36689 459 36723 475
rect 36770 441 36786 475
rect 36820 441 36836 475
rect 36870 459 36904 475
rect 36689 407 36723 425
rect 36963 451 36983 485
rect 37017 451 37037 485
rect 36963 435 37037 451
rect 37071 477 37105 493
rect 36870 407 36904 425
rect 36689 373 36904 407
rect 37071 401 37105 443
rect 37152 484 37326 493
rect 37152 450 37168 484
rect 37202 450 37326 484
rect 37152 425 37326 450
rect 37360 485 37410 527
rect 37394 451 37410 485
rect 37514 485 37658 527
rect 37360 435 37410 451
rect 37444 459 37478 475
rect 36993 367 37105 401
rect 36993 339 37027 367
rect 36727 305 36743 339
rect 36777 305 37027 339
rect 37166 357 37177 391
rect 37211 365 37258 391
rect 37166 333 37208 357
rect 36621 251 36959 271
rect 36621 237 36925 251
rect 36553 163 36574 197
rect 36608 163 36624 197
rect 36553 153 36624 163
rect 36658 95 36692 237
rect 36733 187 36829 203
rect 36767 153 36805 187
rect 36863 169 36891 203
rect 36925 201 36959 217
rect 36839 153 36891 169
rect 36993 167 37027 305
rect 36175 69 36209 85
rect 36075 17 36141 59
rect 36281 55 36297 89
rect 36331 55 36347 89
rect 36381 61 36430 95
rect 36464 61 36480 95
rect 36521 61 36537 95
rect 36571 61 36692 95
rect 36867 93 36933 109
rect 36281 17 36347 55
rect 36867 59 36883 93
rect 36917 59 36933 93
rect 36867 17 36933 59
rect 36975 89 37027 167
rect 37065 331 37208 333
rect 37242 331 37258 365
rect 37292 349 37326 425
rect 37514 451 37530 485
rect 37564 451 37608 485
rect 37642 451 37658 485
rect 37692 477 37773 493
rect 37924 485 37958 527
rect 37444 417 37478 425
rect 37726 443 37773 477
rect 37444 383 37604 417
rect 37065 299 37200 331
rect 37292 315 37486 349
rect 37520 315 37536 349
rect 37065 191 37107 299
rect 37292 297 37326 315
rect 37065 157 37073 191
rect 37065 141 37107 157
rect 37141 255 37211 265
rect 37141 239 37177 255
rect 37141 205 37169 239
rect 37203 205 37211 221
rect 37141 141 37211 205
rect 37245 263 37326 297
rect 37245 107 37279 263
rect 37393 250 37501 281
rect 37570 265 37604 383
rect 37692 409 37773 443
rect 37726 375 37773 409
rect 37692 341 37773 375
rect 37726 307 37773 341
rect 37692 291 37773 307
rect 37570 259 37659 265
rect 37427 241 37501 250
rect 37313 213 37357 229
rect 37347 179 37357 213
rect 37393 207 37409 216
rect 37443 207 37501 241
rect 37313 173 37357 179
rect 37453 187 37501 207
rect 37313 139 37419 173
rect 37089 93 37279 107
rect 36975 55 36995 89
rect 37029 55 37045 89
rect 37089 59 37105 93
rect 37139 59 37279 93
rect 37089 51 37279 59
rect 37313 89 37351 105
rect 37313 55 37317 89
rect 37385 93 37419 139
rect 37487 153 37501 187
rect 37453 127 37501 153
rect 37535 249 37659 259
rect 37535 215 37609 249
rect 37643 215 37659 249
rect 37535 199 37659 215
rect 37535 164 37600 199
rect 37707 165 37773 291
rect 37535 109 37599 164
rect 37385 75 37535 93
rect 37569 75 37599 109
rect 37385 59 37599 75
rect 37639 132 37673 154
rect 37313 17 37351 55
rect 37639 17 37673 98
rect 37707 131 37723 165
rect 37757 131 37773 165
rect 37707 97 37773 131
rect 37707 63 37723 97
rect 37757 63 37773 97
rect 37811 451 37827 485
rect 37861 451 37877 485
rect 37811 417 37877 451
rect 37811 383 37827 417
rect 37861 383 37877 417
rect 37811 265 37877 383
rect 38106 477 38157 493
rect 37924 417 37958 451
rect 37924 349 37958 383
rect 37924 299 37958 315
rect 38008 449 38059 465
rect 38042 415 38059 449
rect 38008 381 38059 415
rect 38042 347 38059 381
rect 38106 443 38123 477
rect 38106 409 38157 443
rect 38191 461 38257 527
rect 38191 427 38207 461
rect 38241 427 38257 461
rect 38291 477 38325 493
rect 38106 375 38123 409
rect 38291 409 38325 443
rect 38157 375 38256 393
rect 38106 359 38256 375
rect 38008 325 38059 347
rect 38008 289 38176 325
rect 38017 274 38176 289
rect 37811 249 37983 265
rect 37811 215 37949 249
rect 37811 199 37983 215
rect 38017 240 38048 274
rect 38086 249 38176 274
rect 38086 240 38120 249
rect 38017 215 38120 240
rect 38154 215 38176 249
rect 37811 119 37861 199
rect 38017 195 38176 215
rect 38210 264 38256 359
rect 38210 255 38222 264
rect 38244 221 38256 230
rect 38017 159 38059 195
rect 38210 161 38256 221
rect 38008 143 38059 159
rect 37811 85 37827 119
rect 37811 69 37861 85
rect 37924 113 37958 136
rect 37707 55 37773 63
rect 37924 17 37958 79
rect 38042 109 38059 143
rect 38008 53 38059 109
rect 38106 127 38256 161
rect 38106 119 38157 127
rect 38106 85 38123 119
rect 38291 119 38325 357
rect 38359 333 38424 490
rect 38458 485 38508 527
rect 38458 451 38474 485
rect 38458 435 38508 451
rect 38542 477 38592 493
rect 38542 443 38558 477
rect 38542 427 38592 443
rect 38635 483 38771 493
rect 38635 449 38651 483
rect 38685 449 38771 483
rect 38886 475 38952 527
rect 39079 485 39153 527
rect 38635 427 38771 449
rect 38542 401 38576 427
rect 38497 367 38576 401
rect 38610 391 38703 393
rect 38371 310 38463 333
rect 38371 276 38429 310
rect 38371 175 38463 276
rect 38371 141 38395 175
rect 38433 141 38463 175
rect 38371 123 38463 141
rect 38106 69 38157 85
rect 38191 59 38207 93
rect 38241 59 38257 93
rect 38497 95 38531 367
rect 38610 365 38669 391
rect 38644 357 38669 365
rect 38644 331 38703 357
rect 38610 315 38703 331
rect 38565 255 38635 277
rect 38565 221 38577 255
rect 38611 221 38635 255
rect 38565 203 38635 221
rect 38565 169 38588 203
rect 38622 169 38635 203
rect 38565 153 38635 169
rect 38669 197 38703 315
rect 38737 271 38771 427
rect 38805 459 38839 475
rect 38886 441 38902 475
rect 38936 441 38952 475
rect 38986 459 39020 475
rect 38805 407 38839 425
rect 39079 451 39099 485
rect 39133 451 39153 485
rect 39079 435 39153 451
rect 39187 477 39221 493
rect 38986 407 39020 425
rect 38805 373 39020 407
rect 39187 401 39221 443
rect 39268 484 39442 493
rect 39268 450 39284 484
rect 39318 450 39442 484
rect 39268 425 39442 450
rect 39476 485 39526 527
rect 39510 451 39526 485
rect 39630 485 39774 527
rect 39476 435 39526 451
rect 39560 459 39594 475
rect 39109 367 39221 401
rect 39109 339 39143 367
rect 38843 305 38859 339
rect 38893 305 39143 339
rect 39282 357 39293 391
rect 39327 365 39374 391
rect 39282 333 39324 357
rect 38737 251 39075 271
rect 38737 237 39041 251
rect 38669 163 38690 197
rect 38724 163 38740 197
rect 38669 153 38740 163
rect 38774 95 38808 237
rect 38849 187 38945 203
rect 38883 153 38921 187
rect 38979 169 39007 203
rect 39041 201 39075 217
rect 38955 153 39007 169
rect 39109 167 39143 305
rect 38291 69 38325 85
rect 38191 17 38257 59
rect 38397 55 38413 89
rect 38447 55 38463 89
rect 38497 61 38546 95
rect 38580 61 38596 95
rect 38637 61 38653 95
rect 38687 61 38808 95
rect 38983 93 39049 109
rect 38397 17 38463 55
rect 38983 59 38999 93
rect 39033 59 39049 93
rect 38983 17 39049 59
rect 39091 89 39143 167
rect 39181 331 39324 333
rect 39358 331 39374 365
rect 39408 349 39442 425
rect 39630 451 39646 485
rect 39680 451 39724 485
rect 39758 451 39774 485
rect 39808 477 39889 493
rect 40040 485 40074 527
rect 39560 417 39594 425
rect 39842 443 39889 477
rect 39560 383 39720 417
rect 39181 299 39316 331
rect 39408 315 39602 349
rect 39636 315 39652 349
rect 39181 191 39223 299
rect 39408 297 39442 315
rect 39181 157 39189 191
rect 39181 141 39223 157
rect 39257 255 39327 265
rect 39257 239 39293 255
rect 39257 205 39285 239
rect 39319 205 39327 221
rect 39257 141 39327 205
rect 39361 263 39442 297
rect 39361 107 39395 263
rect 39509 250 39617 281
rect 39686 265 39720 383
rect 39808 409 39889 443
rect 39842 375 39889 409
rect 39808 341 39889 375
rect 39842 307 39889 341
rect 39808 291 39889 307
rect 39686 259 39775 265
rect 39543 241 39617 250
rect 39429 213 39473 229
rect 39463 179 39473 213
rect 39509 207 39525 216
rect 39559 207 39617 241
rect 39429 173 39473 179
rect 39569 187 39617 207
rect 39429 139 39535 173
rect 39205 93 39395 107
rect 39091 55 39111 89
rect 39145 55 39161 89
rect 39205 59 39221 93
rect 39255 59 39395 93
rect 39205 51 39395 59
rect 39429 89 39467 105
rect 39429 55 39433 89
rect 39501 93 39535 139
rect 39603 153 39617 187
rect 39569 127 39617 153
rect 39651 249 39775 259
rect 39651 215 39725 249
rect 39759 215 39775 249
rect 39651 199 39775 215
rect 39651 164 39716 199
rect 39823 165 39889 291
rect 39651 109 39715 164
rect 39501 75 39651 93
rect 39685 75 39715 109
rect 39501 59 39715 75
rect 39755 132 39789 154
rect 39429 17 39467 55
rect 39755 17 39789 98
rect 39823 131 39839 165
rect 39873 131 39889 165
rect 39823 97 39889 131
rect 39823 63 39839 97
rect 39873 63 39889 97
rect 39927 451 39943 485
rect 39977 451 39993 485
rect 39927 417 39993 451
rect 39927 383 39943 417
rect 39977 383 39993 417
rect 39927 265 39993 383
rect 40222 477 40273 493
rect 40040 417 40074 451
rect 40040 349 40074 383
rect 40040 299 40074 315
rect 40124 449 40175 465
rect 40158 415 40175 449
rect 40124 381 40175 415
rect 40158 347 40175 381
rect 40222 443 40239 477
rect 40222 409 40273 443
rect 40307 461 40373 527
rect 40307 427 40323 461
rect 40357 427 40373 461
rect 40407 477 40441 493
rect 40222 375 40239 409
rect 40407 409 40441 443
rect 40273 375 40372 393
rect 40222 359 40372 375
rect 40124 325 40175 347
rect 40124 289 40292 325
rect 40133 274 40292 289
rect 39927 249 40099 265
rect 39927 215 40065 249
rect 39927 199 40099 215
rect 40133 240 40164 274
rect 40202 249 40292 274
rect 40202 240 40236 249
rect 40133 215 40236 240
rect 40270 215 40292 249
rect 39927 119 39977 199
rect 40133 195 40292 215
rect 40326 264 40372 359
rect 40326 255 40338 264
rect 40360 221 40372 230
rect 40133 159 40175 195
rect 40326 161 40372 221
rect 40124 143 40175 159
rect 39927 85 39943 119
rect 39927 69 39977 85
rect 40040 113 40074 136
rect 39823 55 39889 63
rect 40040 17 40074 79
rect 40158 109 40175 143
rect 40124 53 40175 109
rect 40222 127 40372 161
rect 40222 119 40273 127
rect 40222 85 40239 119
rect 40407 119 40441 357
rect 40475 333 40540 490
rect 40574 485 40624 527
rect 40574 451 40590 485
rect 40574 435 40624 451
rect 40658 477 40708 493
rect 40658 443 40674 477
rect 40658 427 40708 443
rect 40751 483 40887 493
rect 40751 449 40767 483
rect 40801 449 40887 483
rect 41002 475 41068 527
rect 41195 485 41269 527
rect 40751 427 40887 449
rect 40658 401 40692 427
rect 40613 367 40692 401
rect 40726 391 40819 393
rect 40487 310 40579 333
rect 40487 276 40545 310
rect 40487 175 40579 276
rect 40487 141 40511 175
rect 40549 141 40579 175
rect 40487 123 40579 141
rect 40222 69 40273 85
rect 40307 59 40323 93
rect 40357 59 40373 93
rect 40613 95 40647 367
rect 40726 365 40785 391
rect 40760 357 40785 365
rect 40760 331 40819 357
rect 40726 315 40819 331
rect 40681 255 40751 277
rect 40681 221 40693 255
rect 40727 221 40751 255
rect 40681 203 40751 221
rect 40681 169 40704 203
rect 40738 169 40751 203
rect 40681 153 40751 169
rect 40785 197 40819 315
rect 40853 271 40887 427
rect 40921 459 40955 475
rect 41002 441 41018 475
rect 41052 441 41068 475
rect 41102 459 41136 475
rect 40921 407 40955 425
rect 41195 451 41215 485
rect 41249 451 41269 485
rect 41195 435 41269 451
rect 41303 477 41337 493
rect 41102 407 41136 425
rect 40921 373 41136 407
rect 41303 401 41337 443
rect 41384 484 41558 493
rect 41384 450 41400 484
rect 41434 450 41558 484
rect 41384 425 41558 450
rect 41592 485 41642 527
rect 41626 451 41642 485
rect 41746 485 41890 527
rect 41592 435 41642 451
rect 41676 459 41710 475
rect 41225 367 41337 401
rect 41225 339 41259 367
rect 40959 305 40975 339
rect 41009 305 41259 339
rect 41398 357 41409 391
rect 41443 365 41490 391
rect 41398 333 41440 357
rect 40853 251 41191 271
rect 40853 237 41157 251
rect 40785 163 40806 197
rect 40840 163 40856 197
rect 40785 153 40856 163
rect 40890 95 40924 237
rect 40965 187 41061 203
rect 40999 153 41037 187
rect 41095 169 41123 203
rect 41157 201 41191 217
rect 41071 153 41123 169
rect 41225 167 41259 305
rect 40407 69 40441 85
rect 40307 17 40373 59
rect 40513 55 40529 89
rect 40563 55 40579 89
rect 40613 61 40662 95
rect 40696 61 40712 95
rect 40753 61 40769 95
rect 40803 61 40924 95
rect 41099 93 41165 109
rect 40513 17 40579 55
rect 41099 59 41115 93
rect 41149 59 41165 93
rect 41099 17 41165 59
rect 41207 89 41259 167
rect 41297 331 41440 333
rect 41474 331 41490 365
rect 41524 349 41558 425
rect 41746 451 41762 485
rect 41796 451 41840 485
rect 41874 451 41890 485
rect 41924 477 42005 493
rect 42156 485 42190 527
rect 41676 417 41710 425
rect 41958 443 42005 477
rect 41676 383 41836 417
rect 41297 299 41432 331
rect 41524 315 41718 349
rect 41752 315 41768 349
rect 41297 191 41339 299
rect 41524 297 41558 315
rect 41297 157 41305 191
rect 41297 141 41339 157
rect 41373 255 41443 265
rect 41373 239 41409 255
rect 41373 205 41401 239
rect 41435 205 41443 221
rect 41373 141 41443 205
rect 41477 263 41558 297
rect 41477 107 41511 263
rect 41625 250 41733 281
rect 41802 265 41836 383
rect 41924 409 42005 443
rect 41958 375 42005 409
rect 41924 341 42005 375
rect 41958 307 42005 341
rect 41924 291 42005 307
rect 41802 259 41891 265
rect 41659 241 41733 250
rect 41545 213 41589 229
rect 41579 179 41589 213
rect 41625 207 41641 216
rect 41675 207 41733 241
rect 41545 173 41589 179
rect 41685 187 41733 207
rect 41545 139 41651 173
rect 41321 93 41511 107
rect 41207 55 41227 89
rect 41261 55 41277 89
rect 41321 59 41337 93
rect 41371 59 41511 93
rect 41321 51 41511 59
rect 41545 89 41583 105
rect 41545 55 41549 89
rect 41617 93 41651 139
rect 41719 153 41733 187
rect 41685 127 41733 153
rect 41767 249 41891 259
rect 41767 215 41841 249
rect 41875 215 41891 249
rect 41767 199 41891 215
rect 41767 164 41832 199
rect 41939 165 42005 291
rect 41767 109 41831 164
rect 41617 75 41767 93
rect 41801 75 41831 109
rect 41617 59 41831 75
rect 41871 132 41905 154
rect 41545 17 41583 55
rect 41871 17 41905 98
rect 41939 131 41955 165
rect 41989 131 42005 165
rect 41939 97 42005 131
rect 41939 63 41955 97
rect 41989 63 42005 97
rect 42043 451 42059 485
rect 42093 451 42109 485
rect 42043 417 42109 451
rect 42043 383 42059 417
rect 42093 383 42109 417
rect 42043 265 42109 383
rect 42156 417 42190 451
rect 42156 349 42190 383
rect 42156 299 42190 315
rect 42240 449 42291 465
rect 42274 415 42291 449
rect 42240 381 42291 415
rect 42274 347 42291 381
rect 42240 325 42291 347
rect 42240 289 42320 325
rect 42249 274 42320 289
rect 42043 249 42215 265
rect 42043 215 42181 249
rect 42043 199 42215 215
rect 42249 240 42280 274
rect 42318 240 42320 274
rect 42043 119 42093 199
rect 42249 195 42320 240
rect 42249 159 42291 195
rect 42240 143 42291 159
rect 42043 85 42059 119
rect 42043 69 42093 85
rect 42156 113 42190 136
rect 41939 55 42005 63
rect 42156 17 42190 79
rect 42274 109 42291 143
rect 42240 53 42291 109
rect 0 -41 29 17
rect 63 -41 121 17
rect 155 -41 213 17
rect 247 -41 305 17
rect 339 -41 397 17
rect 431 -41 489 17
rect 523 -41 581 17
rect 615 -41 673 17
rect 707 -41 765 17
rect 799 -41 857 17
rect 891 -41 949 17
rect 983 -41 1041 17
rect 1075 -41 1133 17
rect 1167 -41 1225 17
rect 1259 -41 1317 17
rect 1351 -41 1409 17
rect 1443 -41 1501 17
rect 1535 -41 1593 17
rect 1627 -41 1685 17
rect 1719 -41 1777 17
rect 1811 -41 1869 17
rect 1903 -41 1961 17
rect 1995 -41 2053 17
rect 2087 -41 2145 17
rect 2179 -41 2237 17
rect 2271 -41 2329 17
rect 2363 -41 2421 17
rect 2455 -41 2513 17
rect 2547 -41 2605 17
rect 2639 -41 2697 17
rect 2731 -41 2789 17
rect 2823 -41 2881 17
rect 2915 -41 2973 17
rect 3007 -41 3065 17
rect 3099 -41 3157 17
rect 3191 -41 3249 17
rect 3283 -41 3341 17
rect 3375 -41 3433 17
rect 3467 -41 3525 17
rect 3559 -41 3617 17
rect 3651 -41 3709 17
rect 3743 -41 3801 17
rect 3835 -41 3893 17
rect 3927 -41 3985 17
rect 4019 -41 4077 17
rect 4111 -41 4169 17
rect 4203 -41 4261 17
rect 4295 -41 4353 17
rect 4387 -41 4445 17
rect 4479 -41 4537 17
rect 4571 -41 4629 17
rect 4663 -41 4721 17
rect 4755 -41 4813 17
rect 4847 -41 4905 17
rect 4939 -41 4997 17
rect 5031 -41 5089 17
rect 5123 -41 5181 17
rect 5215 -41 5273 17
rect 5307 -41 5365 17
rect 5399 -41 5457 17
rect 5491 -41 5549 17
rect 5583 -41 5641 17
rect 5675 -41 5733 17
rect 5767 -41 5825 17
rect 5859 -41 5917 17
rect 5951 -41 6009 17
rect 6043 -41 6101 17
rect 6135 -41 6193 17
rect 6227 -41 6285 17
rect 6319 -41 6377 17
rect 6411 -41 6469 17
rect 6503 -41 6561 17
rect 6595 -41 6653 17
rect 6687 -41 6745 17
rect 6779 -41 6837 17
rect 6871 -41 6929 17
rect 6963 -41 7021 17
rect 7055 -41 7113 17
rect 7147 -41 7205 17
rect 7239 -41 7297 17
rect 7331 -41 7389 17
rect 7423 -41 7481 17
rect 7515 -41 7573 17
rect 7607 -41 7665 17
rect 7699 -41 7757 17
rect 7791 -41 7849 17
rect 7883 -41 7941 17
rect 7975 -41 8033 17
rect 8067 -41 8125 17
rect 8159 -41 8217 17
rect 8251 -41 8309 17
rect 8343 -41 8401 17
rect 8435 -41 8493 17
rect 8527 -41 8585 17
rect 8619 -41 8677 17
rect 8711 -41 8769 17
rect 8803 -41 8861 17
rect 8895 -41 8953 17
rect 8987 -41 9045 17
rect 9079 -41 9137 17
rect 9171 -41 9229 17
rect 9263 -41 9321 17
rect 9355 -41 9413 17
rect 9447 -41 9505 17
rect 9539 -41 9597 17
rect 9631 -41 9689 17
rect 9723 -41 9781 17
rect 9815 -41 9873 17
rect 9907 -41 9965 17
rect 9999 -41 10057 17
rect 10091 -41 10149 17
rect 10183 -41 10241 17
rect 10275 -41 10333 17
rect 10367 -41 10425 17
rect 10459 -41 10517 17
rect 10551 -41 10609 17
rect 10643 -41 10701 17
rect 10735 -41 10793 17
rect 10827 -41 10885 17
rect 10919 -41 10977 17
rect 11011 -41 11069 17
rect 11103 -41 11161 17
rect 11195 -41 11253 17
rect 11287 -41 11345 17
rect 11379 -41 11437 17
rect 11471 -41 11529 17
rect 11563 -41 11621 17
rect 11655 -41 11713 17
rect 11747 -41 11805 17
rect 11839 -41 11897 17
rect 11931 -41 11989 17
rect 12023 -41 12081 17
rect 12115 -41 12173 17
rect 12207 -41 12265 17
rect 12299 -41 12357 17
rect 12391 -41 12449 17
rect 12483 -41 12541 17
rect 12575 -41 12633 17
rect 12667 -41 12725 17
rect 12759 -41 12817 17
rect 12851 -41 12909 17
rect 12943 -41 13001 17
rect 13035 -41 13093 17
rect 13127 -41 13185 17
rect 13219 -41 13277 17
rect 13311 -41 13369 17
rect 13403 -41 13461 17
rect 13495 -41 13553 17
rect 13587 -41 13645 17
rect 13679 -41 13737 17
rect 13771 -41 13829 17
rect 13863 -41 13921 17
rect 13955 -41 14013 17
rect 14047 -41 14105 17
rect 14139 -41 14197 17
rect 14231 -41 14289 17
rect 14323 -41 14381 17
rect 14415 -41 14473 17
rect 14507 -41 14565 17
rect 14599 -41 14657 17
rect 14691 -41 14749 17
rect 14783 -41 14841 17
rect 14875 -41 14933 17
rect 14967 -41 15025 17
rect 15059 -41 15117 17
rect 15151 -41 15209 17
rect 15243 -41 15301 17
rect 15335 -41 15393 17
rect 15427 -41 15485 17
rect 15519 -41 15577 17
rect 15611 -41 15669 17
rect 15703 -41 15761 17
rect 15795 -41 15853 17
rect 15887 -41 15945 17
rect 15979 -41 16037 17
rect 16071 -41 16129 17
rect 16163 -41 16221 17
rect 16255 -41 16313 17
rect 16347 -41 16405 17
rect 16439 -41 16497 17
rect 16531 -41 16589 17
rect 16623 -41 16681 17
rect 16715 -41 16773 17
rect 16807 -41 16865 17
rect 16899 -41 16957 17
rect 16991 -41 17049 17
rect 17083 -41 17141 17
rect 17175 -41 17233 17
rect 17267 -41 17325 17
rect 17359 -41 17417 17
rect 17451 -41 17509 17
rect 17543 -41 17601 17
rect 17635 -41 17693 17
rect 17727 -41 17785 17
rect 17819 -41 17877 17
rect 17911 -41 17969 17
rect 18003 -41 18061 17
rect 18095 -41 18153 17
rect 18187 -41 18245 17
rect 18279 -41 18337 17
rect 18371 -41 18429 17
rect 18463 -41 18521 17
rect 18555 -41 18613 17
rect 18647 -41 18705 17
rect 18739 -41 18797 17
rect 18831 -41 18889 17
rect 18923 -41 18981 17
rect 19015 -41 19073 17
rect 19107 -41 19165 17
rect 19199 -41 19257 17
rect 19291 -41 19349 17
rect 19383 -41 19441 17
rect 19475 -41 19533 17
rect 19567 -41 19625 17
rect 19659 -41 19717 17
rect 19751 -41 19809 17
rect 19843 -41 19901 17
rect 19935 -41 19993 17
rect 20027 -41 20085 17
rect 20119 -41 20177 17
rect 20211 -41 20269 17
rect 20303 -41 20361 17
rect 20395 -41 20453 17
rect 20487 -41 20545 17
rect 20579 -41 20637 17
rect 20671 -41 20729 17
rect 20763 -41 20821 17
rect 20855 -41 20913 17
rect 20947 -41 21005 17
rect 21039 -41 21097 17
rect 21131 -41 21189 17
rect 21223 -41 21281 17
rect 21315 -41 21373 17
rect 21407 -41 21465 17
rect 21499 -41 21557 17
rect 21591 -41 21649 17
rect 21683 -41 21741 17
rect 21775 -41 21833 17
rect 21867 -41 21925 17
rect 21959 -41 22017 17
rect 22051 -41 22109 17
rect 22143 -41 22201 17
rect 22235 -41 22293 17
rect 22327 -41 22385 17
rect 22419 -41 22477 17
rect 22511 -41 22569 17
rect 22603 -41 22661 17
rect 22695 -41 22753 17
rect 22787 -41 22845 17
rect 22879 -41 22937 17
rect 22971 -41 23029 17
rect 23063 -41 23121 17
rect 23155 -41 23213 17
rect 23247 -41 23305 17
rect 23339 -41 23397 17
rect 23431 -41 23489 17
rect 23523 -41 23581 17
rect 23615 -41 23673 17
rect 23707 -41 23765 17
rect 23799 -41 23857 17
rect 23891 -41 23949 17
rect 23983 -41 24041 17
rect 24075 -41 24133 17
rect 24167 -41 24225 17
rect 24259 -41 24317 17
rect 24351 -41 24409 17
rect 24443 -41 24501 17
rect 24535 -41 24593 17
rect 24627 -41 24685 17
rect 24719 -41 24777 17
rect 24811 -41 24869 17
rect 24903 -41 24961 17
rect 24995 -41 25053 17
rect 25087 -41 25145 17
rect 25179 -41 25237 17
rect 25271 -41 25329 17
rect 25363 -41 25421 17
rect 25455 -41 25513 17
rect 25547 -41 25605 17
rect 25639 -41 25697 17
rect 25731 -41 25789 17
rect 25823 -41 25881 17
rect 25915 -41 25973 17
rect 26007 -41 26065 17
rect 26099 -41 26157 17
rect 26191 -41 26249 17
rect 26283 -41 26341 17
rect 26375 -41 26433 17
rect 26467 -41 26525 17
rect 26559 -41 26617 17
rect 26651 -41 26709 17
rect 26743 -41 26801 17
rect 26835 -41 26893 17
rect 26927 -41 26985 17
rect 27019 -41 27077 17
rect 27111 -41 27169 17
rect 27203 -41 27261 17
rect 27295 -41 27353 17
rect 27387 -41 27445 17
rect 27479 -41 27537 17
rect 27571 -41 27629 17
rect 27663 -41 27721 17
rect 27755 -41 27813 17
rect 27847 -41 27905 17
rect 27939 -41 27997 17
rect 28031 -41 28089 17
rect 28123 -41 28181 17
rect 28215 -41 28273 17
rect 28307 -41 28365 17
rect 28399 -41 28457 17
rect 28491 -41 28549 17
rect 28583 -41 28641 17
rect 28675 -41 28733 17
rect 28767 -41 28825 17
rect 28859 -41 28917 17
rect 28951 -41 29009 17
rect 29043 -41 29101 17
rect 29135 -41 29193 17
rect 29227 -41 29285 17
rect 29319 -41 29377 17
rect 29411 -41 29469 17
rect 29503 -41 29561 17
rect 29595 -41 29653 17
rect 29687 -41 29745 17
rect 29779 -41 29837 17
rect 29871 -41 29929 17
rect 29963 -41 30021 17
rect 30055 -41 30113 17
rect 30147 -41 30205 17
rect 30239 -41 30297 17
rect 30331 -41 30389 17
rect 30423 -41 30481 17
rect 30515 -41 30573 17
rect 30607 -41 30665 17
rect 30699 -41 30757 17
rect 30791 -41 30849 17
rect 30883 -41 30941 17
rect 30975 -41 31033 17
rect 31067 -41 31125 17
rect 31159 -41 31217 17
rect 31251 -41 31309 17
rect 31343 -41 31401 17
rect 31435 -41 31493 17
rect 31527 -41 31585 17
rect 31619 -41 31677 17
rect 31711 -41 31769 17
rect 31803 -41 31861 17
rect 31895 -41 31953 17
rect 31987 -41 32045 17
rect 32079 -41 32137 17
rect 32171 -41 32229 17
rect 32263 -41 32321 17
rect 32355 -41 32413 17
rect 32447 -41 32505 17
rect 32539 -41 32597 17
rect 32631 -41 32689 17
rect 32723 -41 32781 17
rect 32815 -41 32873 17
rect 32907 -41 32965 17
rect 32999 -41 33057 17
rect 33091 -41 33149 17
rect 33183 -41 33241 17
rect 33275 -41 33333 17
rect 33367 -41 33425 17
rect 33459 -41 33517 17
rect 33551 -41 33609 17
rect 33643 -41 33701 17
rect 33735 -41 33793 17
rect 33827 -41 33885 17
rect 33919 -41 33977 17
rect 34011 -41 34069 17
rect 34103 -41 34161 17
rect 34195 -41 34253 17
rect 34287 -41 34345 17
rect 34379 -41 34437 17
rect 34471 -41 34529 17
rect 34563 -41 34621 17
rect 34655 -41 34713 17
rect 34747 -41 34805 17
rect 34839 -41 34897 17
rect 34931 -41 34989 17
rect 35023 -41 35081 17
rect 35115 -41 35173 17
rect 35207 -41 35265 17
rect 35299 -41 35357 17
rect 35391 -41 35449 17
rect 35483 -41 35541 17
rect 35575 -41 35633 17
rect 35667 -41 35725 17
rect 35759 -41 35817 17
rect 35851 -41 35909 17
rect 35943 -41 36001 17
rect 36035 -41 36093 17
rect 36127 -41 36185 17
rect 36219 -41 36277 17
rect 36311 -41 36369 17
rect 36403 -41 36461 17
rect 36495 -41 36553 17
rect 36587 -41 36645 17
rect 36679 -41 36737 17
rect 36771 -41 36829 17
rect 36863 -41 36921 17
rect 36955 -41 37013 17
rect 37047 -41 37105 17
rect 37139 -41 37197 17
rect 37231 -41 37289 17
rect 37323 -41 37381 17
rect 37415 -41 37473 17
rect 37507 -41 37565 17
rect 37599 -41 37657 17
rect 37691 -41 37749 17
rect 37783 -41 37841 17
rect 37875 -41 37933 17
rect 37967 -41 38025 17
rect 38059 -41 38117 17
rect 38151 -41 38209 17
rect 38243 -41 38301 17
rect 38335 -41 38393 17
rect 38427 -41 38485 17
rect 38519 -41 38577 17
rect 38611 -41 38669 17
rect 38703 -41 38761 17
rect 38795 -41 38853 17
rect 38887 -41 38945 17
rect 38979 -41 39037 17
rect 39071 -41 39129 17
rect 39163 -41 39221 17
rect 39255 -41 39313 17
rect 39347 -41 39405 17
rect 39439 -41 39497 17
rect 39531 -41 39589 17
rect 39623 -41 39681 17
rect 39715 -41 39773 17
rect 39807 -41 39865 17
rect 39899 -41 39957 17
rect 39991 -41 40049 17
rect 40083 -41 40141 17
rect 40175 -41 40233 17
rect 40267 -41 40325 17
rect 40359 -41 40417 17
rect 40451 -41 40509 17
rect 40543 -41 40601 17
rect 40635 -41 40693 17
rect 40727 -41 40785 17
rect 40819 -41 40877 17
rect 40911 -41 40969 17
rect 41003 -41 41061 17
rect 41095 -41 41153 17
rect 41187 -41 41245 17
rect 41279 -41 41337 17
rect 41371 -41 41429 17
rect 41463 -41 41521 17
rect 41555 -41 41613 17
rect 41647 -41 41705 17
rect 41739 -41 41797 17
rect 41831 -41 41889 17
rect 41923 -41 41981 17
rect 42015 -41 42073 17
rect 42107 -41 42165 17
rect 42199 -41 42257 17
rect 42291 -41 42320 17
rect 0 -57 42320 -41
<< viali >>
rect 29 551 63 561
rect 29 527 63 551
rect 121 551 155 561
rect 121 527 155 551
rect 213 551 247 561
rect 213 527 247 551
rect 305 551 339 561
rect 305 527 339 551
rect 397 551 431 561
rect 397 527 431 551
rect 489 551 523 561
rect 489 527 523 551
rect 581 551 615 561
rect 581 527 615 551
rect 673 551 707 561
rect 673 527 707 551
rect 765 551 799 561
rect 765 527 799 551
rect 857 551 891 561
rect 857 527 891 551
rect 949 551 983 561
rect 949 527 983 551
rect 1041 551 1075 561
rect 1041 527 1075 551
rect 1133 551 1167 561
rect 1133 527 1167 551
rect 1225 551 1259 561
rect 1225 527 1259 551
rect 1317 551 1351 561
rect 1317 527 1351 551
rect 1409 551 1443 561
rect 1409 527 1443 551
rect 1501 551 1535 561
rect 1501 527 1535 551
rect 1593 551 1627 561
rect 1593 527 1627 551
rect 1685 551 1719 561
rect 1685 527 1719 551
rect 1777 551 1811 561
rect 1777 527 1811 551
rect 1869 551 1903 561
rect 1869 527 1903 551
rect 1961 551 1995 561
rect 1961 527 1995 551
rect 2053 551 2087 561
rect 2053 527 2087 551
rect 2145 551 2179 561
rect 2145 527 2179 551
rect 2237 551 2271 561
rect 2237 527 2271 551
rect 2329 551 2363 561
rect 2329 527 2363 551
rect 2421 551 2455 561
rect 2421 527 2455 551
rect 2513 551 2547 561
rect 2513 527 2547 551
rect 2605 551 2639 561
rect 2605 527 2639 551
rect 2697 551 2731 561
rect 2697 527 2731 551
rect 2789 551 2823 561
rect 2789 527 2823 551
rect 2881 551 2915 561
rect 2881 527 2915 551
rect 2973 551 3007 561
rect 2973 527 3007 551
rect 3065 551 3099 561
rect 3065 527 3099 551
rect 3157 551 3191 561
rect 3157 527 3191 551
rect 3249 551 3283 561
rect 3249 527 3283 551
rect 3341 551 3375 561
rect 3341 527 3375 551
rect 3433 551 3467 561
rect 3433 527 3467 551
rect 3525 551 3559 561
rect 3525 527 3559 551
rect 3617 551 3651 561
rect 3617 527 3651 551
rect 3709 551 3743 561
rect 3709 527 3743 551
rect 3801 551 3835 561
rect 3801 527 3835 551
rect 3893 551 3927 561
rect 3893 527 3927 551
rect 3985 551 4019 561
rect 3985 527 4019 551
rect 4077 551 4111 561
rect 4077 527 4111 551
rect 4169 551 4203 561
rect 4169 527 4203 551
rect 4261 551 4295 561
rect 4261 527 4295 551
rect 4353 551 4387 561
rect 4353 527 4387 551
rect 4445 551 4479 561
rect 4445 527 4479 551
rect 4537 551 4571 561
rect 4537 527 4571 551
rect 4629 551 4663 561
rect 4629 527 4663 551
rect 4721 551 4755 561
rect 4721 527 4755 551
rect 4813 551 4847 561
rect 4813 527 4847 551
rect 4905 551 4939 561
rect 4905 527 4939 551
rect 4997 551 5031 561
rect 4997 527 5031 551
rect 5089 551 5123 561
rect 5089 527 5123 551
rect 5181 551 5215 561
rect 5181 527 5215 551
rect 5273 551 5307 561
rect 5273 527 5307 551
rect 5365 551 5399 561
rect 5365 527 5399 551
rect 5457 551 5491 561
rect 5457 527 5491 551
rect 5549 551 5583 561
rect 5549 527 5583 551
rect 5641 551 5675 561
rect 5641 527 5675 551
rect 5733 551 5767 561
rect 5733 527 5767 551
rect 5825 551 5859 561
rect 5825 527 5859 551
rect 5917 551 5951 561
rect 5917 527 5951 551
rect 6009 551 6043 561
rect 6009 527 6043 551
rect 6101 551 6135 561
rect 6101 527 6135 551
rect 6193 551 6227 561
rect 6193 527 6227 551
rect 6285 551 6319 561
rect 6285 527 6319 551
rect 6377 551 6411 561
rect 6377 527 6411 551
rect 6469 551 6503 561
rect 6469 527 6503 551
rect 6561 551 6595 561
rect 6561 527 6595 551
rect 6653 551 6687 561
rect 6653 527 6687 551
rect 6745 551 6779 561
rect 6745 527 6779 551
rect 6837 551 6871 561
rect 6837 527 6871 551
rect 6929 551 6963 561
rect 6929 527 6963 551
rect 7021 551 7055 561
rect 7021 527 7055 551
rect 7113 551 7147 561
rect 7113 527 7147 551
rect 7205 551 7239 561
rect 7205 527 7239 551
rect 7297 551 7331 561
rect 7297 527 7331 551
rect 7389 551 7423 561
rect 7389 527 7423 551
rect 7481 551 7515 561
rect 7481 527 7515 551
rect 7573 551 7607 561
rect 7573 527 7607 551
rect 7665 551 7699 561
rect 7665 527 7699 551
rect 7757 551 7791 561
rect 7757 527 7791 551
rect 7849 551 7883 561
rect 7849 527 7883 551
rect 7941 551 7975 561
rect 7941 527 7975 551
rect 8033 551 8067 561
rect 8033 527 8067 551
rect 8125 551 8159 561
rect 8125 527 8159 551
rect 8217 551 8251 561
rect 8217 527 8251 551
rect 8309 551 8343 561
rect 8309 527 8343 551
rect 8401 551 8435 561
rect 8401 527 8435 551
rect 8493 551 8527 561
rect 8493 527 8527 551
rect 8585 551 8619 561
rect 8585 527 8619 551
rect 8677 551 8711 561
rect 8677 527 8711 551
rect 8769 551 8803 561
rect 8769 527 8803 551
rect 8861 551 8895 561
rect 8861 527 8895 551
rect 8953 551 8987 561
rect 8953 527 8987 551
rect 9045 551 9079 561
rect 9045 527 9079 551
rect 9137 551 9171 561
rect 9137 527 9171 551
rect 9229 551 9263 561
rect 9229 527 9263 551
rect 9321 551 9355 561
rect 9321 527 9355 551
rect 9413 551 9447 561
rect 9413 527 9447 551
rect 9505 551 9539 561
rect 9505 527 9539 551
rect 9597 551 9631 561
rect 9597 527 9631 551
rect 9689 551 9723 561
rect 9689 527 9723 551
rect 9781 551 9815 561
rect 9781 527 9815 551
rect 9873 551 9907 561
rect 9873 527 9907 551
rect 9965 551 9999 561
rect 9965 527 9999 551
rect 10057 551 10091 561
rect 10057 527 10091 551
rect 10149 551 10183 561
rect 10149 527 10183 551
rect 10241 551 10275 561
rect 10241 527 10275 551
rect 10333 551 10367 561
rect 10333 527 10367 551
rect 10425 551 10459 561
rect 10425 527 10459 551
rect 10517 551 10551 561
rect 10517 527 10551 551
rect 10609 551 10643 561
rect 10609 527 10643 551
rect 10701 551 10735 561
rect 10701 527 10735 551
rect 10793 551 10827 561
rect 10793 527 10827 551
rect 10885 551 10919 561
rect 10885 527 10919 551
rect 10977 551 11011 561
rect 10977 527 11011 551
rect 11069 551 11103 561
rect 11069 527 11103 551
rect 11161 551 11195 561
rect 11161 527 11195 551
rect 11253 551 11287 561
rect 11253 527 11287 551
rect 11345 551 11379 561
rect 11345 527 11379 551
rect 11437 551 11471 561
rect 11437 527 11471 551
rect 11529 551 11563 561
rect 11529 527 11563 551
rect 11621 551 11655 561
rect 11621 527 11655 551
rect 11713 551 11747 561
rect 11713 527 11747 551
rect 11805 551 11839 561
rect 11805 527 11839 551
rect 11897 551 11931 561
rect 11897 527 11931 551
rect 11989 551 12023 561
rect 11989 527 12023 551
rect 12081 551 12115 561
rect 12081 527 12115 551
rect 12173 551 12207 561
rect 12173 527 12207 551
rect 12265 551 12299 561
rect 12265 527 12299 551
rect 12357 551 12391 561
rect 12357 527 12391 551
rect 12449 551 12483 561
rect 12449 527 12483 551
rect 12541 551 12575 561
rect 12541 527 12575 551
rect 12633 551 12667 561
rect 12633 527 12667 551
rect 12725 551 12759 561
rect 12725 527 12759 551
rect 12817 551 12851 561
rect 12817 527 12851 551
rect 12909 551 12943 561
rect 12909 527 12943 551
rect 13001 551 13035 561
rect 13001 527 13035 551
rect 13093 551 13127 561
rect 13093 527 13127 551
rect 13185 551 13219 561
rect 13185 527 13219 551
rect 13277 551 13311 561
rect 13277 527 13311 551
rect 13369 551 13403 561
rect 13369 527 13403 551
rect 13461 551 13495 561
rect 13461 527 13495 551
rect 13553 551 13587 561
rect 13553 527 13587 551
rect 13645 551 13679 561
rect 13645 527 13679 551
rect 13737 551 13771 561
rect 13737 527 13771 551
rect 13829 551 13863 561
rect 13829 527 13863 551
rect 13921 551 13955 561
rect 13921 527 13955 551
rect 14013 551 14047 561
rect 14013 527 14047 551
rect 14105 551 14139 561
rect 14105 527 14139 551
rect 14197 551 14231 561
rect 14197 527 14231 551
rect 14289 551 14323 561
rect 14289 527 14323 551
rect 14381 551 14415 561
rect 14381 527 14415 551
rect 14473 551 14507 561
rect 14473 527 14507 551
rect 14565 551 14599 561
rect 14565 527 14599 551
rect 14657 551 14691 561
rect 14657 527 14691 551
rect 14749 551 14783 561
rect 14749 527 14783 551
rect 14841 551 14875 561
rect 14841 527 14875 551
rect 14933 551 14967 561
rect 14933 527 14967 551
rect 15025 551 15059 561
rect 15025 527 15059 551
rect 15117 551 15151 561
rect 15117 527 15151 551
rect 15209 551 15243 561
rect 15209 527 15243 551
rect 15301 551 15335 561
rect 15301 527 15335 551
rect 15393 551 15427 561
rect 15393 527 15427 551
rect 15485 551 15519 561
rect 15485 527 15519 551
rect 15577 551 15611 561
rect 15577 527 15611 551
rect 15669 551 15703 561
rect 15669 527 15703 551
rect 15761 551 15795 561
rect 15761 527 15795 551
rect 15853 551 15887 561
rect 15853 527 15887 551
rect 15945 551 15979 561
rect 15945 527 15979 551
rect 16037 551 16071 561
rect 16037 527 16071 551
rect 16129 551 16163 561
rect 16129 527 16163 551
rect 16221 551 16255 561
rect 16221 527 16255 551
rect 16313 551 16347 561
rect 16313 527 16347 551
rect 16405 551 16439 561
rect 16405 527 16439 551
rect 16497 551 16531 561
rect 16497 527 16531 551
rect 16589 551 16623 561
rect 16589 527 16623 551
rect 16681 551 16715 561
rect 16681 527 16715 551
rect 16773 551 16807 561
rect 16773 527 16807 551
rect 16865 551 16899 561
rect 16865 527 16899 551
rect 16957 551 16991 561
rect 16957 527 16991 551
rect 17049 551 17083 561
rect 17049 527 17083 551
rect 17141 551 17175 561
rect 17141 527 17175 551
rect 17233 551 17267 561
rect 17233 527 17267 551
rect 17325 551 17359 561
rect 17325 527 17359 551
rect 17417 551 17451 561
rect 17417 527 17451 551
rect 17509 551 17543 561
rect 17509 527 17543 551
rect 17601 551 17635 561
rect 17601 527 17635 551
rect 17693 551 17727 561
rect 17693 527 17727 551
rect 17785 551 17819 561
rect 17785 527 17819 551
rect 17877 551 17911 561
rect 17877 527 17911 551
rect 17969 551 18003 561
rect 17969 527 18003 551
rect 18061 551 18095 561
rect 18061 527 18095 551
rect 18153 551 18187 561
rect 18153 527 18187 551
rect 18245 551 18279 561
rect 18245 527 18279 551
rect 18337 551 18371 561
rect 18337 527 18371 551
rect 18429 551 18463 561
rect 18429 527 18463 551
rect 18521 551 18555 561
rect 18521 527 18555 551
rect 18613 551 18647 561
rect 18613 527 18647 551
rect 18705 551 18739 561
rect 18705 527 18739 551
rect 18797 551 18831 561
rect 18797 527 18831 551
rect 18889 551 18923 561
rect 18889 527 18923 551
rect 18981 551 19015 561
rect 18981 527 19015 551
rect 19073 551 19107 561
rect 19073 527 19107 551
rect 19165 551 19199 561
rect 19165 527 19199 551
rect 19257 551 19291 561
rect 19257 527 19291 551
rect 19349 551 19383 561
rect 19349 527 19383 551
rect 19441 551 19475 561
rect 19441 527 19475 551
rect 19533 551 19567 561
rect 19533 527 19567 551
rect 19625 551 19659 561
rect 19625 527 19659 551
rect 19717 551 19751 561
rect 19717 527 19751 551
rect 19809 551 19843 561
rect 19809 527 19843 551
rect 19901 551 19935 561
rect 19901 527 19935 551
rect 19993 551 20027 561
rect 19993 527 20027 551
rect 20085 551 20119 561
rect 20085 527 20119 551
rect 20177 551 20211 561
rect 20177 527 20211 551
rect 20269 551 20303 561
rect 20269 527 20303 551
rect 20361 551 20395 561
rect 20361 527 20395 551
rect 20453 551 20487 561
rect 20453 527 20487 551
rect 20545 551 20579 561
rect 20545 527 20579 551
rect 20637 551 20671 561
rect 20637 527 20671 551
rect 20729 551 20763 561
rect 20729 527 20763 551
rect 20821 551 20855 561
rect 20821 527 20855 551
rect 20913 551 20947 561
rect 20913 527 20947 551
rect 21005 551 21039 561
rect 21005 527 21039 551
rect 21097 551 21131 561
rect 21097 527 21131 551
rect 21189 551 21223 561
rect 21189 527 21223 551
rect 21281 551 21315 561
rect 21281 527 21315 551
rect 21373 551 21407 561
rect 21373 527 21407 551
rect 21465 551 21499 561
rect 21465 527 21499 551
rect 21557 551 21591 561
rect 21557 527 21591 551
rect 21649 551 21683 561
rect 21649 527 21683 551
rect 21741 551 21775 561
rect 21741 527 21775 551
rect 21833 551 21867 561
rect 21833 527 21867 551
rect 21925 551 21959 561
rect 21925 527 21959 551
rect 22017 551 22051 561
rect 22017 527 22051 551
rect 22109 551 22143 561
rect 22109 527 22143 551
rect 22201 551 22235 561
rect 22201 527 22235 551
rect 22293 551 22327 561
rect 22293 527 22327 551
rect 22385 551 22419 561
rect 22385 527 22419 551
rect 22477 551 22511 561
rect 22477 527 22511 551
rect 22569 551 22603 561
rect 22569 527 22603 551
rect 22661 551 22695 561
rect 22661 527 22695 551
rect 22753 551 22787 561
rect 22753 527 22787 551
rect 22845 551 22879 561
rect 22845 527 22879 551
rect 22937 551 22971 561
rect 22937 527 22971 551
rect 23029 551 23063 561
rect 23029 527 23063 551
rect 23121 551 23155 561
rect 23121 527 23155 551
rect 23213 551 23247 561
rect 23213 527 23247 551
rect 23305 551 23339 561
rect 23305 527 23339 551
rect 23397 551 23431 561
rect 23397 527 23431 551
rect 23489 551 23523 561
rect 23489 527 23523 551
rect 23581 551 23615 561
rect 23581 527 23615 551
rect 23673 551 23707 561
rect 23673 527 23707 551
rect 23765 551 23799 561
rect 23765 527 23799 551
rect 23857 551 23891 561
rect 23857 527 23891 551
rect 23949 551 23983 561
rect 23949 527 23983 551
rect 24041 551 24075 561
rect 24041 527 24075 551
rect 24133 551 24167 561
rect 24133 527 24167 551
rect 24225 551 24259 561
rect 24225 527 24259 551
rect 24317 551 24351 561
rect 24317 527 24351 551
rect 24409 551 24443 561
rect 24409 527 24443 551
rect 24501 551 24535 561
rect 24501 527 24535 551
rect 24593 551 24627 561
rect 24593 527 24627 551
rect 24685 551 24719 561
rect 24685 527 24719 551
rect 24777 551 24811 561
rect 24777 527 24811 551
rect 24869 551 24903 561
rect 24869 527 24903 551
rect 24961 551 24995 561
rect 24961 527 24995 551
rect 25053 551 25087 561
rect 25053 527 25087 551
rect 25145 551 25179 561
rect 25145 527 25179 551
rect 25237 551 25271 561
rect 25237 527 25271 551
rect 25329 551 25363 561
rect 25329 527 25363 551
rect 25421 551 25455 561
rect 25421 527 25455 551
rect 25513 551 25547 561
rect 25513 527 25547 551
rect 25605 551 25639 561
rect 25605 527 25639 551
rect 25697 551 25731 561
rect 25697 527 25731 551
rect 25789 551 25823 561
rect 25789 527 25823 551
rect 25881 551 25915 561
rect 25881 527 25915 551
rect 25973 551 26007 561
rect 25973 527 26007 551
rect 26065 551 26099 561
rect 26065 527 26099 551
rect 26157 551 26191 561
rect 26157 527 26191 551
rect 26249 551 26283 561
rect 26249 527 26283 551
rect 26341 551 26375 561
rect 26341 527 26375 551
rect 26433 551 26467 561
rect 26433 527 26467 551
rect 26525 551 26559 561
rect 26525 527 26559 551
rect 26617 551 26651 561
rect 26617 527 26651 551
rect 26709 551 26743 561
rect 26709 527 26743 551
rect 26801 551 26835 561
rect 26801 527 26835 551
rect 26893 551 26927 561
rect 26893 527 26927 551
rect 26985 551 27019 561
rect 26985 527 27019 551
rect 27077 551 27111 561
rect 27077 527 27111 551
rect 27169 551 27203 561
rect 27169 527 27203 551
rect 27261 551 27295 561
rect 27261 527 27295 551
rect 27353 551 27387 561
rect 27353 527 27387 551
rect 27445 551 27479 561
rect 27445 527 27479 551
rect 27537 551 27571 561
rect 27537 527 27571 551
rect 27629 551 27663 561
rect 27629 527 27663 551
rect 27721 551 27755 561
rect 27721 527 27755 551
rect 27813 551 27847 561
rect 27813 527 27847 551
rect 27905 551 27939 561
rect 27905 527 27939 551
rect 27997 551 28031 561
rect 27997 527 28031 551
rect 28089 551 28123 561
rect 28089 527 28123 551
rect 28181 551 28215 561
rect 28181 527 28215 551
rect 28273 551 28307 561
rect 28273 527 28307 551
rect 28365 551 28399 561
rect 28365 527 28399 551
rect 28457 551 28491 561
rect 28457 527 28491 551
rect 28549 551 28583 561
rect 28549 527 28583 551
rect 28641 551 28675 561
rect 28641 527 28675 551
rect 28733 551 28767 561
rect 28733 527 28767 551
rect 28825 551 28859 561
rect 28825 527 28859 551
rect 28917 551 28951 561
rect 28917 527 28951 551
rect 29009 551 29043 561
rect 29009 527 29043 551
rect 29101 551 29135 561
rect 29101 527 29135 551
rect 29193 551 29227 561
rect 29193 527 29227 551
rect 29285 551 29319 561
rect 29285 527 29319 551
rect 29377 551 29411 561
rect 29377 527 29411 551
rect 29469 551 29503 561
rect 29469 527 29503 551
rect 29561 551 29595 561
rect 29561 527 29595 551
rect 29653 551 29687 561
rect 29653 527 29687 551
rect 29745 551 29779 561
rect 29745 527 29779 551
rect 29837 551 29871 561
rect 29837 527 29871 551
rect 29929 551 29963 561
rect 29929 527 29963 551
rect 30021 551 30055 561
rect 30021 527 30055 551
rect 30113 551 30147 561
rect 30113 527 30147 551
rect 30205 551 30239 561
rect 30205 527 30239 551
rect 30297 551 30331 561
rect 30297 527 30331 551
rect 30389 551 30423 561
rect 30389 527 30423 551
rect 30481 551 30515 561
rect 30481 527 30515 551
rect 30573 551 30607 561
rect 30573 527 30607 551
rect 30665 551 30699 561
rect 30665 527 30699 551
rect 30757 551 30791 561
rect 30757 527 30791 551
rect 30849 551 30883 561
rect 30849 527 30883 551
rect 30941 551 30975 561
rect 30941 527 30975 551
rect 31033 551 31067 561
rect 31033 527 31067 551
rect 31125 551 31159 561
rect 31125 527 31159 551
rect 31217 551 31251 561
rect 31217 527 31251 551
rect 31309 551 31343 561
rect 31309 527 31343 551
rect 31401 551 31435 561
rect 31401 527 31435 551
rect 31493 551 31527 561
rect 31493 527 31527 551
rect 31585 551 31619 561
rect 31585 527 31619 551
rect 31677 551 31711 561
rect 31677 527 31711 551
rect 31769 551 31803 561
rect 31769 527 31803 551
rect 31861 551 31895 561
rect 31861 527 31895 551
rect 31953 551 31987 561
rect 31953 527 31987 551
rect 32045 551 32079 561
rect 32045 527 32079 551
rect 32137 551 32171 561
rect 32137 527 32171 551
rect 32229 551 32263 561
rect 32229 527 32263 551
rect 32321 551 32355 561
rect 32321 527 32355 551
rect 32413 551 32447 561
rect 32413 527 32447 551
rect 32505 551 32539 561
rect 32505 527 32539 551
rect 32597 551 32631 561
rect 32597 527 32631 551
rect 32689 551 32723 561
rect 32689 527 32723 551
rect 32781 551 32815 561
rect 32781 527 32815 551
rect 32873 551 32907 561
rect 32873 527 32907 551
rect 32965 551 32999 561
rect 32965 527 32999 551
rect 33057 551 33091 561
rect 33057 527 33091 551
rect 33149 551 33183 561
rect 33149 527 33183 551
rect 33241 551 33275 561
rect 33241 527 33275 551
rect 33333 551 33367 561
rect 33333 527 33367 551
rect 33425 551 33459 561
rect 33425 527 33459 551
rect 33517 551 33551 561
rect 33517 527 33551 551
rect 33609 551 33643 561
rect 33609 527 33643 551
rect 33701 551 33735 561
rect 33701 527 33735 551
rect 33793 551 33827 561
rect 33793 527 33827 551
rect 33885 551 33919 561
rect 33885 527 33919 551
rect 33977 551 34011 561
rect 33977 527 34011 551
rect 34069 551 34103 561
rect 34069 527 34103 551
rect 34161 551 34195 561
rect 34161 527 34195 551
rect 34253 551 34287 561
rect 34253 527 34287 551
rect 34345 551 34379 561
rect 34345 527 34379 551
rect 34437 551 34471 561
rect 34437 527 34471 551
rect 34529 551 34563 561
rect 34529 527 34563 551
rect 34621 551 34655 561
rect 34621 527 34655 551
rect 34713 551 34747 561
rect 34713 527 34747 551
rect 34805 551 34839 561
rect 34805 527 34839 551
rect 34897 551 34931 561
rect 34897 527 34931 551
rect 34989 551 35023 561
rect 34989 527 35023 551
rect 35081 551 35115 561
rect 35081 527 35115 551
rect 35173 551 35207 561
rect 35173 527 35207 551
rect 35265 551 35299 561
rect 35265 527 35299 551
rect 35357 551 35391 561
rect 35357 527 35391 551
rect 35449 551 35483 561
rect 35449 527 35483 551
rect 35541 551 35575 561
rect 35541 527 35575 551
rect 35633 551 35667 561
rect 35633 527 35667 551
rect 35725 551 35759 561
rect 35725 527 35759 551
rect 35817 551 35851 561
rect 35817 527 35851 551
rect 35909 551 35943 561
rect 35909 527 35943 551
rect 36001 551 36035 561
rect 36001 527 36035 551
rect 36093 551 36127 561
rect 36093 527 36127 551
rect 36185 551 36219 561
rect 36185 527 36219 551
rect 36277 551 36311 561
rect 36277 527 36311 551
rect 36369 551 36403 561
rect 36369 527 36403 551
rect 36461 551 36495 561
rect 36461 527 36495 551
rect 36553 551 36587 561
rect 36553 527 36587 551
rect 36645 551 36679 561
rect 36645 527 36679 551
rect 36737 551 36771 561
rect 36737 527 36771 551
rect 36829 551 36863 561
rect 36829 527 36863 551
rect 36921 551 36955 561
rect 36921 527 36955 551
rect 37013 551 37047 561
rect 37013 527 37047 551
rect 37105 551 37139 561
rect 37105 527 37139 551
rect 37197 551 37231 561
rect 37197 527 37231 551
rect 37289 551 37323 561
rect 37289 527 37323 551
rect 37381 551 37415 561
rect 37381 527 37415 551
rect 37473 551 37507 561
rect 37473 527 37507 551
rect 37565 551 37599 561
rect 37565 527 37599 551
rect 37657 551 37691 561
rect 37657 527 37691 551
rect 37749 551 37783 561
rect 37749 527 37783 551
rect 37841 551 37875 561
rect 37841 527 37875 551
rect 37933 551 37967 561
rect 37933 527 37967 551
rect 38025 551 38059 561
rect 38025 527 38059 551
rect 38117 551 38151 561
rect 38117 527 38151 551
rect 38209 551 38243 561
rect 38209 527 38243 551
rect 38301 551 38335 561
rect 38301 527 38335 551
rect 38393 551 38427 561
rect 38393 527 38427 551
rect 38485 551 38519 561
rect 38485 527 38519 551
rect 38577 551 38611 561
rect 38577 527 38611 551
rect 38669 551 38703 561
rect 38669 527 38703 551
rect 38761 551 38795 561
rect 38761 527 38795 551
rect 38853 551 38887 561
rect 38853 527 38887 551
rect 38945 551 38979 561
rect 38945 527 38979 551
rect 39037 551 39071 561
rect 39037 527 39071 551
rect 39129 551 39163 561
rect 39129 527 39163 551
rect 39221 551 39255 561
rect 39221 527 39255 551
rect 39313 551 39347 561
rect 39313 527 39347 551
rect 39405 551 39439 561
rect 39405 527 39439 551
rect 39497 551 39531 561
rect 39497 527 39531 551
rect 39589 551 39623 561
rect 39589 527 39623 551
rect 39681 551 39715 561
rect 39681 527 39715 551
rect 39773 551 39807 561
rect 39773 527 39807 551
rect 39865 551 39899 561
rect 39865 527 39899 551
rect 39957 551 39991 561
rect 39957 527 39991 551
rect 40049 551 40083 561
rect 40049 527 40083 551
rect 40141 551 40175 561
rect 40141 527 40175 551
rect 40233 551 40267 561
rect 40233 527 40267 551
rect 40325 551 40359 561
rect 40325 527 40359 551
rect 40417 551 40451 561
rect 40417 527 40451 551
rect 40509 551 40543 561
rect 40509 527 40543 551
rect 40601 551 40635 561
rect 40601 527 40635 551
rect 40693 551 40727 561
rect 40693 527 40727 551
rect 40785 551 40819 561
rect 40785 527 40819 551
rect 40877 551 40911 561
rect 40877 527 40911 551
rect 40969 551 41003 561
rect 40969 527 41003 551
rect 41061 551 41095 561
rect 41061 527 41095 551
rect 41153 551 41187 561
rect 41153 527 41187 551
rect 41245 551 41279 561
rect 41245 527 41279 551
rect 41337 551 41371 561
rect 41337 527 41371 551
rect 41429 551 41463 561
rect 41429 527 41463 551
rect 41521 551 41555 561
rect 41521 527 41555 551
rect 41613 551 41647 561
rect 41613 527 41647 551
rect 41705 551 41739 561
rect 41705 527 41739 551
rect 41797 551 41831 561
rect 41797 527 41831 551
rect 41889 551 41923 561
rect 41889 527 41923 551
rect 41981 551 42015 561
rect 41981 527 42015 551
rect 42073 551 42107 561
rect 42073 527 42107 551
rect 42165 551 42199 561
rect 42165 527 42199 551
rect 42257 551 42291 561
rect 42257 527 42291 551
rect 122 230 134 255
rect 134 230 156 255
rect 122 221 156 230
rect 203 375 237 391
rect 203 357 237 375
rect 307 141 345 175
rect 581 357 615 391
rect 489 221 523 255
rect 1205 365 1239 391
rect 1205 357 1236 365
rect 1236 357 1239 365
rect 761 153 795 187
rect 833 169 857 187
rect 857 169 867 187
rect 833 153 867 169
rect 1205 239 1239 255
rect 1205 221 1231 239
rect 1231 221 1239 239
rect 1421 241 1455 250
rect 1421 216 1437 241
rect 1437 216 1455 241
rect 1481 153 1515 187
rect 2076 240 2114 274
rect 2238 230 2250 255
rect 2250 230 2272 255
rect 2238 221 2272 230
rect 2319 375 2353 391
rect 2319 357 2353 375
rect 2423 141 2461 175
rect 2697 357 2731 391
rect 2605 221 2639 255
rect 3321 365 3355 391
rect 3321 357 3352 365
rect 3352 357 3355 365
rect 2877 153 2911 187
rect 2949 169 2973 187
rect 2973 169 2983 187
rect 2949 153 2983 169
rect 3321 239 3355 255
rect 3321 221 3347 239
rect 3347 221 3355 239
rect 3537 241 3571 250
rect 3537 216 3553 241
rect 3553 216 3571 241
rect 3597 153 3631 187
rect 4192 240 4230 274
rect 4354 230 4366 255
rect 4366 230 4388 255
rect 4354 221 4388 230
rect 4435 375 4469 391
rect 4435 357 4469 375
rect 4539 141 4577 175
rect 4813 357 4847 391
rect 4721 221 4755 255
rect 5437 365 5471 391
rect 5437 357 5468 365
rect 5468 357 5471 365
rect 4993 153 5027 187
rect 5065 169 5089 187
rect 5089 169 5099 187
rect 5065 153 5099 169
rect 5437 239 5471 255
rect 5437 221 5463 239
rect 5463 221 5471 239
rect 5653 241 5687 250
rect 5653 216 5669 241
rect 5669 216 5687 241
rect 5713 153 5747 187
rect 6308 240 6346 274
rect 6470 230 6482 255
rect 6482 230 6504 255
rect 6470 221 6504 230
rect 6551 375 6585 391
rect 6551 357 6585 375
rect 6655 141 6693 175
rect 6929 357 6963 391
rect 6837 221 6871 255
rect 7553 365 7587 391
rect 7553 357 7584 365
rect 7584 357 7587 365
rect 7109 153 7143 187
rect 7181 169 7205 187
rect 7205 169 7215 187
rect 7181 153 7215 169
rect 7553 239 7587 255
rect 7553 221 7579 239
rect 7579 221 7587 239
rect 7769 241 7803 250
rect 7769 216 7785 241
rect 7785 216 7803 241
rect 7829 153 7863 187
rect 8424 240 8462 274
rect 8586 230 8598 255
rect 8598 230 8620 255
rect 8586 221 8620 230
rect 8667 375 8701 391
rect 8667 357 8701 375
rect 8771 141 8809 175
rect 9045 357 9079 391
rect 8953 221 8987 255
rect 9669 365 9703 391
rect 9669 357 9700 365
rect 9700 357 9703 365
rect 9225 153 9259 187
rect 9297 169 9321 187
rect 9321 169 9331 187
rect 9297 153 9331 169
rect 9669 239 9703 255
rect 9669 221 9695 239
rect 9695 221 9703 239
rect 9885 241 9919 250
rect 9885 216 9901 241
rect 9901 216 9919 241
rect 9945 153 9979 187
rect 10540 240 10578 274
rect 10702 230 10714 255
rect 10714 230 10736 255
rect 10702 221 10736 230
rect 10783 375 10817 391
rect 10783 357 10817 375
rect 10887 141 10925 175
rect 11161 357 11195 391
rect 11069 221 11103 255
rect 11785 365 11819 391
rect 11785 357 11816 365
rect 11816 357 11819 365
rect 11341 153 11375 187
rect 11413 169 11437 187
rect 11437 169 11447 187
rect 11413 153 11447 169
rect 11785 239 11819 255
rect 11785 221 11811 239
rect 11811 221 11819 239
rect 12001 241 12035 250
rect 12001 216 12017 241
rect 12017 216 12035 241
rect 12061 153 12095 187
rect 12656 240 12694 274
rect 12818 230 12830 255
rect 12830 230 12852 255
rect 12818 221 12852 230
rect 12899 375 12933 391
rect 12899 357 12933 375
rect 13003 141 13041 175
rect 13277 357 13311 391
rect 13185 221 13219 255
rect 13901 365 13935 391
rect 13901 357 13932 365
rect 13932 357 13935 365
rect 13457 153 13491 187
rect 13529 169 13553 187
rect 13553 169 13563 187
rect 13529 153 13563 169
rect 13901 239 13935 255
rect 13901 221 13927 239
rect 13927 221 13935 239
rect 14117 241 14151 250
rect 14117 216 14133 241
rect 14133 216 14151 241
rect 14177 153 14211 187
rect 14772 240 14810 274
rect 14934 230 14946 255
rect 14946 230 14968 255
rect 14934 221 14968 230
rect 15015 375 15049 391
rect 15015 357 15049 375
rect 15119 141 15157 175
rect 15393 357 15427 391
rect 15301 221 15335 255
rect 16017 365 16051 391
rect 16017 357 16048 365
rect 16048 357 16051 365
rect 15573 153 15607 187
rect 15645 169 15669 187
rect 15669 169 15679 187
rect 15645 153 15679 169
rect 16017 239 16051 255
rect 16017 221 16043 239
rect 16043 221 16051 239
rect 16233 241 16267 250
rect 16233 216 16249 241
rect 16249 216 16267 241
rect 16293 153 16327 187
rect 16888 240 16926 274
rect 17050 230 17062 255
rect 17062 230 17084 255
rect 17050 221 17084 230
rect 17131 375 17165 391
rect 17131 357 17165 375
rect 17235 141 17273 175
rect 17509 357 17543 391
rect 17417 221 17451 255
rect 18133 365 18167 391
rect 18133 357 18164 365
rect 18164 357 18167 365
rect 17689 153 17723 187
rect 17761 169 17785 187
rect 17785 169 17795 187
rect 17761 153 17795 169
rect 18133 239 18167 255
rect 18133 221 18159 239
rect 18159 221 18167 239
rect 18349 241 18383 250
rect 18349 216 18365 241
rect 18365 216 18383 241
rect 18409 153 18443 187
rect 19004 240 19042 274
rect 19166 230 19178 255
rect 19178 230 19200 255
rect 19166 221 19200 230
rect 19247 375 19281 391
rect 19247 357 19281 375
rect 19351 141 19389 175
rect 19625 357 19659 391
rect 19533 221 19567 255
rect 20249 365 20283 391
rect 20249 357 20280 365
rect 20280 357 20283 365
rect 19805 153 19839 187
rect 19877 169 19901 187
rect 19901 169 19911 187
rect 19877 153 19911 169
rect 20249 239 20283 255
rect 20249 221 20275 239
rect 20275 221 20283 239
rect 20465 241 20499 250
rect 20465 216 20481 241
rect 20481 216 20499 241
rect 20525 153 20559 187
rect 21120 240 21158 274
rect 21282 230 21294 255
rect 21294 230 21316 255
rect 21282 221 21316 230
rect 21363 375 21397 391
rect 21363 357 21397 375
rect 21467 141 21505 175
rect 21741 357 21775 391
rect 21649 221 21683 255
rect 22365 365 22399 391
rect 22365 357 22396 365
rect 22396 357 22399 365
rect 21921 153 21955 187
rect 21993 169 22017 187
rect 22017 169 22027 187
rect 21993 153 22027 169
rect 22365 239 22399 255
rect 22365 221 22391 239
rect 22391 221 22399 239
rect 22581 241 22615 250
rect 22581 216 22597 241
rect 22597 216 22615 241
rect 22641 153 22675 187
rect 23236 240 23274 274
rect 23398 230 23410 255
rect 23410 230 23432 255
rect 23398 221 23432 230
rect 23479 375 23513 391
rect 23479 357 23513 375
rect 23583 141 23621 175
rect 23857 357 23891 391
rect 23765 221 23799 255
rect 24481 365 24515 391
rect 24481 357 24512 365
rect 24512 357 24515 365
rect 24037 153 24071 187
rect 24109 169 24133 187
rect 24133 169 24143 187
rect 24109 153 24143 169
rect 24481 239 24515 255
rect 24481 221 24507 239
rect 24507 221 24515 239
rect 24697 241 24731 250
rect 24697 216 24713 241
rect 24713 216 24731 241
rect 24757 153 24791 187
rect 25352 240 25390 274
rect 25514 230 25526 255
rect 25526 230 25548 255
rect 25514 221 25548 230
rect 25595 375 25629 391
rect 25595 357 25629 375
rect 25699 141 25737 175
rect 25973 357 26007 391
rect 25881 221 25915 255
rect 26597 365 26631 391
rect 26597 357 26628 365
rect 26628 357 26631 365
rect 26153 153 26187 187
rect 26225 169 26249 187
rect 26249 169 26259 187
rect 26225 153 26259 169
rect 26597 239 26631 255
rect 26597 221 26623 239
rect 26623 221 26631 239
rect 26813 241 26847 250
rect 26813 216 26829 241
rect 26829 216 26847 241
rect 26873 153 26907 187
rect 27468 240 27506 274
rect 27630 230 27642 255
rect 27642 230 27664 255
rect 27630 221 27664 230
rect 27711 375 27745 391
rect 27711 357 27745 375
rect 27815 141 27853 175
rect 28089 357 28123 391
rect 27997 221 28031 255
rect 28713 365 28747 391
rect 28713 357 28744 365
rect 28744 357 28747 365
rect 28269 153 28303 187
rect 28341 169 28365 187
rect 28365 169 28375 187
rect 28341 153 28375 169
rect 28713 239 28747 255
rect 28713 221 28739 239
rect 28739 221 28747 239
rect 28929 241 28963 250
rect 28929 216 28945 241
rect 28945 216 28963 241
rect 28989 153 29023 187
rect 29584 240 29622 274
rect 29746 230 29758 255
rect 29758 230 29780 255
rect 29746 221 29780 230
rect 29827 375 29861 391
rect 29827 357 29861 375
rect 29931 141 29969 175
rect 30205 357 30239 391
rect 30113 221 30147 255
rect 30829 365 30863 391
rect 30829 357 30860 365
rect 30860 357 30863 365
rect 30385 153 30419 187
rect 30457 169 30481 187
rect 30481 169 30491 187
rect 30457 153 30491 169
rect 30829 239 30863 255
rect 30829 221 30855 239
rect 30855 221 30863 239
rect 31045 241 31079 250
rect 31045 216 31061 241
rect 31061 216 31079 241
rect 31105 153 31139 187
rect 31700 240 31738 274
rect 31862 230 31874 255
rect 31874 230 31896 255
rect 31862 221 31896 230
rect 31943 375 31977 391
rect 31943 357 31977 375
rect 32047 141 32085 175
rect 32321 357 32355 391
rect 32229 221 32263 255
rect 32945 365 32979 391
rect 32945 357 32976 365
rect 32976 357 32979 365
rect 32501 153 32535 187
rect 32573 169 32597 187
rect 32597 169 32607 187
rect 32573 153 32607 169
rect 32945 239 32979 255
rect 32945 221 32971 239
rect 32971 221 32979 239
rect 33161 241 33195 250
rect 33161 216 33177 241
rect 33177 216 33195 241
rect 33221 153 33255 187
rect 33816 240 33854 274
rect 33978 230 33990 255
rect 33990 230 34012 255
rect 33978 221 34012 230
rect 34059 375 34093 391
rect 34059 357 34093 375
rect 34163 141 34201 175
rect 34437 357 34471 391
rect 34345 221 34379 255
rect 35061 365 35095 391
rect 35061 357 35092 365
rect 35092 357 35095 365
rect 34617 153 34651 187
rect 34689 169 34713 187
rect 34713 169 34723 187
rect 34689 153 34723 169
rect 35061 239 35095 255
rect 35061 221 35087 239
rect 35087 221 35095 239
rect 35277 241 35311 250
rect 35277 216 35293 241
rect 35293 216 35311 241
rect 35337 153 35371 187
rect 35932 240 35970 274
rect 36094 230 36106 255
rect 36106 230 36128 255
rect 36094 221 36128 230
rect 36175 375 36209 391
rect 36175 357 36209 375
rect 36279 141 36317 175
rect 36553 357 36587 391
rect 36461 221 36495 255
rect 37177 365 37211 391
rect 37177 357 37208 365
rect 37208 357 37211 365
rect 36733 153 36767 187
rect 36805 169 36829 187
rect 36829 169 36839 187
rect 36805 153 36839 169
rect 37177 239 37211 255
rect 37177 221 37203 239
rect 37203 221 37211 239
rect 37393 241 37427 250
rect 37393 216 37409 241
rect 37409 216 37427 241
rect 37453 153 37487 187
rect 38048 240 38086 274
rect 38210 230 38222 255
rect 38222 230 38244 255
rect 38210 221 38244 230
rect 38291 375 38325 391
rect 38291 357 38325 375
rect 38395 141 38433 175
rect 38669 357 38703 391
rect 38577 221 38611 255
rect 39293 365 39327 391
rect 39293 357 39324 365
rect 39324 357 39327 365
rect 38849 153 38883 187
rect 38921 169 38945 187
rect 38945 169 38955 187
rect 38921 153 38955 169
rect 39293 239 39327 255
rect 39293 221 39319 239
rect 39319 221 39327 239
rect 39509 241 39543 250
rect 39509 216 39525 241
rect 39525 216 39543 241
rect 39569 153 39603 187
rect 40164 240 40202 274
rect 40326 230 40338 255
rect 40338 230 40360 255
rect 40326 221 40360 230
rect 40407 375 40441 391
rect 40407 357 40441 375
rect 40511 141 40549 175
rect 40785 357 40819 391
rect 40693 221 40727 255
rect 41409 365 41443 391
rect 41409 357 41440 365
rect 41440 357 41443 365
rect 40965 153 40999 187
rect 41037 169 41061 187
rect 41061 169 41071 187
rect 41037 153 41071 169
rect 41409 239 41443 255
rect 41409 221 41435 239
rect 41435 221 41443 239
rect 41625 241 41659 250
rect 41625 216 41641 241
rect 41641 216 41659 241
rect 41685 153 41719 187
rect 42280 240 42318 274
rect 29 -7 63 17
rect 29 -17 63 -7
rect 121 -7 155 17
rect 121 -17 155 -7
rect 213 -7 247 17
rect 213 -17 247 -7
rect 305 -7 339 17
rect 305 -17 339 -7
rect 397 -7 431 17
rect 397 -17 431 -7
rect 489 -7 523 17
rect 489 -17 523 -7
rect 581 -7 615 17
rect 581 -17 615 -7
rect 673 -7 707 17
rect 673 -17 707 -7
rect 765 -7 799 17
rect 765 -17 799 -7
rect 857 -7 891 17
rect 857 -17 891 -7
rect 949 -7 983 17
rect 949 -17 983 -7
rect 1041 -7 1075 17
rect 1041 -17 1075 -7
rect 1133 -7 1167 17
rect 1133 -17 1167 -7
rect 1225 -7 1259 17
rect 1225 -17 1259 -7
rect 1317 -7 1351 17
rect 1317 -17 1351 -7
rect 1409 -7 1443 17
rect 1409 -17 1443 -7
rect 1501 -7 1535 17
rect 1501 -17 1535 -7
rect 1593 -7 1627 17
rect 1593 -17 1627 -7
rect 1685 -7 1719 17
rect 1685 -17 1719 -7
rect 1777 -7 1811 17
rect 1777 -17 1811 -7
rect 1869 -7 1903 17
rect 1869 -17 1903 -7
rect 1961 -7 1995 17
rect 1961 -17 1995 -7
rect 2053 -7 2087 17
rect 2053 -17 2087 -7
rect 2145 -7 2179 17
rect 2145 -17 2179 -7
rect 2237 -7 2271 17
rect 2237 -17 2271 -7
rect 2329 -7 2363 17
rect 2329 -17 2363 -7
rect 2421 -7 2455 17
rect 2421 -17 2455 -7
rect 2513 -7 2547 17
rect 2513 -17 2547 -7
rect 2605 -7 2639 17
rect 2605 -17 2639 -7
rect 2697 -7 2731 17
rect 2697 -17 2731 -7
rect 2789 -7 2823 17
rect 2789 -17 2823 -7
rect 2881 -7 2915 17
rect 2881 -17 2915 -7
rect 2973 -7 3007 17
rect 2973 -17 3007 -7
rect 3065 -7 3099 17
rect 3065 -17 3099 -7
rect 3157 -7 3191 17
rect 3157 -17 3191 -7
rect 3249 -7 3283 17
rect 3249 -17 3283 -7
rect 3341 -7 3375 17
rect 3341 -17 3375 -7
rect 3433 -7 3467 17
rect 3433 -17 3467 -7
rect 3525 -7 3559 17
rect 3525 -17 3559 -7
rect 3617 -7 3651 17
rect 3617 -17 3651 -7
rect 3709 -7 3743 17
rect 3709 -17 3743 -7
rect 3801 -7 3835 17
rect 3801 -17 3835 -7
rect 3893 -7 3927 17
rect 3893 -17 3927 -7
rect 3985 -7 4019 17
rect 3985 -17 4019 -7
rect 4077 -7 4111 17
rect 4077 -17 4111 -7
rect 4169 -7 4203 17
rect 4169 -17 4203 -7
rect 4261 -7 4295 17
rect 4261 -17 4295 -7
rect 4353 -7 4387 17
rect 4353 -17 4387 -7
rect 4445 -7 4479 17
rect 4445 -17 4479 -7
rect 4537 -7 4571 17
rect 4537 -17 4571 -7
rect 4629 -7 4663 17
rect 4629 -17 4663 -7
rect 4721 -7 4755 17
rect 4721 -17 4755 -7
rect 4813 -7 4847 17
rect 4813 -17 4847 -7
rect 4905 -7 4939 17
rect 4905 -17 4939 -7
rect 4997 -7 5031 17
rect 4997 -17 5031 -7
rect 5089 -7 5123 17
rect 5089 -17 5123 -7
rect 5181 -7 5215 17
rect 5181 -17 5215 -7
rect 5273 -7 5307 17
rect 5273 -17 5307 -7
rect 5365 -7 5399 17
rect 5365 -17 5399 -7
rect 5457 -7 5491 17
rect 5457 -17 5491 -7
rect 5549 -7 5583 17
rect 5549 -17 5583 -7
rect 5641 -7 5675 17
rect 5641 -17 5675 -7
rect 5733 -7 5767 17
rect 5733 -17 5767 -7
rect 5825 -7 5859 17
rect 5825 -17 5859 -7
rect 5917 -7 5951 17
rect 5917 -17 5951 -7
rect 6009 -7 6043 17
rect 6009 -17 6043 -7
rect 6101 -7 6135 17
rect 6101 -17 6135 -7
rect 6193 -7 6227 17
rect 6193 -17 6227 -7
rect 6285 -7 6319 17
rect 6285 -17 6319 -7
rect 6377 -7 6411 17
rect 6377 -17 6411 -7
rect 6469 -7 6503 17
rect 6469 -17 6503 -7
rect 6561 -7 6595 17
rect 6561 -17 6595 -7
rect 6653 -7 6687 17
rect 6653 -17 6687 -7
rect 6745 -7 6779 17
rect 6745 -17 6779 -7
rect 6837 -7 6871 17
rect 6837 -17 6871 -7
rect 6929 -7 6963 17
rect 6929 -17 6963 -7
rect 7021 -7 7055 17
rect 7021 -17 7055 -7
rect 7113 -7 7147 17
rect 7113 -17 7147 -7
rect 7205 -7 7239 17
rect 7205 -17 7239 -7
rect 7297 -7 7331 17
rect 7297 -17 7331 -7
rect 7389 -7 7423 17
rect 7389 -17 7423 -7
rect 7481 -7 7515 17
rect 7481 -17 7515 -7
rect 7573 -7 7607 17
rect 7573 -17 7607 -7
rect 7665 -7 7699 17
rect 7665 -17 7699 -7
rect 7757 -7 7791 17
rect 7757 -17 7791 -7
rect 7849 -7 7883 17
rect 7849 -17 7883 -7
rect 7941 -7 7975 17
rect 7941 -17 7975 -7
rect 8033 -7 8067 17
rect 8033 -17 8067 -7
rect 8125 -7 8159 17
rect 8125 -17 8159 -7
rect 8217 -7 8251 17
rect 8217 -17 8251 -7
rect 8309 -7 8343 17
rect 8309 -17 8343 -7
rect 8401 -7 8435 17
rect 8401 -17 8435 -7
rect 8493 -7 8527 17
rect 8493 -17 8527 -7
rect 8585 -7 8619 17
rect 8585 -17 8619 -7
rect 8677 -7 8711 17
rect 8677 -17 8711 -7
rect 8769 -7 8803 17
rect 8769 -17 8803 -7
rect 8861 -7 8895 17
rect 8861 -17 8895 -7
rect 8953 -7 8987 17
rect 8953 -17 8987 -7
rect 9045 -7 9079 17
rect 9045 -17 9079 -7
rect 9137 -7 9171 17
rect 9137 -17 9171 -7
rect 9229 -7 9263 17
rect 9229 -17 9263 -7
rect 9321 -7 9355 17
rect 9321 -17 9355 -7
rect 9413 -7 9447 17
rect 9413 -17 9447 -7
rect 9505 -7 9539 17
rect 9505 -17 9539 -7
rect 9597 -7 9631 17
rect 9597 -17 9631 -7
rect 9689 -7 9723 17
rect 9689 -17 9723 -7
rect 9781 -7 9815 17
rect 9781 -17 9815 -7
rect 9873 -7 9907 17
rect 9873 -17 9907 -7
rect 9965 -7 9999 17
rect 9965 -17 9999 -7
rect 10057 -7 10091 17
rect 10057 -17 10091 -7
rect 10149 -7 10183 17
rect 10149 -17 10183 -7
rect 10241 -7 10275 17
rect 10241 -17 10275 -7
rect 10333 -7 10367 17
rect 10333 -17 10367 -7
rect 10425 -7 10459 17
rect 10425 -17 10459 -7
rect 10517 -7 10551 17
rect 10517 -17 10551 -7
rect 10609 -7 10643 17
rect 10609 -17 10643 -7
rect 10701 -7 10735 17
rect 10701 -17 10735 -7
rect 10793 -7 10827 17
rect 10793 -17 10827 -7
rect 10885 -7 10919 17
rect 10885 -17 10919 -7
rect 10977 -7 11011 17
rect 10977 -17 11011 -7
rect 11069 -7 11103 17
rect 11069 -17 11103 -7
rect 11161 -7 11195 17
rect 11161 -17 11195 -7
rect 11253 -7 11287 17
rect 11253 -17 11287 -7
rect 11345 -7 11379 17
rect 11345 -17 11379 -7
rect 11437 -7 11471 17
rect 11437 -17 11471 -7
rect 11529 -7 11563 17
rect 11529 -17 11563 -7
rect 11621 -7 11655 17
rect 11621 -17 11655 -7
rect 11713 -7 11747 17
rect 11713 -17 11747 -7
rect 11805 -7 11839 17
rect 11805 -17 11839 -7
rect 11897 -7 11931 17
rect 11897 -17 11931 -7
rect 11989 -7 12023 17
rect 11989 -17 12023 -7
rect 12081 -7 12115 17
rect 12081 -17 12115 -7
rect 12173 -7 12207 17
rect 12173 -17 12207 -7
rect 12265 -7 12299 17
rect 12265 -17 12299 -7
rect 12357 -7 12391 17
rect 12357 -17 12391 -7
rect 12449 -7 12483 17
rect 12449 -17 12483 -7
rect 12541 -7 12575 17
rect 12541 -17 12575 -7
rect 12633 -7 12667 17
rect 12633 -17 12667 -7
rect 12725 -7 12759 17
rect 12725 -17 12759 -7
rect 12817 -7 12851 17
rect 12817 -17 12851 -7
rect 12909 -7 12943 17
rect 12909 -17 12943 -7
rect 13001 -7 13035 17
rect 13001 -17 13035 -7
rect 13093 -7 13127 17
rect 13093 -17 13127 -7
rect 13185 -7 13219 17
rect 13185 -17 13219 -7
rect 13277 -7 13311 17
rect 13277 -17 13311 -7
rect 13369 -7 13403 17
rect 13369 -17 13403 -7
rect 13461 -7 13495 17
rect 13461 -17 13495 -7
rect 13553 -7 13587 17
rect 13553 -17 13587 -7
rect 13645 -7 13679 17
rect 13645 -17 13679 -7
rect 13737 -7 13771 17
rect 13737 -17 13771 -7
rect 13829 -7 13863 17
rect 13829 -17 13863 -7
rect 13921 -7 13955 17
rect 13921 -17 13955 -7
rect 14013 -7 14047 17
rect 14013 -17 14047 -7
rect 14105 -7 14139 17
rect 14105 -17 14139 -7
rect 14197 -7 14231 17
rect 14197 -17 14231 -7
rect 14289 -7 14323 17
rect 14289 -17 14323 -7
rect 14381 -7 14415 17
rect 14381 -17 14415 -7
rect 14473 -7 14507 17
rect 14473 -17 14507 -7
rect 14565 -7 14599 17
rect 14565 -17 14599 -7
rect 14657 -7 14691 17
rect 14657 -17 14691 -7
rect 14749 -7 14783 17
rect 14749 -17 14783 -7
rect 14841 -7 14875 17
rect 14841 -17 14875 -7
rect 14933 -7 14967 17
rect 14933 -17 14967 -7
rect 15025 -7 15059 17
rect 15025 -17 15059 -7
rect 15117 -7 15151 17
rect 15117 -17 15151 -7
rect 15209 -7 15243 17
rect 15209 -17 15243 -7
rect 15301 -7 15335 17
rect 15301 -17 15335 -7
rect 15393 -7 15427 17
rect 15393 -17 15427 -7
rect 15485 -7 15519 17
rect 15485 -17 15519 -7
rect 15577 -7 15611 17
rect 15577 -17 15611 -7
rect 15669 -7 15703 17
rect 15669 -17 15703 -7
rect 15761 -7 15795 17
rect 15761 -17 15795 -7
rect 15853 -7 15887 17
rect 15853 -17 15887 -7
rect 15945 -7 15979 17
rect 15945 -17 15979 -7
rect 16037 -7 16071 17
rect 16037 -17 16071 -7
rect 16129 -7 16163 17
rect 16129 -17 16163 -7
rect 16221 -7 16255 17
rect 16221 -17 16255 -7
rect 16313 -7 16347 17
rect 16313 -17 16347 -7
rect 16405 -7 16439 17
rect 16405 -17 16439 -7
rect 16497 -7 16531 17
rect 16497 -17 16531 -7
rect 16589 -7 16623 17
rect 16589 -17 16623 -7
rect 16681 -7 16715 17
rect 16681 -17 16715 -7
rect 16773 -7 16807 17
rect 16773 -17 16807 -7
rect 16865 -7 16899 17
rect 16865 -17 16899 -7
rect 16957 -7 16991 17
rect 16957 -17 16991 -7
rect 17049 -7 17083 17
rect 17049 -17 17083 -7
rect 17141 -7 17175 17
rect 17141 -17 17175 -7
rect 17233 -7 17267 17
rect 17233 -17 17267 -7
rect 17325 -7 17359 17
rect 17325 -17 17359 -7
rect 17417 -7 17451 17
rect 17417 -17 17451 -7
rect 17509 -7 17543 17
rect 17509 -17 17543 -7
rect 17601 -7 17635 17
rect 17601 -17 17635 -7
rect 17693 -7 17727 17
rect 17693 -17 17727 -7
rect 17785 -7 17819 17
rect 17785 -17 17819 -7
rect 17877 -7 17911 17
rect 17877 -17 17911 -7
rect 17969 -7 18003 17
rect 17969 -17 18003 -7
rect 18061 -7 18095 17
rect 18061 -17 18095 -7
rect 18153 -7 18187 17
rect 18153 -17 18187 -7
rect 18245 -7 18279 17
rect 18245 -17 18279 -7
rect 18337 -7 18371 17
rect 18337 -17 18371 -7
rect 18429 -7 18463 17
rect 18429 -17 18463 -7
rect 18521 -7 18555 17
rect 18521 -17 18555 -7
rect 18613 -7 18647 17
rect 18613 -17 18647 -7
rect 18705 -7 18739 17
rect 18705 -17 18739 -7
rect 18797 -7 18831 17
rect 18797 -17 18831 -7
rect 18889 -7 18923 17
rect 18889 -17 18923 -7
rect 18981 -7 19015 17
rect 18981 -17 19015 -7
rect 19073 -7 19107 17
rect 19073 -17 19107 -7
rect 19165 -7 19199 17
rect 19165 -17 19199 -7
rect 19257 -7 19291 17
rect 19257 -17 19291 -7
rect 19349 -7 19383 17
rect 19349 -17 19383 -7
rect 19441 -7 19475 17
rect 19441 -17 19475 -7
rect 19533 -7 19567 17
rect 19533 -17 19567 -7
rect 19625 -7 19659 17
rect 19625 -17 19659 -7
rect 19717 -7 19751 17
rect 19717 -17 19751 -7
rect 19809 -7 19843 17
rect 19809 -17 19843 -7
rect 19901 -7 19935 17
rect 19901 -17 19935 -7
rect 19993 -7 20027 17
rect 19993 -17 20027 -7
rect 20085 -7 20119 17
rect 20085 -17 20119 -7
rect 20177 -7 20211 17
rect 20177 -17 20211 -7
rect 20269 -7 20303 17
rect 20269 -17 20303 -7
rect 20361 -7 20395 17
rect 20361 -17 20395 -7
rect 20453 -7 20487 17
rect 20453 -17 20487 -7
rect 20545 -7 20579 17
rect 20545 -17 20579 -7
rect 20637 -7 20671 17
rect 20637 -17 20671 -7
rect 20729 -7 20763 17
rect 20729 -17 20763 -7
rect 20821 -7 20855 17
rect 20821 -17 20855 -7
rect 20913 -7 20947 17
rect 20913 -17 20947 -7
rect 21005 -7 21039 17
rect 21005 -17 21039 -7
rect 21097 -7 21131 17
rect 21097 -17 21131 -7
rect 21189 -7 21223 17
rect 21189 -17 21223 -7
rect 21281 -7 21315 17
rect 21281 -17 21315 -7
rect 21373 -7 21407 17
rect 21373 -17 21407 -7
rect 21465 -7 21499 17
rect 21465 -17 21499 -7
rect 21557 -7 21591 17
rect 21557 -17 21591 -7
rect 21649 -7 21683 17
rect 21649 -17 21683 -7
rect 21741 -7 21775 17
rect 21741 -17 21775 -7
rect 21833 -7 21867 17
rect 21833 -17 21867 -7
rect 21925 -7 21959 17
rect 21925 -17 21959 -7
rect 22017 -7 22051 17
rect 22017 -17 22051 -7
rect 22109 -7 22143 17
rect 22109 -17 22143 -7
rect 22201 -7 22235 17
rect 22201 -17 22235 -7
rect 22293 -7 22327 17
rect 22293 -17 22327 -7
rect 22385 -7 22419 17
rect 22385 -17 22419 -7
rect 22477 -7 22511 17
rect 22477 -17 22511 -7
rect 22569 -7 22603 17
rect 22569 -17 22603 -7
rect 22661 -7 22695 17
rect 22661 -17 22695 -7
rect 22753 -7 22787 17
rect 22753 -17 22787 -7
rect 22845 -7 22879 17
rect 22845 -17 22879 -7
rect 22937 -7 22971 17
rect 22937 -17 22971 -7
rect 23029 -7 23063 17
rect 23029 -17 23063 -7
rect 23121 -7 23155 17
rect 23121 -17 23155 -7
rect 23213 -7 23247 17
rect 23213 -17 23247 -7
rect 23305 -7 23339 17
rect 23305 -17 23339 -7
rect 23397 -7 23431 17
rect 23397 -17 23431 -7
rect 23489 -7 23523 17
rect 23489 -17 23523 -7
rect 23581 -7 23615 17
rect 23581 -17 23615 -7
rect 23673 -7 23707 17
rect 23673 -17 23707 -7
rect 23765 -7 23799 17
rect 23765 -17 23799 -7
rect 23857 -7 23891 17
rect 23857 -17 23891 -7
rect 23949 -7 23983 17
rect 23949 -17 23983 -7
rect 24041 -7 24075 17
rect 24041 -17 24075 -7
rect 24133 -7 24167 17
rect 24133 -17 24167 -7
rect 24225 -7 24259 17
rect 24225 -17 24259 -7
rect 24317 -7 24351 17
rect 24317 -17 24351 -7
rect 24409 -7 24443 17
rect 24409 -17 24443 -7
rect 24501 -7 24535 17
rect 24501 -17 24535 -7
rect 24593 -7 24627 17
rect 24593 -17 24627 -7
rect 24685 -7 24719 17
rect 24685 -17 24719 -7
rect 24777 -7 24811 17
rect 24777 -17 24811 -7
rect 24869 -7 24903 17
rect 24869 -17 24903 -7
rect 24961 -7 24995 17
rect 24961 -17 24995 -7
rect 25053 -7 25087 17
rect 25053 -17 25087 -7
rect 25145 -7 25179 17
rect 25145 -17 25179 -7
rect 25237 -7 25271 17
rect 25237 -17 25271 -7
rect 25329 -7 25363 17
rect 25329 -17 25363 -7
rect 25421 -7 25455 17
rect 25421 -17 25455 -7
rect 25513 -7 25547 17
rect 25513 -17 25547 -7
rect 25605 -7 25639 17
rect 25605 -17 25639 -7
rect 25697 -7 25731 17
rect 25697 -17 25731 -7
rect 25789 -7 25823 17
rect 25789 -17 25823 -7
rect 25881 -7 25915 17
rect 25881 -17 25915 -7
rect 25973 -7 26007 17
rect 25973 -17 26007 -7
rect 26065 -7 26099 17
rect 26065 -17 26099 -7
rect 26157 -7 26191 17
rect 26157 -17 26191 -7
rect 26249 -7 26283 17
rect 26249 -17 26283 -7
rect 26341 -7 26375 17
rect 26341 -17 26375 -7
rect 26433 -7 26467 17
rect 26433 -17 26467 -7
rect 26525 -7 26559 17
rect 26525 -17 26559 -7
rect 26617 -7 26651 17
rect 26617 -17 26651 -7
rect 26709 -7 26743 17
rect 26709 -17 26743 -7
rect 26801 -7 26835 17
rect 26801 -17 26835 -7
rect 26893 -7 26927 17
rect 26893 -17 26927 -7
rect 26985 -7 27019 17
rect 26985 -17 27019 -7
rect 27077 -7 27111 17
rect 27077 -17 27111 -7
rect 27169 -7 27203 17
rect 27169 -17 27203 -7
rect 27261 -7 27295 17
rect 27261 -17 27295 -7
rect 27353 -7 27387 17
rect 27353 -17 27387 -7
rect 27445 -7 27479 17
rect 27445 -17 27479 -7
rect 27537 -7 27571 17
rect 27537 -17 27571 -7
rect 27629 -7 27663 17
rect 27629 -17 27663 -7
rect 27721 -7 27755 17
rect 27721 -17 27755 -7
rect 27813 -7 27847 17
rect 27813 -17 27847 -7
rect 27905 -7 27939 17
rect 27905 -17 27939 -7
rect 27997 -7 28031 17
rect 27997 -17 28031 -7
rect 28089 -7 28123 17
rect 28089 -17 28123 -7
rect 28181 -7 28215 17
rect 28181 -17 28215 -7
rect 28273 -7 28307 17
rect 28273 -17 28307 -7
rect 28365 -7 28399 17
rect 28365 -17 28399 -7
rect 28457 -7 28491 17
rect 28457 -17 28491 -7
rect 28549 -7 28583 17
rect 28549 -17 28583 -7
rect 28641 -7 28675 17
rect 28641 -17 28675 -7
rect 28733 -7 28767 17
rect 28733 -17 28767 -7
rect 28825 -7 28859 17
rect 28825 -17 28859 -7
rect 28917 -7 28951 17
rect 28917 -17 28951 -7
rect 29009 -7 29043 17
rect 29009 -17 29043 -7
rect 29101 -7 29135 17
rect 29101 -17 29135 -7
rect 29193 -7 29227 17
rect 29193 -17 29227 -7
rect 29285 -7 29319 17
rect 29285 -17 29319 -7
rect 29377 -7 29411 17
rect 29377 -17 29411 -7
rect 29469 -7 29503 17
rect 29469 -17 29503 -7
rect 29561 -7 29595 17
rect 29561 -17 29595 -7
rect 29653 -7 29687 17
rect 29653 -17 29687 -7
rect 29745 -7 29779 17
rect 29745 -17 29779 -7
rect 29837 -7 29871 17
rect 29837 -17 29871 -7
rect 29929 -7 29963 17
rect 29929 -17 29963 -7
rect 30021 -7 30055 17
rect 30021 -17 30055 -7
rect 30113 -7 30147 17
rect 30113 -17 30147 -7
rect 30205 -7 30239 17
rect 30205 -17 30239 -7
rect 30297 -7 30331 17
rect 30297 -17 30331 -7
rect 30389 -7 30423 17
rect 30389 -17 30423 -7
rect 30481 -7 30515 17
rect 30481 -17 30515 -7
rect 30573 -7 30607 17
rect 30573 -17 30607 -7
rect 30665 -7 30699 17
rect 30665 -17 30699 -7
rect 30757 -7 30791 17
rect 30757 -17 30791 -7
rect 30849 -7 30883 17
rect 30849 -17 30883 -7
rect 30941 -7 30975 17
rect 30941 -17 30975 -7
rect 31033 -7 31067 17
rect 31033 -17 31067 -7
rect 31125 -7 31159 17
rect 31125 -17 31159 -7
rect 31217 -7 31251 17
rect 31217 -17 31251 -7
rect 31309 -7 31343 17
rect 31309 -17 31343 -7
rect 31401 -7 31435 17
rect 31401 -17 31435 -7
rect 31493 -7 31527 17
rect 31493 -17 31527 -7
rect 31585 -7 31619 17
rect 31585 -17 31619 -7
rect 31677 -7 31711 17
rect 31677 -17 31711 -7
rect 31769 -7 31803 17
rect 31769 -17 31803 -7
rect 31861 -7 31895 17
rect 31861 -17 31895 -7
rect 31953 -7 31987 17
rect 31953 -17 31987 -7
rect 32045 -7 32079 17
rect 32045 -17 32079 -7
rect 32137 -7 32171 17
rect 32137 -17 32171 -7
rect 32229 -7 32263 17
rect 32229 -17 32263 -7
rect 32321 -7 32355 17
rect 32321 -17 32355 -7
rect 32413 -7 32447 17
rect 32413 -17 32447 -7
rect 32505 -7 32539 17
rect 32505 -17 32539 -7
rect 32597 -7 32631 17
rect 32597 -17 32631 -7
rect 32689 -7 32723 17
rect 32689 -17 32723 -7
rect 32781 -7 32815 17
rect 32781 -17 32815 -7
rect 32873 -7 32907 17
rect 32873 -17 32907 -7
rect 32965 -7 32999 17
rect 32965 -17 32999 -7
rect 33057 -7 33091 17
rect 33057 -17 33091 -7
rect 33149 -7 33183 17
rect 33149 -17 33183 -7
rect 33241 -7 33275 17
rect 33241 -17 33275 -7
rect 33333 -7 33367 17
rect 33333 -17 33367 -7
rect 33425 -7 33459 17
rect 33425 -17 33459 -7
rect 33517 -7 33551 17
rect 33517 -17 33551 -7
rect 33609 -7 33643 17
rect 33609 -17 33643 -7
rect 33701 -7 33735 17
rect 33701 -17 33735 -7
rect 33793 -7 33827 17
rect 33793 -17 33827 -7
rect 33885 -7 33919 17
rect 33885 -17 33919 -7
rect 33977 -7 34011 17
rect 33977 -17 34011 -7
rect 34069 -7 34103 17
rect 34069 -17 34103 -7
rect 34161 -7 34195 17
rect 34161 -17 34195 -7
rect 34253 -7 34287 17
rect 34253 -17 34287 -7
rect 34345 -7 34379 17
rect 34345 -17 34379 -7
rect 34437 -7 34471 17
rect 34437 -17 34471 -7
rect 34529 -7 34563 17
rect 34529 -17 34563 -7
rect 34621 -7 34655 17
rect 34621 -17 34655 -7
rect 34713 -7 34747 17
rect 34713 -17 34747 -7
rect 34805 -7 34839 17
rect 34805 -17 34839 -7
rect 34897 -7 34931 17
rect 34897 -17 34931 -7
rect 34989 -7 35023 17
rect 34989 -17 35023 -7
rect 35081 -7 35115 17
rect 35081 -17 35115 -7
rect 35173 -7 35207 17
rect 35173 -17 35207 -7
rect 35265 -7 35299 17
rect 35265 -17 35299 -7
rect 35357 -7 35391 17
rect 35357 -17 35391 -7
rect 35449 -7 35483 17
rect 35449 -17 35483 -7
rect 35541 -7 35575 17
rect 35541 -17 35575 -7
rect 35633 -7 35667 17
rect 35633 -17 35667 -7
rect 35725 -7 35759 17
rect 35725 -17 35759 -7
rect 35817 -7 35851 17
rect 35817 -17 35851 -7
rect 35909 -7 35943 17
rect 35909 -17 35943 -7
rect 36001 -7 36035 17
rect 36001 -17 36035 -7
rect 36093 -7 36127 17
rect 36093 -17 36127 -7
rect 36185 -7 36219 17
rect 36185 -17 36219 -7
rect 36277 -7 36311 17
rect 36277 -17 36311 -7
rect 36369 -7 36403 17
rect 36369 -17 36403 -7
rect 36461 -7 36495 17
rect 36461 -17 36495 -7
rect 36553 -7 36587 17
rect 36553 -17 36587 -7
rect 36645 -7 36679 17
rect 36645 -17 36679 -7
rect 36737 -7 36771 17
rect 36737 -17 36771 -7
rect 36829 -7 36863 17
rect 36829 -17 36863 -7
rect 36921 -7 36955 17
rect 36921 -17 36955 -7
rect 37013 -7 37047 17
rect 37013 -17 37047 -7
rect 37105 -7 37139 17
rect 37105 -17 37139 -7
rect 37197 -7 37231 17
rect 37197 -17 37231 -7
rect 37289 -7 37323 17
rect 37289 -17 37323 -7
rect 37381 -7 37415 17
rect 37381 -17 37415 -7
rect 37473 -7 37507 17
rect 37473 -17 37507 -7
rect 37565 -7 37599 17
rect 37565 -17 37599 -7
rect 37657 -7 37691 17
rect 37657 -17 37691 -7
rect 37749 -7 37783 17
rect 37749 -17 37783 -7
rect 37841 -7 37875 17
rect 37841 -17 37875 -7
rect 37933 -7 37967 17
rect 37933 -17 37967 -7
rect 38025 -7 38059 17
rect 38025 -17 38059 -7
rect 38117 -7 38151 17
rect 38117 -17 38151 -7
rect 38209 -7 38243 17
rect 38209 -17 38243 -7
rect 38301 -7 38335 17
rect 38301 -17 38335 -7
rect 38393 -7 38427 17
rect 38393 -17 38427 -7
rect 38485 -7 38519 17
rect 38485 -17 38519 -7
rect 38577 -7 38611 17
rect 38577 -17 38611 -7
rect 38669 -7 38703 17
rect 38669 -17 38703 -7
rect 38761 -7 38795 17
rect 38761 -17 38795 -7
rect 38853 -7 38887 17
rect 38853 -17 38887 -7
rect 38945 -7 38979 17
rect 38945 -17 38979 -7
rect 39037 -7 39071 17
rect 39037 -17 39071 -7
rect 39129 -7 39163 17
rect 39129 -17 39163 -7
rect 39221 -7 39255 17
rect 39221 -17 39255 -7
rect 39313 -7 39347 17
rect 39313 -17 39347 -7
rect 39405 -7 39439 17
rect 39405 -17 39439 -7
rect 39497 -7 39531 17
rect 39497 -17 39531 -7
rect 39589 -7 39623 17
rect 39589 -17 39623 -7
rect 39681 -7 39715 17
rect 39681 -17 39715 -7
rect 39773 -7 39807 17
rect 39773 -17 39807 -7
rect 39865 -7 39899 17
rect 39865 -17 39899 -7
rect 39957 -7 39991 17
rect 39957 -17 39991 -7
rect 40049 -7 40083 17
rect 40049 -17 40083 -7
rect 40141 -7 40175 17
rect 40141 -17 40175 -7
rect 40233 -7 40267 17
rect 40233 -17 40267 -7
rect 40325 -7 40359 17
rect 40325 -17 40359 -7
rect 40417 -7 40451 17
rect 40417 -17 40451 -7
rect 40509 -7 40543 17
rect 40509 -17 40543 -7
rect 40601 -7 40635 17
rect 40601 -17 40635 -7
rect 40693 -7 40727 17
rect 40693 -17 40727 -7
rect 40785 -7 40819 17
rect 40785 -17 40819 -7
rect 40877 -7 40911 17
rect 40877 -17 40911 -7
rect 40969 -7 41003 17
rect 40969 -17 41003 -7
rect 41061 -7 41095 17
rect 41061 -17 41095 -7
rect 41153 -7 41187 17
rect 41153 -17 41187 -7
rect 41245 -7 41279 17
rect 41245 -17 41279 -7
rect 41337 -7 41371 17
rect 41337 -17 41371 -7
rect 41429 -7 41463 17
rect 41429 -17 41463 -7
rect 41521 -7 41555 17
rect 41521 -17 41555 -7
rect 41613 -7 41647 17
rect 41613 -17 41647 -7
rect 41705 -7 41739 17
rect 41705 -17 41739 -7
rect 41797 -7 41831 17
rect 41797 -17 41831 -7
rect 41889 -7 41923 17
rect 41889 -17 41923 -7
rect 41981 -7 42015 17
rect 41981 -17 42015 -7
rect 42073 -7 42107 17
rect 42073 -17 42107 -7
rect 42165 -7 42199 17
rect 42165 -17 42199 -7
rect 42257 -7 42291 17
rect 42257 -17 42291 -7
<< metal1 >>
rect 0 561 42320 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2697 561
rect 2731 527 2789 561
rect 2823 527 2881 561
rect 2915 527 2973 561
rect 3007 527 3065 561
rect 3099 527 3157 561
rect 3191 527 3249 561
rect 3283 527 3341 561
rect 3375 527 3433 561
rect 3467 527 3525 561
rect 3559 527 3617 561
rect 3651 527 3709 561
rect 3743 527 3801 561
rect 3835 527 3893 561
rect 3927 527 3985 561
rect 4019 527 4077 561
rect 4111 527 4169 561
rect 4203 527 4261 561
rect 4295 527 4353 561
rect 4387 527 4445 561
rect 4479 527 4537 561
rect 4571 527 4629 561
rect 4663 527 4721 561
rect 4755 527 4813 561
rect 4847 527 4905 561
rect 4939 527 4997 561
rect 5031 527 5089 561
rect 5123 527 5181 561
rect 5215 527 5273 561
rect 5307 527 5365 561
rect 5399 527 5457 561
rect 5491 527 5549 561
rect 5583 527 5641 561
rect 5675 527 5733 561
rect 5767 527 5825 561
rect 5859 527 5917 561
rect 5951 527 6009 561
rect 6043 527 6101 561
rect 6135 527 6193 561
rect 6227 527 6285 561
rect 6319 527 6377 561
rect 6411 527 6469 561
rect 6503 527 6561 561
rect 6595 527 6653 561
rect 6687 527 6745 561
rect 6779 527 6837 561
rect 6871 527 6929 561
rect 6963 527 7021 561
rect 7055 527 7113 561
rect 7147 527 7205 561
rect 7239 527 7297 561
rect 7331 527 7389 561
rect 7423 527 7481 561
rect 7515 527 7573 561
rect 7607 527 7665 561
rect 7699 527 7757 561
rect 7791 527 7849 561
rect 7883 527 7941 561
rect 7975 527 8033 561
rect 8067 527 8125 561
rect 8159 527 8217 561
rect 8251 527 8309 561
rect 8343 527 8401 561
rect 8435 527 8493 561
rect 8527 527 8585 561
rect 8619 527 8677 561
rect 8711 527 8769 561
rect 8803 527 8861 561
rect 8895 527 8953 561
rect 8987 527 9045 561
rect 9079 527 9137 561
rect 9171 527 9229 561
rect 9263 527 9321 561
rect 9355 527 9413 561
rect 9447 527 9505 561
rect 9539 527 9597 561
rect 9631 527 9689 561
rect 9723 527 9781 561
rect 9815 527 9873 561
rect 9907 527 9965 561
rect 9999 527 10057 561
rect 10091 527 10149 561
rect 10183 527 10241 561
rect 10275 527 10333 561
rect 10367 527 10425 561
rect 10459 527 10517 561
rect 10551 527 10609 561
rect 10643 527 10701 561
rect 10735 527 10793 561
rect 10827 527 10885 561
rect 10919 527 10977 561
rect 11011 527 11069 561
rect 11103 527 11161 561
rect 11195 527 11253 561
rect 11287 527 11345 561
rect 11379 527 11437 561
rect 11471 527 11529 561
rect 11563 527 11621 561
rect 11655 527 11713 561
rect 11747 527 11805 561
rect 11839 527 11897 561
rect 11931 527 11989 561
rect 12023 527 12081 561
rect 12115 527 12173 561
rect 12207 527 12265 561
rect 12299 527 12357 561
rect 12391 527 12449 561
rect 12483 527 12541 561
rect 12575 527 12633 561
rect 12667 527 12725 561
rect 12759 527 12817 561
rect 12851 527 12909 561
rect 12943 527 13001 561
rect 13035 527 13093 561
rect 13127 527 13185 561
rect 13219 527 13277 561
rect 13311 527 13369 561
rect 13403 527 13461 561
rect 13495 527 13553 561
rect 13587 527 13645 561
rect 13679 527 13737 561
rect 13771 527 13829 561
rect 13863 527 13921 561
rect 13955 527 14013 561
rect 14047 527 14105 561
rect 14139 527 14197 561
rect 14231 527 14289 561
rect 14323 527 14381 561
rect 14415 527 14473 561
rect 14507 527 14565 561
rect 14599 527 14657 561
rect 14691 527 14749 561
rect 14783 527 14841 561
rect 14875 527 14933 561
rect 14967 527 15025 561
rect 15059 527 15117 561
rect 15151 527 15209 561
rect 15243 527 15301 561
rect 15335 527 15393 561
rect 15427 527 15485 561
rect 15519 527 15577 561
rect 15611 527 15669 561
rect 15703 527 15761 561
rect 15795 527 15853 561
rect 15887 527 15945 561
rect 15979 527 16037 561
rect 16071 527 16129 561
rect 16163 527 16221 561
rect 16255 527 16313 561
rect 16347 527 16405 561
rect 16439 527 16497 561
rect 16531 527 16589 561
rect 16623 527 16681 561
rect 16715 527 16773 561
rect 16807 527 16865 561
rect 16899 527 16957 561
rect 16991 527 17049 561
rect 17083 527 17141 561
rect 17175 527 17233 561
rect 17267 527 17325 561
rect 17359 527 17417 561
rect 17451 527 17509 561
rect 17543 527 17601 561
rect 17635 527 17693 561
rect 17727 527 17785 561
rect 17819 527 17877 561
rect 17911 527 17969 561
rect 18003 527 18061 561
rect 18095 527 18153 561
rect 18187 527 18245 561
rect 18279 527 18337 561
rect 18371 527 18429 561
rect 18463 527 18521 561
rect 18555 527 18613 561
rect 18647 527 18705 561
rect 18739 527 18797 561
rect 18831 527 18889 561
rect 18923 527 18981 561
rect 19015 527 19073 561
rect 19107 527 19165 561
rect 19199 527 19257 561
rect 19291 527 19349 561
rect 19383 527 19441 561
rect 19475 527 19533 561
rect 19567 527 19625 561
rect 19659 527 19717 561
rect 19751 527 19809 561
rect 19843 527 19901 561
rect 19935 527 19993 561
rect 20027 527 20085 561
rect 20119 527 20177 561
rect 20211 527 20269 561
rect 20303 527 20361 561
rect 20395 527 20453 561
rect 20487 527 20545 561
rect 20579 527 20637 561
rect 20671 527 20729 561
rect 20763 527 20821 561
rect 20855 527 20913 561
rect 20947 527 21005 561
rect 21039 527 21097 561
rect 21131 527 21189 561
rect 21223 527 21281 561
rect 21315 527 21373 561
rect 21407 527 21465 561
rect 21499 527 21557 561
rect 21591 527 21649 561
rect 21683 527 21741 561
rect 21775 527 21833 561
rect 21867 527 21925 561
rect 21959 527 22017 561
rect 22051 527 22109 561
rect 22143 527 22201 561
rect 22235 527 22293 561
rect 22327 527 22385 561
rect 22419 527 22477 561
rect 22511 527 22569 561
rect 22603 527 22661 561
rect 22695 527 22753 561
rect 22787 527 22845 561
rect 22879 527 22937 561
rect 22971 527 23029 561
rect 23063 527 23121 561
rect 23155 527 23213 561
rect 23247 527 23305 561
rect 23339 527 23397 561
rect 23431 527 23489 561
rect 23523 527 23581 561
rect 23615 527 23673 561
rect 23707 527 23765 561
rect 23799 527 23857 561
rect 23891 527 23949 561
rect 23983 527 24041 561
rect 24075 527 24133 561
rect 24167 527 24225 561
rect 24259 527 24317 561
rect 24351 527 24409 561
rect 24443 527 24501 561
rect 24535 527 24593 561
rect 24627 527 24685 561
rect 24719 527 24777 561
rect 24811 527 24869 561
rect 24903 527 24961 561
rect 24995 527 25053 561
rect 25087 527 25145 561
rect 25179 527 25237 561
rect 25271 527 25329 561
rect 25363 527 25421 561
rect 25455 527 25513 561
rect 25547 527 25605 561
rect 25639 527 25697 561
rect 25731 527 25789 561
rect 25823 527 25881 561
rect 25915 527 25973 561
rect 26007 527 26065 561
rect 26099 527 26157 561
rect 26191 527 26249 561
rect 26283 527 26341 561
rect 26375 527 26433 561
rect 26467 527 26525 561
rect 26559 527 26617 561
rect 26651 527 26709 561
rect 26743 527 26801 561
rect 26835 527 26893 561
rect 26927 527 26985 561
rect 27019 527 27077 561
rect 27111 527 27169 561
rect 27203 527 27261 561
rect 27295 527 27353 561
rect 27387 527 27445 561
rect 27479 527 27537 561
rect 27571 527 27629 561
rect 27663 527 27721 561
rect 27755 527 27813 561
rect 27847 527 27905 561
rect 27939 527 27997 561
rect 28031 527 28089 561
rect 28123 527 28181 561
rect 28215 527 28273 561
rect 28307 527 28365 561
rect 28399 527 28457 561
rect 28491 527 28549 561
rect 28583 527 28641 561
rect 28675 527 28733 561
rect 28767 527 28825 561
rect 28859 527 28917 561
rect 28951 527 29009 561
rect 29043 527 29101 561
rect 29135 527 29193 561
rect 29227 527 29285 561
rect 29319 527 29377 561
rect 29411 527 29469 561
rect 29503 527 29561 561
rect 29595 527 29653 561
rect 29687 527 29745 561
rect 29779 527 29837 561
rect 29871 527 29929 561
rect 29963 527 30021 561
rect 30055 527 30113 561
rect 30147 527 30205 561
rect 30239 527 30297 561
rect 30331 527 30389 561
rect 30423 527 30481 561
rect 30515 527 30573 561
rect 30607 527 30665 561
rect 30699 527 30757 561
rect 30791 527 30849 561
rect 30883 527 30941 561
rect 30975 527 31033 561
rect 31067 527 31125 561
rect 31159 527 31217 561
rect 31251 527 31309 561
rect 31343 527 31401 561
rect 31435 527 31493 561
rect 31527 527 31585 561
rect 31619 527 31677 561
rect 31711 527 31769 561
rect 31803 527 31861 561
rect 31895 527 31953 561
rect 31987 527 32045 561
rect 32079 527 32137 561
rect 32171 527 32229 561
rect 32263 527 32321 561
rect 32355 527 32413 561
rect 32447 527 32505 561
rect 32539 527 32597 561
rect 32631 527 32689 561
rect 32723 527 32781 561
rect 32815 527 32873 561
rect 32907 527 32965 561
rect 32999 527 33057 561
rect 33091 527 33149 561
rect 33183 527 33241 561
rect 33275 527 33333 561
rect 33367 527 33425 561
rect 33459 527 33517 561
rect 33551 527 33609 561
rect 33643 527 33701 561
rect 33735 527 33793 561
rect 33827 527 33885 561
rect 33919 527 33977 561
rect 34011 527 34069 561
rect 34103 527 34161 561
rect 34195 527 34253 561
rect 34287 527 34345 561
rect 34379 527 34437 561
rect 34471 527 34529 561
rect 34563 527 34621 561
rect 34655 527 34713 561
rect 34747 527 34805 561
rect 34839 527 34897 561
rect 34931 527 34989 561
rect 35023 527 35081 561
rect 35115 527 35173 561
rect 35207 527 35265 561
rect 35299 527 35357 561
rect 35391 527 35449 561
rect 35483 527 35541 561
rect 35575 527 35633 561
rect 35667 527 35725 561
rect 35759 527 35817 561
rect 35851 527 35909 561
rect 35943 527 36001 561
rect 36035 527 36093 561
rect 36127 527 36185 561
rect 36219 527 36277 561
rect 36311 527 36369 561
rect 36403 527 36461 561
rect 36495 527 36553 561
rect 36587 527 36645 561
rect 36679 527 36737 561
rect 36771 527 36829 561
rect 36863 527 36921 561
rect 36955 527 37013 561
rect 37047 527 37105 561
rect 37139 527 37197 561
rect 37231 527 37289 561
rect 37323 527 37381 561
rect 37415 527 37473 561
rect 37507 527 37565 561
rect 37599 527 37657 561
rect 37691 527 37749 561
rect 37783 527 37841 561
rect 37875 527 37933 561
rect 37967 527 38025 561
rect 38059 527 38117 561
rect 38151 527 38209 561
rect 38243 527 38301 561
rect 38335 527 38393 561
rect 38427 527 38485 561
rect 38519 527 38577 561
rect 38611 527 38669 561
rect 38703 527 38761 561
rect 38795 527 38853 561
rect 38887 527 38945 561
rect 38979 527 39037 561
rect 39071 527 39129 561
rect 39163 527 39221 561
rect 39255 527 39313 561
rect 39347 527 39405 561
rect 39439 527 39497 561
rect 39531 527 39589 561
rect 39623 527 39681 561
rect 39715 527 39773 561
rect 39807 527 39865 561
rect 39899 527 39957 561
rect 39991 527 40049 561
rect 40083 527 40141 561
rect 40175 527 40233 561
rect 40267 527 40325 561
rect 40359 527 40417 561
rect 40451 527 40509 561
rect 40543 527 40601 561
rect 40635 527 40693 561
rect 40727 527 40785 561
rect 40819 527 40877 561
rect 40911 527 40969 561
rect 41003 527 41061 561
rect 41095 527 41153 561
rect 41187 527 41245 561
rect 41279 527 41337 561
rect 41371 527 41429 561
rect 41463 527 41521 561
rect 41555 527 41613 561
rect 41647 527 41705 561
rect 41739 527 41797 561
rect 41831 527 41889 561
rect 41923 527 41981 561
rect 42015 527 42073 561
rect 42107 527 42165 561
rect 42199 527 42257 561
rect 42291 527 42320 561
rect 0 496 42320 527
rect 191 391 249 397
rect 191 357 203 391
rect 237 388 249 391
rect 569 391 627 397
rect 569 388 581 391
rect 237 360 581 388
rect 237 357 249 360
rect 191 351 249 357
rect 569 357 581 360
rect 615 388 627 391
rect 1193 391 1251 397
rect 1193 388 1205 391
rect 615 360 1205 388
rect 615 357 627 360
rect 569 351 627 357
rect 1193 357 1205 360
rect 1239 357 1251 391
rect 1193 351 1251 357
rect 2307 391 2365 397
rect 2307 357 2319 391
rect 2353 388 2365 391
rect 2685 391 2743 397
rect 2685 388 2697 391
rect 2353 360 2697 388
rect 2353 357 2365 360
rect 2307 351 2365 357
rect 2685 357 2697 360
rect 2731 388 2743 391
rect 3309 391 3367 397
rect 3309 388 3321 391
rect 2731 360 3321 388
rect 2731 357 2743 360
rect 2685 351 2743 357
rect 3309 357 3321 360
rect 3355 357 3367 391
rect 3309 351 3367 357
rect 4423 391 4481 397
rect 4423 357 4435 391
rect 4469 388 4481 391
rect 4801 391 4859 397
rect 4801 388 4813 391
rect 4469 360 4813 388
rect 4469 357 4481 360
rect 4423 351 4481 357
rect 4801 357 4813 360
rect 4847 388 4859 391
rect 5425 391 5483 397
rect 5425 388 5437 391
rect 4847 360 5437 388
rect 4847 357 4859 360
rect 4801 351 4859 357
rect 5425 357 5437 360
rect 5471 357 5483 391
rect 5425 351 5483 357
rect 6539 391 6597 397
rect 6539 357 6551 391
rect 6585 388 6597 391
rect 6917 391 6975 397
rect 6917 388 6929 391
rect 6585 360 6929 388
rect 6585 357 6597 360
rect 6539 351 6597 357
rect 6917 357 6929 360
rect 6963 388 6975 391
rect 7541 391 7599 397
rect 7541 388 7553 391
rect 6963 360 7553 388
rect 6963 357 6975 360
rect 6917 351 6975 357
rect 7541 357 7553 360
rect 7587 357 7599 391
rect 7541 351 7599 357
rect 8655 391 8713 397
rect 8655 357 8667 391
rect 8701 388 8713 391
rect 9033 391 9091 397
rect 9033 388 9045 391
rect 8701 360 9045 388
rect 8701 357 8713 360
rect 8655 351 8713 357
rect 9033 357 9045 360
rect 9079 388 9091 391
rect 9657 391 9715 397
rect 9657 388 9669 391
rect 9079 360 9669 388
rect 9079 357 9091 360
rect 9033 351 9091 357
rect 9657 357 9669 360
rect 9703 357 9715 391
rect 9657 351 9715 357
rect 10771 391 10829 397
rect 10771 357 10783 391
rect 10817 388 10829 391
rect 11149 391 11207 397
rect 11149 388 11161 391
rect 10817 360 11161 388
rect 10817 357 10829 360
rect 10771 351 10829 357
rect 11149 357 11161 360
rect 11195 388 11207 391
rect 11773 391 11831 397
rect 11773 388 11785 391
rect 11195 360 11785 388
rect 11195 357 11207 360
rect 11149 351 11207 357
rect 11773 357 11785 360
rect 11819 357 11831 391
rect 11773 351 11831 357
rect 12887 391 12945 397
rect 12887 357 12899 391
rect 12933 388 12945 391
rect 13265 391 13323 397
rect 13265 388 13277 391
rect 12933 360 13277 388
rect 12933 357 12945 360
rect 12887 351 12945 357
rect 13265 357 13277 360
rect 13311 388 13323 391
rect 13889 391 13947 397
rect 13889 388 13901 391
rect 13311 360 13901 388
rect 13311 357 13323 360
rect 13265 351 13323 357
rect 13889 357 13901 360
rect 13935 357 13947 391
rect 13889 351 13947 357
rect 15003 391 15061 397
rect 15003 357 15015 391
rect 15049 388 15061 391
rect 15381 391 15439 397
rect 15381 388 15393 391
rect 15049 360 15393 388
rect 15049 357 15061 360
rect 15003 351 15061 357
rect 15381 357 15393 360
rect 15427 388 15439 391
rect 16005 391 16063 397
rect 16005 388 16017 391
rect 15427 360 16017 388
rect 15427 357 15439 360
rect 15381 351 15439 357
rect 16005 357 16017 360
rect 16051 357 16063 391
rect 16005 351 16063 357
rect 17119 391 17177 397
rect 17119 357 17131 391
rect 17165 388 17177 391
rect 17497 391 17555 397
rect 17497 388 17509 391
rect 17165 360 17509 388
rect 17165 357 17177 360
rect 17119 351 17177 357
rect 17497 357 17509 360
rect 17543 388 17555 391
rect 18121 391 18179 397
rect 18121 388 18133 391
rect 17543 360 18133 388
rect 17543 357 17555 360
rect 17497 351 17555 357
rect 18121 357 18133 360
rect 18167 357 18179 391
rect 18121 351 18179 357
rect 19235 391 19293 397
rect 19235 357 19247 391
rect 19281 388 19293 391
rect 19613 391 19671 397
rect 19613 388 19625 391
rect 19281 360 19625 388
rect 19281 357 19293 360
rect 19235 351 19293 357
rect 19613 357 19625 360
rect 19659 388 19671 391
rect 20237 391 20295 397
rect 20237 388 20249 391
rect 19659 360 20249 388
rect 19659 357 19671 360
rect 19613 351 19671 357
rect 20237 357 20249 360
rect 20283 357 20295 391
rect 20237 351 20295 357
rect 21351 391 21409 397
rect 21351 357 21363 391
rect 21397 388 21409 391
rect 21729 391 21787 397
rect 21729 388 21741 391
rect 21397 360 21741 388
rect 21397 357 21409 360
rect 21351 351 21409 357
rect 21729 357 21741 360
rect 21775 388 21787 391
rect 22353 391 22411 397
rect 22353 388 22365 391
rect 21775 360 22365 388
rect 21775 357 21787 360
rect 21729 351 21787 357
rect 22353 357 22365 360
rect 22399 357 22411 391
rect 22353 351 22411 357
rect 23467 391 23525 397
rect 23467 357 23479 391
rect 23513 388 23525 391
rect 23845 391 23903 397
rect 23845 388 23857 391
rect 23513 360 23857 388
rect 23513 357 23525 360
rect 23467 351 23525 357
rect 23845 357 23857 360
rect 23891 388 23903 391
rect 24469 391 24527 397
rect 24469 388 24481 391
rect 23891 360 24481 388
rect 23891 357 23903 360
rect 23845 351 23903 357
rect 24469 357 24481 360
rect 24515 357 24527 391
rect 24469 351 24527 357
rect 25583 391 25641 397
rect 25583 357 25595 391
rect 25629 388 25641 391
rect 25961 391 26019 397
rect 25961 388 25973 391
rect 25629 360 25973 388
rect 25629 357 25641 360
rect 25583 351 25641 357
rect 25961 357 25973 360
rect 26007 388 26019 391
rect 26585 391 26643 397
rect 26585 388 26597 391
rect 26007 360 26597 388
rect 26007 357 26019 360
rect 25961 351 26019 357
rect 26585 357 26597 360
rect 26631 357 26643 391
rect 26585 351 26643 357
rect 27699 391 27757 397
rect 27699 357 27711 391
rect 27745 388 27757 391
rect 28077 391 28135 397
rect 28077 388 28089 391
rect 27745 360 28089 388
rect 27745 357 27757 360
rect 27699 351 27757 357
rect 28077 357 28089 360
rect 28123 388 28135 391
rect 28701 391 28759 397
rect 28701 388 28713 391
rect 28123 360 28713 388
rect 28123 357 28135 360
rect 28077 351 28135 357
rect 28701 357 28713 360
rect 28747 357 28759 391
rect 28701 351 28759 357
rect 29815 391 29873 397
rect 29815 357 29827 391
rect 29861 388 29873 391
rect 30193 391 30251 397
rect 30193 388 30205 391
rect 29861 360 30205 388
rect 29861 357 29873 360
rect 29815 351 29873 357
rect 30193 357 30205 360
rect 30239 388 30251 391
rect 30817 391 30875 397
rect 30817 388 30829 391
rect 30239 360 30829 388
rect 30239 357 30251 360
rect 30193 351 30251 357
rect 30817 357 30829 360
rect 30863 357 30875 391
rect 30817 351 30875 357
rect 31931 391 31989 397
rect 31931 357 31943 391
rect 31977 388 31989 391
rect 32309 391 32367 397
rect 32309 388 32321 391
rect 31977 360 32321 388
rect 31977 357 31989 360
rect 31931 351 31989 357
rect 32309 357 32321 360
rect 32355 388 32367 391
rect 32933 391 32991 397
rect 32933 388 32945 391
rect 32355 360 32945 388
rect 32355 357 32367 360
rect 32309 351 32367 357
rect 32933 357 32945 360
rect 32979 357 32991 391
rect 32933 351 32991 357
rect 34047 391 34105 397
rect 34047 357 34059 391
rect 34093 388 34105 391
rect 34425 391 34483 397
rect 34425 388 34437 391
rect 34093 360 34437 388
rect 34093 357 34105 360
rect 34047 351 34105 357
rect 34425 357 34437 360
rect 34471 388 34483 391
rect 35049 391 35107 397
rect 35049 388 35061 391
rect 34471 360 35061 388
rect 34471 357 34483 360
rect 34425 351 34483 357
rect 35049 357 35061 360
rect 35095 357 35107 391
rect 35049 351 35107 357
rect 36163 391 36221 397
rect 36163 357 36175 391
rect 36209 388 36221 391
rect 36541 391 36599 397
rect 36541 388 36553 391
rect 36209 360 36553 388
rect 36209 357 36221 360
rect 36163 351 36221 357
rect 36541 357 36553 360
rect 36587 388 36599 391
rect 37165 391 37223 397
rect 37165 388 37177 391
rect 36587 360 37177 388
rect 36587 357 36599 360
rect 36541 351 36599 357
rect 37165 357 37177 360
rect 37211 357 37223 391
rect 37165 351 37223 357
rect 38279 391 38337 397
rect 38279 357 38291 391
rect 38325 388 38337 391
rect 38657 391 38715 397
rect 38657 388 38669 391
rect 38325 360 38669 388
rect 38325 357 38337 360
rect 38279 351 38337 357
rect 38657 357 38669 360
rect 38703 388 38715 391
rect 39281 391 39339 397
rect 39281 388 39293 391
rect 38703 360 39293 388
rect 38703 357 38715 360
rect 38657 351 38715 357
rect 39281 357 39293 360
rect 39327 357 39339 391
rect 39281 351 39339 357
rect 40395 391 40453 397
rect 40395 357 40407 391
rect 40441 388 40453 391
rect 40773 391 40831 397
rect 40773 388 40785 391
rect 40441 360 40785 388
rect 40441 357 40453 360
rect 40395 351 40453 357
rect 40773 357 40785 360
rect 40819 388 40831 391
rect 41397 391 41455 397
rect 41397 388 41409 391
rect 40819 360 41409 388
rect 40819 357 40831 360
rect 40773 351 40831 357
rect 41397 357 41409 360
rect 41443 357 41455 391
rect 41397 351 41455 357
rect 1409 294 1529 300
rect 110 255 168 261
rect 110 221 122 255
rect 156 252 168 255
rect 477 255 535 261
rect 477 252 489 255
rect 156 224 489 252
rect 156 221 168 224
rect 110 215 168 221
rect 477 221 489 224
rect 523 252 535 255
rect 1193 255 1251 261
rect 1193 252 1205 255
rect 523 224 1205 252
rect 523 221 535 224
rect 477 215 535 221
rect 1193 221 1205 224
rect 1239 221 1251 255
rect 1193 215 1251 221
rect 1409 250 1433 294
rect 1409 216 1421 250
rect 1485 242 1529 294
rect 1455 216 1529 242
rect 249 183 418 191
rect 249 131 300 183
rect 352 131 418 183
rect 749 187 879 193
rect 749 153 761 187
rect 795 153 833 187
rect 867 184 879 187
rect 1409 187 1529 216
rect 2045 282 2138 309
rect 2045 230 2069 282
rect 2121 230 2138 282
rect 3525 294 3645 300
rect 2045 208 2138 230
rect 2226 255 2284 261
rect 2226 221 2238 255
rect 2272 252 2284 255
rect 2593 255 2651 261
rect 2593 252 2605 255
rect 2272 224 2605 252
rect 2272 221 2284 224
rect 2226 215 2284 221
rect 2593 221 2605 224
rect 2639 252 2651 255
rect 3309 255 3367 261
rect 3309 252 3321 255
rect 2639 224 3321 252
rect 2639 221 2651 224
rect 2593 215 2651 221
rect 3309 221 3321 224
rect 3355 221 3367 255
rect 3309 215 3367 221
rect 3525 250 3549 294
rect 3525 216 3537 250
rect 3601 242 3645 294
rect 3571 216 3645 242
rect 1409 184 1481 187
rect 867 156 1481 184
rect 867 153 879 156
rect 749 147 879 153
rect 1469 153 1481 156
rect 1515 184 1529 187
rect 1515 153 1527 184
rect 1469 147 1527 153
rect 2365 183 2534 191
rect 249 122 418 131
rect 2365 131 2416 183
rect 2468 131 2534 183
rect 2865 187 2995 193
rect 2865 153 2877 187
rect 2911 153 2949 187
rect 2983 184 2995 187
rect 3525 187 3645 216
rect 4161 282 4254 309
rect 4161 230 4185 282
rect 4237 230 4254 282
rect 5641 294 5761 300
rect 4161 208 4254 230
rect 4342 255 4400 261
rect 4342 221 4354 255
rect 4388 252 4400 255
rect 4709 255 4767 261
rect 4709 252 4721 255
rect 4388 224 4721 252
rect 4388 221 4400 224
rect 4342 215 4400 221
rect 4709 221 4721 224
rect 4755 252 4767 255
rect 5425 255 5483 261
rect 5425 252 5437 255
rect 4755 224 5437 252
rect 4755 221 4767 224
rect 4709 215 4767 221
rect 5425 221 5437 224
rect 5471 221 5483 255
rect 5425 215 5483 221
rect 5641 250 5665 294
rect 5641 216 5653 250
rect 5717 242 5761 294
rect 5687 216 5761 242
rect 3525 184 3597 187
rect 2983 156 3597 184
rect 2983 153 2995 156
rect 2865 147 2995 153
rect 3585 153 3597 156
rect 3631 184 3645 187
rect 3631 153 3643 184
rect 3585 147 3643 153
rect 4481 183 4650 191
rect 2365 122 2534 131
rect 4481 131 4532 183
rect 4584 131 4650 183
rect 4981 187 5111 193
rect 4981 153 4993 187
rect 5027 153 5065 187
rect 5099 184 5111 187
rect 5641 187 5761 216
rect 6277 282 6370 309
rect 6277 230 6301 282
rect 6353 230 6370 282
rect 7757 294 7877 300
rect 6277 208 6370 230
rect 6458 255 6516 261
rect 6458 221 6470 255
rect 6504 252 6516 255
rect 6825 255 6883 261
rect 6825 252 6837 255
rect 6504 224 6837 252
rect 6504 221 6516 224
rect 6458 215 6516 221
rect 6825 221 6837 224
rect 6871 252 6883 255
rect 7541 255 7599 261
rect 7541 252 7553 255
rect 6871 224 7553 252
rect 6871 221 6883 224
rect 6825 215 6883 221
rect 7541 221 7553 224
rect 7587 221 7599 255
rect 7541 215 7599 221
rect 7757 250 7781 294
rect 7757 216 7769 250
rect 7833 242 7877 294
rect 7803 216 7877 242
rect 5641 184 5713 187
rect 5099 156 5713 184
rect 5099 153 5111 156
rect 4981 147 5111 153
rect 5701 153 5713 156
rect 5747 184 5761 187
rect 5747 153 5759 184
rect 5701 147 5759 153
rect 6597 183 6766 191
rect 4481 122 4650 131
rect 6597 131 6648 183
rect 6700 131 6766 183
rect 7097 187 7227 193
rect 7097 153 7109 187
rect 7143 153 7181 187
rect 7215 184 7227 187
rect 7757 187 7877 216
rect 8393 282 8486 309
rect 8393 230 8417 282
rect 8469 230 8486 282
rect 9873 294 9993 300
rect 8393 208 8486 230
rect 8574 255 8632 261
rect 8574 221 8586 255
rect 8620 252 8632 255
rect 8941 255 8999 261
rect 8941 252 8953 255
rect 8620 224 8953 252
rect 8620 221 8632 224
rect 8574 215 8632 221
rect 8941 221 8953 224
rect 8987 252 8999 255
rect 9657 255 9715 261
rect 9657 252 9669 255
rect 8987 224 9669 252
rect 8987 221 8999 224
rect 8941 215 8999 221
rect 9657 221 9669 224
rect 9703 221 9715 255
rect 9657 215 9715 221
rect 9873 250 9897 294
rect 9873 216 9885 250
rect 9949 242 9993 294
rect 9919 216 9993 242
rect 7757 184 7829 187
rect 7215 156 7829 184
rect 7215 153 7227 156
rect 7097 147 7227 153
rect 7817 153 7829 156
rect 7863 184 7877 187
rect 7863 153 7875 184
rect 7817 147 7875 153
rect 8713 183 8882 191
rect 6597 122 6766 131
rect 8713 131 8764 183
rect 8816 131 8882 183
rect 9213 187 9343 193
rect 9213 153 9225 187
rect 9259 153 9297 187
rect 9331 184 9343 187
rect 9873 187 9993 216
rect 10509 282 10602 309
rect 10509 230 10533 282
rect 10585 230 10602 282
rect 11989 294 12109 300
rect 10509 208 10602 230
rect 10690 255 10748 261
rect 10690 221 10702 255
rect 10736 252 10748 255
rect 11057 255 11115 261
rect 11057 252 11069 255
rect 10736 224 11069 252
rect 10736 221 10748 224
rect 10690 215 10748 221
rect 11057 221 11069 224
rect 11103 252 11115 255
rect 11773 255 11831 261
rect 11773 252 11785 255
rect 11103 224 11785 252
rect 11103 221 11115 224
rect 11057 215 11115 221
rect 11773 221 11785 224
rect 11819 221 11831 255
rect 11773 215 11831 221
rect 11989 250 12013 294
rect 11989 216 12001 250
rect 12065 242 12109 294
rect 12035 216 12109 242
rect 9873 184 9945 187
rect 9331 156 9945 184
rect 9331 153 9343 156
rect 9213 147 9343 153
rect 9933 153 9945 156
rect 9979 184 9993 187
rect 9979 153 9991 184
rect 9933 147 9991 153
rect 10829 183 10998 191
rect 8713 122 8882 131
rect 10829 131 10880 183
rect 10932 131 10998 183
rect 11329 187 11459 193
rect 11329 153 11341 187
rect 11375 153 11413 187
rect 11447 184 11459 187
rect 11989 187 12109 216
rect 12625 282 12718 309
rect 12625 230 12649 282
rect 12701 230 12718 282
rect 14105 294 14225 300
rect 12625 208 12718 230
rect 12806 255 12864 261
rect 12806 221 12818 255
rect 12852 252 12864 255
rect 13173 255 13231 261
rect 13173 252 13185 255
rect 12852 224 13185 252
rect 12852 221 12864 224
rect 12806 215 12864 221
rect 13173 221 13185 224
rect 13219 252 13231 255
rect 13889 255 13947 261
rect 13889 252 13901 255
rect 13219 224 13901 252
rect 13219 221 13231 224
rect 13173 215 13231 221
rect 13889 221 13901 224
rect 13935 221 13947 255
rect 13889 215 13947 221
rect 14105 250 14129 294
rect 14105 216 14117 250
rect 14181 242 14225 294
rect 14151 216 14225 242
rect 11989 184 12061 187
rect 11447 156 12061 184
rect 11447 153 11459 156
rect 11329 147 11459 153
rect 12049 153 12061 156
rect 12095 184 12109 187
rect 12095 153 12107 184
rect 12049 147 12107 153
rect 12945 183 13114 191
rect 10829 122 10998 131
rect 12945 131 12996 183
rect 13048 131 13114 183
rect 13445 187 13575 193
rect 13445 153 13457 187
rect 13491 153 13529 187
rect 13563 184 13575 187
rect 14105 187 14225 216
rect 14741 282 14834 309
rect 14741 230 14765 282
rect 14817 230 14834 282
rect 16221 294 16341 300
rect 14741 208 14834 230
rect 14922 255 14980 261
rect 14922 221 14934 255
rect 14968 252 14980 255
rect 15289 255 15347 261
rect 15289 252 15301 255
rect 14968 224 15301 252
rect 14968 221 14980 224
rect 14922 215 14980 221
rect 15289 221 15301 224
rect 15335 252 15347 255
rect 16005 255 16063 261
rect 16005 252 16017 255
rect 15335 224 16017 252
rect 15335 221 15347 224
rect 15289 215 15347 221
rect 16005 221 16017 224
rect 16051 221 16063 255
rect 16005 215 16063 221
rect 16221 250 16245 294
rect 16221 216 16233 250
rect 16297 242 16341 294
rect 16267 216 16341 242
rect 14105 184 14177 187
rect 13563 156 14177 184
rect 13563 153 13575 156
rect 13445 147 13575 153
rect 14165 153 14177 156
rect 14211 184 14225 187
rect 14211 153 14223 184
rect 14165 147 14223 153
rect 15061 183 15230 191
rect 12945 122 13114 131
rect 15061 131 15112 183
rect 15164 131 15230 183
rect 15561 187 15691 193
rect 15561 153 15573 187
rect 15607 153 15645 187
rect 15679 184 15691 187
rect 16221 187 16341 216
rect 16857 282 16950 309
rect 16857 230 16881 282
rect 16933 230 16950 282
rect 18337 294 18457 300
rect 16857 208 16950 230
rect 17038 255 17096 261
rect 17038 221 17050 255
rect 17084 252 17096 255
rect 17405 255 17463 261
rect 17405 252 17417 255
rect 17084 224 17417 252
rect 17084 221 17096 224
rect 17038 215 17096 221
rect 17405 221 17417 224
rect 17451 252 17463 255
rect 18121 255 18179 261
rect 18121 252 18133 255
rect 17451 224 18133 252
rect 17451 221 17463 224
rect 17405 215 17463 221
rect 18121 221 18133 224
rect 18167 221 18179 255
rect 18121 215 18179 221
rect 18337 250 18361 294
rect 18337 216 18349 250
rect 18413 242 18457 294
rect 18383 216 18457 242
rect 16221 184 16293 187
rect 15679 156 16293 184
rect 15679 153 15691 156
rect 15561 147 15691 153
rect 16281 153 16293 156
rect 16327 184 16341 187
rect 16327 153 16339 184
rect 16281 147 16339 153
rect 17177 183 17346 191
rect 15061 122 15230 131
rect 17177 131 17228 183
rect 17280 131 17346 183
rect 17677 187 17807 193
rect 17677 153 17689 187
rect 17723 153 17761 187
rect 17795 184 17807 187
rect 18337 187 18457 216
rect 18973 282 19066 309
rect 18973 230 18997 282
rect 19049 230 19066 282
rect 20453 294 20573 300
rect 18973 208 19066 230
rect 19154 255 19212 261
rect 19154 221 19166 255
rect 19200 252 19212 255
rect 19521 255 19579 261
rect 19521 252 19533 255
rect 19200 224 19533 252
rect 19200 221 19212 224
rect 19154 215 19212 221
rect 19521 221 19533 224
rect 19567 252 19579 255
rect 20237 255 20295 261
rect 20237 252 20249 255
rect 19567 224 20249 252
rect 19567 221 19579 224
rect 19521 215 19579 221
rect 20237 221 20249 224
rect 20283 221 20295 255
rect 20237 215 20295 221
rect 20453 250 20477 294
rect 20453 216 20465 250
rect 20529 242 20573 294
rect 20499 216 20573 242
rect 18337 184 18409 187
rect 17795 156 18409 184
rect 17795 153 17807 156
rect 17677 147 17807 153
rect 18397 153 18409 156
rect 18443 184 18457 187
rect 18443 153 18455 184
rect 18397 147 18455 153
rect 19293 183 19462 191
rect 17177 122 17346 131
rect 19293 131 19344 183
rect 19396 131 19462 183
rect 19793 187 19923 193
rect 19793 153 19805 187
rect 19839 153 19877 187
rect 19911 184 19923 187
rect 20453 187 20573 216
rect 21089 282 21182 309
rect 21089 230 21113 282
rect 21165 230 21182 282
rect 22569 294 22689 300
rect 21089 208 21182 230
rect 21270 255 21328 261
rect 21270 221 21282 255
rect 21316 252 21328 255
rect 21637 255 21695 261
rect 21637 252 21649 255
rect 21316 224 21649 252
rect 21316 221 21328 224
rect 21270 215 21328 221
rect 21637 221 21649 224
rect 21683 252 21695 255
rect 22353 255 22411 261
rect 22353 252 22365 255
rect 21683 224 22365 252
rect 21683 221 21695 224
rect 21637 215 21695 221
rect 22353 221 22365 224
rect 22399 221 22411 255
rect 22353 215 22411 221
rect 22569 250 22593 294
rect 22569 216 22581 250
rect 22645 242 22689 294
rect 22615 216 22689 242
rect 20453 184 20525 187
rect 19911 156 20525 184
rect 19911 153 19923 156
rect 19793 147 19923 153
rect 20513 153 20525 156
rect 20559 184 20573 187
rect 20559 153 20571 184
rect 20513 147 20571 153
rect 21409 183 21578 191
rect 19293 122 19462 131
rect 21409 131 21460 183
rect 21512 131 21578 183
rect 21909 187 22039 193
rect 21909 153 21921 187
rect 21955 153 21993 187
rect 22027 184 22039 187
rect 22569 187 22689 216
rect 23205 282 23298 309
rect 23205 230 23229 282
rect 23281 230 23298 282
rect 24685 294 24805 300
rect 23205 208 23298 230
rect 23386 255 23444 261
rect 23386 221 23398 255
rect 23432 252 23444 255
rect 23753 255 23811 261
rect 23753 252 23765 255
rect 23432 224 23765 252
rect 23432 221 23444 224
rect 23386 215 23444 221
rect 23753 221 23765 224
rect 23799 252 23811 255
rect 24469 255 24527 261
rect 24469 252 24481 255
rect 23799 224 24481 252
rect 23799 221 23811 224
rect 23753 215 23811 221
rect 24469 221 24481 224
rect 24515 221 24527 255
rect 24469 215 24527 221
rect 24685 250 24709 294
rect 24685 216 24697 250
rect 24761 242 24805 294
rect 24731 216 24805 242
rect 22569 184 22641 187
rect 22027 156 22641 184
rect 22027 153 22039 156
rect 21909 147 22039 153
rect 22629 153 22641 156
rect 22675 184 22689 187
rect 22675 153 22687 184
rect 22629 147 22687 153
rect 23525 183 23694 191
rect 21409 122 21578 131
rect 23525 131 23576 183
rect 23628 131 23694 183
rect 24025 187 24155 193
rect 24025 153 24037 187
rect 24071 153 24109 187
rect 24143 184 24155 187
rect 24685 187 24805 216
rect 25321 282 25414 309
rect 25321 230 25345 282
rect 25397 230 25414 282
rect 26801 294 26921 300
rect 25321 208 25414 230
rect 25502 255 25560 261
rect 25502 221 25514 255
rect 25548 252 25560 255
rect 25869 255 25927 261
rect 25869 252 25881 255
rect 25548 224 25881 252
rect 25548 221 25560 224
rect 25502 215 25560 221
rect 25869 221 25881 224
rect 25915 252 25927 255
rect 26585 255 26643 261
rect 26585 252 26597 255
rect 25915 224 26597 252
rect 25915 221 25927 224
rect 25869 215 25927 221
rect 26585 221 26597 224
rect 26631 221 26643 255
rect 26585 215 26643 221
rect 26801 250 26825 294
rect 26801 216 26813 250
rect 26877 242 26921 294
rect 26847 216 26921 242
rect 24685 184 24757 187
rect 24143 156 24757 184
rect 24143 153 24155 156
rect 24025 147 24155 153
rect 24745 153 24757 156
rect 24791 184 24805 187
rect 24791 153 24803 184
rect 24745 147 24803 153
rect 25641 183 25810 191
rect 23525 122 23694 131
rect 25641 131 25692 183
rect 25744 131 25810 183
rect 26141 187 26271 193
rect 26141 153 26153 187
rect 26187 153 26225 187
rect 26259 184 26271 187
rect 26801 187 26921 216
rect 27437 282 27530 309
rect 27437 230 27461 282
rect 27513 230 27530 282
rect 28917 294 29037 300
rect 27437 208 27530 230
rect 27618 255 27676 261
rect 27618 221 27630 255
rect 27664 252 27676 255
rect 27985 255 28043 261
rect 27985 252 27997 255
rect 27664 224 27997 252
rect 27664 221 27676 224
rect 27618 215 27676 221
rect 27985 221 27997 224
rect 28031 252 28043 255
rect 28701 255 28759 261
rect 28701 252 28713 255
rect 28031 224 28713 252
rect 28031 221 28043 224
rect 27985 215 28043 221
rect 28701 221 28713 224
rect 28747 221 28759 255
rect 28701 215 28759 221
rect 28917 250 28941 294
rect 28917 216 28929 250
rect 28993 242 29037 294
rect 28963 216 29037 242
rect 26801 184 26873 187
rect 26259 156 26873 184
rect 26259 153 26271 156
rect 26141 147 26271 153
rect 26861 153 26873 156
rect 26907 184 26921 187
rect 26907 153 26919 184
rect 26861 147 26919 153
rect 27757 183 27926 191
rect 25641 122 25810 131
rect 27757 131 27808 183
rect 27860 131 27926 183
rect 28257 187 28387 193
rect 28257 153 28269 187
rect 28303 153 28341 187
rect 28375 184 28387 187
rect 28917 187 29037 216
rect 29553 282 29646 309
rect 29553 230 29577 282
rect 29629 230 29646 282
rect 31033 294 31153 300
rect 29553 208 29646 230
rect 29734 255 29792 261
rect 29734 221 29746 255
rect 29780 252 29792 255
rect 30101 255 30159 261
rect 30101 252 30113 255
rect 29780 224 30113 252
rect 29780 221 29792 224
rect 29734 215 29792 221
rect 30101 221 30113 224
rect 30147 252 30159 255
rect 30817 255 30875 261
rect 30817 252 30829 255
rect 30147 224 30829 252
rect 30147 221 30159 224
rect 30101 215 30159 221
rect 30817 221 30829 224
rect 30863 221 30875 255
rect 30817 215 30875 221
rect 31033 250 31057 294
rect 31033 216 31045 250
rect 31109 242 31153 294
rect 31079 216 31153 242
rect 28917 184 28989 187
rect 28375 156 28989 184
rect 28375 153 28387 156
rect 28257 147 28387 153
rect 28977 153 28989 156
rect 29023 184 29037 187
rect 29023 153 29035 184
rect 28977 147 29035 153
rect 29873 183 30042 191
rect 27757 122 27926 131
rect 29873 131 29924 183
rect 29976 131 30042 183
rect 30373 187 30503 193
rect 30373 153 30385 187
rect 30419 153 30457 187
rect 30491 184 30503 187
rect 31033 187 31153 216
rect 31669 282 31762 309
rect 31669 230 31693 282
rect 31745 230 31762 282
rect 33149 294 33269 300
rect 31669 208 31762 230
rect 31850 255 31908 261
rect 31850 221 31862 255
rect 31896 252 31908 255
rect 32217 255 32275 261
rect 32217 252 32229 255
rect 31896 224 32229 252
rect 31896 221 31908 224
rect 31850 215 31908 221
rect 32217 221 32229 224
rect 32263 252 32275 255
rect 32933 255 32991 261
rect 32933 252 32945 255
rect 32263 224 32945 252
rect 32263 221 32275 224
rect 32217 215 32275 221
rect 32933 221 32945 224
rect 32979 221 32991 255
rect 32933 215 32991 221
rect 33149 250 33173 294
rect 33149 216 33161 250
rect 33225 242 33269 294
rect 33195 216 33269 242
rect 31033 184 31105 187
rect 30491 156 31105 184
rect 30491 153 30503 156
rect 30373 147 30503 153
rect 31093 153 31105 156
rect 31139 184 31153 187
rect 31139 153 31151 184
rect 31093 147 31151 153
rect 31989 183 32158 191
rect 29873 122 30042 131
rect 31989 131 32040 183
rect 32092 131 32158 183
rect 32489 187 32619 193
rect 32489 153 32501 187
rect 32535 153 32573 187
rect 32607 184 32619 187
rect 33149 187 33269 216
rect 33785 282 33878 309
rect 33785 230 33809 282
rect 33861 230 33878 282
rect 35265 294 35385 300
rect 33785 208 33878 230
rect 33966 255 34024 261
rect 33966 221 33978 255
rect 34012 252 34024 255
rect 34333 255 34391 261
rect 34333 252 34345 255
rect 34012 224 34345 252
rect 34012 221 34024 224
rect 33966 215 34024 221
rect 34333 221 34345 224
rect 34379 252 34391 255
rect 35049 255 35107 261
rect 35049 252 35061 255
rect 34379 224 35061 252
rect 34379 221 34391 224
rect 34333 215 34391 221
rect 35049 221 35061 224
rect 35095 221 35107 255
rect 35049 215 35107 221
rect 35265 250 35289 294
rect 35265 216 35277 250
rect 35341 242 35385 294
rect 35311 216 35385 242
rect 33149 184 33221 187
rect 32607 156 33221 184
rect 32607 153 32619 156
rect 32489 147 32619 153
rect 33209 153 33221 156
rect 33255 184 33269 187
rect 33255 153 33267 184
rect 33209 147 33267 153
rect 34105 183 34274 191
rect 31989 122 32158 131
rect 34105 131 34156 183
rect 34208 131 34274 183
rect 34605 187 34735 193
rect 34605 153 34617 187
rect 34651 153 34689 187
rect 34723 184 34735 187
rect 35265 187 35385 216
rect 35901 282 35994 309
rect 35901 230 35925 282
rect 35977 230 35994 282
rect 37381 294 37501 300
rect 35901 208 35994 230
rect 36082 255 36140 261
rect 36082 221 36094 255
rect 36128 252 36140 255
rect 36449 255 36507 261
rect 36449 252 36461 255
rect 36128 224 36461 252
rect 36128 221 36140 224
rect 36082 215 36140 221
rect 36449 221 36461 224
rect 36495 252 36507 255
rect 37165 255 37223 261
rect 37165 252 37177 255
rect 36495 224 37177 252
rect 36495 221 36507 224
rect 36449 215 36507 221
rect 37165 221 37177 224
rect 37211 221 37223 255
rect 37165 215 37223 221
rect 37381 250 37405 294
rect 37381 216 37393 250
rect 37457 242 37501 294
rect 37427 216 37501 242
rect 35265 184 35337 187
rect 34723 156 35337 184
rect 34723 153 34735 156
rect 34605 147 34735 153
rect 35325 153 35337 156
rect 35371 184 35385 187
rect 35371 153 35383 184
rect 35325 147 35383 153
rect 36221 183 36390 191
rect 34105 122 34274 131
rect 36221 131 36272 183
rect 36324 131 36390 183
rect 36721 187 36851 193
rect 36721 153 36733 187
rect 36767 153 36805 187
rect 36839 184 36851 187
rect 37381 187 37501 216
rect 38017 282 38110 309
rect 38017 230 38041 282
rect 38093 230 38110 282
rect 39497 294 39617 300
rect 38017 208 38110 230
rect 38198 255 38256 261
rect 38198 221 38210 255
rect 38244 252 38256 255
rect 38565 255 38623 261
rect 38565 252 38577 255
rect 38244 224 38577 252
rect 38244 221 38256 224
rect 38198 215 38256 221
rect 38565 221 38577 224
rect 38611 252 38623 255
rect 39281 255 39339 261
rect 39281 252 39293 255
rect 38611 224 39293 252
rect 38611 221 38623 224
rect 38565 215 38623 221
rect 39281 221 39293 224
rect 39327 221 39339 255
rect 39281 215 39339 221
rect 39497 250 39521 294
rect 39497 216 39509 250
rect 39573 242 39617 294
rect 39543 216 39617 242
rect 37381 184 37453 187
rect 36839 156 37453 184
rect 36839 153 36851 156
rect 36721 147 36851 153
rect 37441 153 37453 156
rect 37487 184 37501 187
rect 37487 153 37499 184
rect 37441 147 37499 153
rect 38337 183 38506 191
rect 36221 122 36390 131
rect 38337 131 38388 183
rect 38440 131 38506 183
rect 38837 187 38967 193
rect 38837 153 38849 187
rect 38883 153 38921 187
rect 38955 184 38967 187
rect 39497 187 39617 216
rect 40133 282 40226 309
rect 40133 230 40157 282
rect 40209 230 40226 282
rect 41613 294 41733 300
rect 40133 208 40226 230
rect 40314 255 40372 261
rect 40314 221 40326 255
rect 40360 252 40372 255
rect 40681 255 40739 261
rect 40681 252 40693 255
rect 40360 224 40693 252
rect 40360 221 40372 224
rect 40314 215 40372 221
rect 40681 221 40693 224
rect 40727 252 40739 255
rect 41397 255 41455 261
rect 41397 252 41409 255
rect 40727 224 41409 252
rect 40727 221 40739 224
rect 40681 215 40739 221
rect 41397 221 41409 224
rect 41443 221 41455 255
rect 41397 215 41455 221
rect 41613 250 41637 294
rect 41613 216 41625 250
rect 41689 242 41733 294
rect 41659 216 41733 242
rect 39497 184 39569 187
rect 38955 156 39569 184
rect 38955 153 38967 156
rect 38837 147 38967 153
rect 39557 153 39569 156
rect 39603 184 39617 187
rect 39603 153 39615 184
rect 39557 147 39615 153
rect 40453 183 40622 191
rect 38337 122 38506 131
rect 40453 131 40504 183
rect 40556 131 40622 183
rect 40953 187 41083 193
rect 40953 153 40965 187
rect 40999 153 41037 187
rect 41071 184 41083 187
rect 41613 187 41733 216
rect 42249 282 42342 309
rect 42249 230 42273 282
rect 42325 230 42342 282
rect 42249 208 42342 230
rect 41613 184 41685 187
rect 41071 156 41685 184
rect 41071 153 41083 156
rect 40953 147 41083 153
rect 41673 153 41685 156
rect 41719 184 41733 187
rect 41719 153 41731 184
rect 41673 147 41731 153
rect 40453 122 40622 131
rect 0 17 42320 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2697 17
rect 2731 -17 2789 17
rect 2823 -17 2881 17
rect 2915 -17 2973 17
rect 3007 -17 3065 17
rect 3099 -17 3157 17
rect 3191 -17 3249 17
rect 3283 -17 3341 17
rect 3375 -17 3433 17
rect 3467 -17 3525 17
rect 3559 -17 3617 17
rect 3651 -17 3709 17
rect 3743 -17 3801 17
rect 3835 -17 3893 17
rect 3927 -17 3985 17
rect 4019 -17 4077 17
rect 4111 -17 4169 17
rect 4203 -17 4261 17
rect 4295 -17 4353 17
rect 4387 -17 4445 17
rect 4479 -17 4537 17
rect 4571 -17 4629 17
rect 4663 -17 4721 17
rect 4755 -17 4813 17
rect 4847 -17 4905 17
rect 4939 -17 4997 17
rect 5031 -17 5089 17
rect 5123 -17 5181 17
rect 5215 -17 5273 17
rect 5307 -17 5365 17
rect 5399 -17 5457 17
rect 5491 -17 5549 17
rect 5583 -17 5641 17
rect 5675 -17 5733 17
rect 5767 -17 5825 17
rect 5859 -17 5917 17
rect 5951 -17 6009 17
rect 6043 -17 6101 17
rect 6135 -17 6193 17
rect 6227 -17 6285 17
rect 6319 -17 6377 17
rect 6411 -17 6469 17
rect 6503 -17 6561 17
rect 6595 -17 6653 17
rect 6687 -17 6745 17
rect 6779 -17 6837 17
rect 6871 -17 6929 17
rect 6963 -17 7021 17
rect 7055 -17 7113 17
rect 7147 -17 7205 17
rect 7239 -17 7297 17
rect 7331 -17 7389 17
rect 7423 -17 7481 17
rect 7515 -17 7573 17
rect 7607 -17 7665 17
rect 7699 -17 7757 17
rect 7791 -17 7849 17
rect 7883 -17 7941 17
rect 7975 -17 8033 17
rect 8067 -17 8125 17
rect 8159 -17 8217 17
rect 8251 -17 8309 17
rect 8343 -17 8401 17
rect 8435 -17 8493 17
rect 8527 -17 8585 17
rect 8619 -17 8677 17
rect 8711 -17 8769 17
rect 8803 -17 8861 17
rect 8895 -17 8953 17
rect 8987 -17 9045 17
rect 9079 -17 9137 17
rect 9171 -17 9229 17
rect 9263 -17 9321 17
rect 9355 -17 9413 17
rect 9447 -17 9505 17
rect 9539 -17 9597 17
rect 9631 -17 9689 17
rect 9723 -17 9781 17
rect 9815 -17 9873 17
rect 9907 -17 9965 17
rect 9999 -17 10057 17
rect 10091 -17 10149 17
rect 10183 -17 10241 17
rect 10275 -17 10333 17
rect 10367 -17 10425 17
rect 10459 -17 10517 17
rect 10551 -17 10609 17
rect 10643 -17 10701 17
rect 10735 -17 10793 17
rect 10827 -17 10885 17
rect 10919 -17 10977 17
rect 11011 -17 11069 17
rect 11103 -17 11161 17
rect 11195 -17 11253 17
rect 11287 -17 11345 17
rect 11379 -17 11437 17
rect 11471 -17 11529 17
rect 11563 -17 11621 17
rect 11655 -17 11713 17
rect 11747 -17 11805 17
rect 11839 -17 11897 17
rect 11931 -17 11989 17
rect 12023 -17 12081 17
rect 12115 -17 12173 17
rect 12207 -17 12265 17
rect 12299 -17 12357 17
rect 12391 -17 12449 17
rect 12483 -17 12541 17
rect 12575 -17 12633 17
rect 12667 -17 12725 17
rect 12759 -17 12817 17
rect 12851 -17 12909 17
rect 12943 -17 13001 17
rect 13035 -17 13093 17
rect 13127 -17 13185 17
rect 13219 -17 13277 17
rect 13311 -17 13369 17
rect 13403 -17 13461 17
rect 13495 -17 13553 17
rect 13587 -17 13645 17
rect 13679 -17 13737 17
rect 13771 -17 13829 17
rect 13863 -17 13921 17
rect 13955 -17 14013 17
rect 14047 -17 14105 17
rect 14139 -17 14197 17
rect 14231 -17 14289 17
rect 14323 -17 14381 17
rect 14415 -17 14473 17
rect 14507 -17 14565 17
rect 14599 -17 14657 17
rect 14691 -17 14749 17
rect 14783 -17 14841 17
rect 14875 -17 14933 17
rect 14967 -17 15025 17
rect 15059 -17 15117 17
rect 15151 -17 15209 17
rect 15243 -17 15301 17
rect 15335 -17 15393 17
rect 15427 -17 15485 17
rect 15519 -17 15577 17
rect 15611 -17 15669 17
rect 15703 -17 15761 17
rect 15795 -17 15853 17
rect 15887 -17 15945 17
rect 15979 -17 16037 17
rect 16071 -17 16129 17
rect 16163 -17 16221 17
rect 16255 -17 16313 17
rect 16347 -17 16405 17
rect 16439 -17 16497 17
rect 16531 -17 16589 17
rect 16623 -17 16681 17
rect 16715 -17 16773 17
rect 16807 -17 16865 17
rect 16899 -17 16957 17
rect 16991 -17 17049 17
rect 17083 -17 17141 17
rect 17175 -17 17233 17
rect 17267 -17 17325 17
rect 17359 -17 17417 17
rect 17451 -17 17509 17
rect 17543 -17 17601 17
rect 17635 -17 17693 17
rect 17727 -17 17785 17
rect 17819 -17 17877 17
rect 17911 -17 17969 17
rect 18003 -17 18061 17
rect 18095 -17 18153 17
rect 18187 -17 18245 17
rect 18279 -17 18337 17
rect 18371 -17 18429 17
rect 18463 -17 18521 17
rect 18555 -17 18613 17
rect 18647 -17 18705 17
rect 18739 -17 18797 17
rect 18831 -17 18889 17
rect 18923 -17 18981 17
rect 19015 -17 19073 17
rect 19107 -17 19165 17
rect 19199 -17 19257 17
rect 19291 -17 19349 17
rect 19383 -17 19441 17
rect 19475 -17 19533 17
rect 19567 -17 19625 17
rect 19659 -17 19717 17
rect 19751 -17 19809 17
rect 19843 -17 19901 17
rect 19935 -17 19993 17
rect 20027 -17 20085 17
rect 20119 -17 20177 17
rect 20211 -17 20269 17
rect 20303 -17 20361 17
rect 20395 -17 20453 17
rect 20487 -17 20545 17
rect 20579 -17 20637 17
rect 20671 -17 20729 17
rect 20763 -17 20821 17
rect 20855 -17 20913 17
rect 20947 -17 21005 17
rect 21039 -17 21097 17
rect 21131 -17 21189 17
rect 21223 -17 21281 17
rect 21315 -17 21373 17
rect 21407 -17 21465 17
rect 21499 -17 21557 17
rect 21591 -17 21649 17
rect 21683 -17 21741 17
rect 21775 -17 21833 17
rect 21867 -17 21925 17
rect 21959 -17 22017 17
rect 22051 -17 22109 17
rect 22143 -17 22201 17
rect 22235 -17 22293 17
rect 22327 -17 22385 17
rect 22419 -17 22477 17
rect 22511 -17 22569 17
rect 22603 -17 22661 17
rect 22695 -17 22753 17
rect 22787 -17 22845 17
rect 22879 -17 22937 17
rect 22971 -17 23029 17
rect 23063 -17 23121 17
rect 23155 -17 23213 17
rect 23247 -17 23305 17
rect 23339 -17 23397 17
rect 23431 -17 23489 17
rect 23523 -17 23581 17
rect 23615 -17 23673 17
rect 23707 -17 23765 17
rect 23799 -17 23857 17
rect 23891 -17 23949 17
rect 23983 -17 24041 17
rect 24075 -17 24133 17
rect 24167 -17 24225 17
rect 24259 -17 24317 17
rect 24351 -17 24409 17
rect 24443 -17 24501 17
rect 24535 -17 24593 17
rect 24627 -17 24685 17
rect 24719 -17 24777 17
rect 24811 -17 24869 17
rect 24903 -17 24961 17
rect 24995 -17 25053 17
rect 25087 -17 25145 17
rect 25179 -17 25237 17
rect 25271 -17 25329 17
rect 25363 -17 25421 17
rect 25455 -17 25513 17
rect 25547 -17 25605 17
rect 25639 -17 25697 17
rect 25731 -17 25789 17
rect 25823 -17 25881 17
rect 25915 -17 25973 17
rect 26007 -17 26065 17
rect 26099 -17 26157 17
rect 26191 -17 26249 17
rect 26283 -17 26341 17
rect 26375 -17 26433 17
rect 26467 -17 26525 17
rect 26559 -17 26617 17
rect 26651 -17 26709 17
rect 26743 -17 26801 17
rect 26835 -17 26893 17
rect 26927 -17 26985 17
rect 27019 -17 27077 17
rect 27111 -17 27169 17
rect 27203 -17 27261 17
rect 27295 -17 27353 17
rect 27387 -17 27445 17
rect 27479 -17 27537 17
rect 27571 -17 27629 17
rect 27663 -17 27721 17
rect 27755 -17 27813 17
rect 27847 -17 27905 17
rect 27939 -17 27997 17
rect 28031 -17 28089 17
rect 28123 -17 28181 17
rect 28215 -17 28273 17
rect 28307 -17 28365 17
rect 28399 -17 28457 17
rect 28491 -17 28549 17
rect 28583 -17 28641 17
rect 28675 -17 28733 17
rect 28767 -17 28825 17
rect 28859 -17 28917 17
rect 28951 -17 29009 17
rect 29043 -17 29101 17
rect 29135 -17 29193 17
rect 29227 -17 29285 17
rect 29319 -17 29377 17
rect 29411 -17 29469 17
rect 29503 -17 29561 17
rect 29595 -17 29653 17
rect 29687 -17 29745 17
rect 29779 -17 29837 17
rect 29871 -17 29929 17
rect 29963 -17 30021 17
rect 30055 -17 30113 17
rect 30147 -17 30205 17
rect 30239 -17 30297 17
rect 30331 -17 30389 17
rect 30423 -17 30481 17
rect 30515 -17 30573 17
rect 30607 -17 30665 17
rect 30699 -17 30757 17
rect 30791 -17 30849 17
rect 30883 -17 30941 17
rect 30975 -17 31033 17
rect 31067 -17 31125 17
rect 31159 -17 31217 17
rect 31251 -17 31309 17
rect 31343 -17 31401 17
rect 31435 -17 31493 17
rect 31527 -17 31585 17
rect 31619 -17 31677 17
rect 31711 -17 31769 17
rect 31803 -17 31861 17
rect 31895 -17 31953 17
rect 31987 -17 32045 17
rect 32079 -17 32137 17
rect 32171 -17 32229 17
rect 32263 -17 32321 17
rect 32355 -17 32413 17
rect 32447 -17 32505 17
rect 32539 -17 32597 17
rect 32631 -17 32689 17
rect 32723 -17 32781 17
rect 32815 -17 32873 17
rect 32907 -17 32965 17
rect 32999 -17 33057 17
rect 33091 -17 33149 17
rect 33183 -17 33241 17
rect 33275 -17 33333 17
rect 33367 -17 33425 17
rect 33459 -17 33517 17
rect 33551 -17 33609 17
rect 33643 -17 33701 17
rect 33735 -17 33793 17
rect 33827 -17 33885 17
rect 33919 -17 33977 17
rect 34011 -17 34069 17
rect 34103 -17 34161 17
rect 34195 -17 34253 17
rect 34287 -17 34345 17
rect 34379 -17 34437 17
rect 34471 -17 34529 17
rect 34563 -17 34621 17
rect 34655 -17 34713 17
rect 34747 -17 34805 17
rect 34839 -17 34897 17
rect 34931 -17 34989 17
rect 35023 -17 35081 17
rect 35115 -17 35173 17
rect 35207 -17 35265 17
rect 35299 -17 35357 17
rect 35391 -17 35449 17
rect 35483 -17 35541 17
rect 35575 -17 35633 17
rect 35667 -17 35725 17
rect 35759 -17 35817 17
rect 35851 -17 35909 17
rect 35943 -17 36001 17
rect 36035 -17 36093 17
rect 36127 -17 36185 17
rect 36219 -17 36277 17
rect 36311 -17 36369 17
rect 36403 -17 36461 17
rect 36495 -17 36553 17
rect 36587 -17 36645 17
rect 36679 -17 36737 17
rect 36771 -17 36829 17
rect 36863 -17 36921 17
rect 36955 -17 37013 17
rect 37047 -17 37105 17
rect 37139 -17 37197 17
rect 37231 -17 37289 17
rect 37323 -17 37381 17
rect 37415 -17 37473 17
rect 37507 -17 37565 17
rect 37599 -17 37657 17
rect 37691 -17 37749 17
rect 37783 -17 37841 17
rect 37875 -17 37933 17
rect 37967 -17 38025 17
rect 38059 -17 38117 17
rect 38151 -17 38209 17
rect 38243 -17 38301 17
rect 38335 -17 38393 17
rect 38427 -17 38485 17
rect 38519 -17 38577 17
rect 38611 -17 38669 17
rect 38703 -17 38761 17
rect 38795 -17 38853 17
rect 38887 -17 38945 17
rect 38979 -17 39037 17
rect 39071 -17 39129 17
rect 39163 -17 39221 17
rect 39255 -17 39313 17
rect 39347 -17 39405 17
rect 39439 -17 39497 17
rect 39531 -17 39589 17
rect 39623 -17 39681 17
rect 39715 -17 39773 17
rect 39807 -17 39865 17
rect 39899 -17 39957 17
rect 39991 -17 40049 17
rect 40083 -17 40141 17
rect 40175 -17 40233 17
rect 40267 -17 40325 17
rect 40359 -17 40417 17
rect 40451 -17 40509 17
rect 40543 -17 40601 17
rect 40635 -17 40693 17
rect 40727 -17 40785 17
rect 40819 -17 40877 17
rect 40911 -17 40969 17
rect 41003 -17 41061 17
rect 41095 -17 41153 17
rect 41187 -17 41245 17
rect 41279 -17 41337 17
rect 41371 -17 41429 17
rect 41463 -17 41521 17
rect 41555 -17 41613 17
rect 41647 -17 41705 17
rect 41739 -17 41797 17
rect 41831 -17 41889 17
rect 41923 -17 41981 17
rect 42015 -17 42073 17
rect 42107 -17 42165 17
rect 42199 -17 42257 17
rect 42291 -17 42320 17
rect 0 -48 42320 -17
<< via1 >>
rect 1433 250 1485 294
rect 1433 242 1455 250
rect 1455 242 1485 250
rect 300 175 352 183
rect 300 141 307 175
rect 307 141 345 175
rect 345 141 352 175
rect 300 131 352 141
rect 2069 274 2121 282
rect 2069 240 2076 274
rect 2076 240 2114 274
rect 2114 240 2121 274
rect 2069 230 2121 240
rect 3549 250 3601 294
rect 3549 242 3571 250
rect 3571 242 3601 250
rect 2416 175 2468 183
rect 2416 141 2423 175
rect 2423 141 2461 175
rect 2461 141 2468 175
rect 2416 131 2468 141
rect 4185 274 4237 282
rect 4185 240 4192 274
rect 4192 240 4230 274
rect 4230 240 4237 274
rect 4185 230 4237 240
rect 5665 250 5717 294
rect 5665 242 5687 250
rect 5687 242 5717 250
rect 4532 175 4584 183
rect 4532 141 4539 175
rect 4539 141 4577 175
rect 4577 141 4584 175
rect 4532 131 4584 141
rect 6301 274 6353 282
rect 6301 240 6308 274
rect 6308 240 6346 274
rect 6346 240 6353 274
rect 6301 230 6353 240
rect 7781 250 7833 294
rect 7781 242 7803 250
rect 7803 242 7833 250
rect 6648 175 6700 183
rect 6648 141 6655 175
rect 6655 141 6693 175
rect 6693 141 6700 175
rect 6648 131 6700 141
rect 8417 274 8469 282
rect 8417 240 8424 274
rect 8424 240 8462 274
rect 8462 240 8469 274
rect 8417 230 8469 240
rect 9897 250 9949 294
rect 9897 242 9919 250
rect 9919 242 9949 250
rect 8764 175 8816 183
rect 8764 141 8771 175
rect 8771 141 8809 175
rect 8809 141 8816 175
rect 8764 131 8816 141
rect 10533 274 10585 282
rect 10533 240 10540 274
rect 10540 240 10578 274
rect 10578 240 10585 274
rect 10533 230 10585 240
rect 12013 250 12065 294
rect 12013 242 12035 250
rect 12035 242 12065 250
rect 10880 175 10932 183
rect 10880 141 10887 175
rect 10887 141 10925 175
rect 10925 141 10932 175
rect 10880 131 10932 141
rect 12649 274 12701 282
rect 12649 240 12656 274
rect 12656 240 12694 274
rect 12694 240 12701 274
rect 12649 230 12701 240
rect 14129 250 14181 294
rect 14129 242 14151 250
rect 14151 242 14181 250
rect 12996 175 13048 183
rect 12996 141 13003 175
rect 13003 141 13041 175
rect 13041 141 13048 175
rect 12996 131 13048 141
rect 14765 274 14817 282
rect 14765 240 14772 274
rect 14772 240 14810 274
rect 14810 240 14817 274
rect 14765 230 14817 240
rect 16245 250 16297 294
rect 16245 242 16267 250
rect 16267 242 16297 250
rect 15112 175 15164 183
rect 15112 141 15119 175
rect 15119 141 15157 175
rect 15157 141 15164 175
rect 15112 131 15164 141
rect 16881 274 16933 282
rect 16881 240 16888 274
rect 16888 240 16926 274
rect 16926 240 16933 274
rect 16881 230 16933 240
rect 18361 250 18413 294
rect 18361 242 18383 250
rect 18383 242 18413 250
rect 17228 175 17280 183
rect 17228 141 17235 175
rect 17235 141 17273 175
rect 17273 141 17280 175
rect 17228 131 17280 141
rect 18997 274 19049 282
rect 18997 240 19004 274
rect 19004 240 19042 274
rect 19042 240 19049 274
rect 18997 230 19049 240
rect 20477 250 20529 294
rect 20477 242 20499 250
rect 20499 242 20529 250
rect 19344 175 19396 183
rect 19344 141 19351 175
rect 19351 141 19389 175
rect 19389 141 19396 175
rect 19344 131 19396 141
rect 21113 274 21165 282
rect 21113 240 21120 274
rect 21120 240 21158 274
rect 21158 240 21165 274
rect 21113 230 21165 240
rect 22593 250 22645 294
rect 22593 242 22615 250
rect 22615 242 22645 250
rect 21460 175 21512 183
rect 21460 141 21467 175
rect 21467 141 21505 175
rect 21505 141 21512 175
rect 21460 131 21512 141
rect 23229 274 23281 282
rect 23229 240 23236 274
rect 23236 240 23274 274
rect 23274 240 23281 274
rect 23229 230 23281 240
rect 24709 250 24761 294
rect 24709 242 24731 250
rect 24731 242 24761 250
rect 23576 175 23628 183
rect 23576 141 23583 175
rect 23583 141 23621 175
rect 23621 141 23628 175
rect 23576 131 23628 141
rect 25345 274 25397 282
rect 25345 240 25352 274
rect 25352 240 25390 274
rect 25390 240 25397 274
rect 25345 230 25397 240
rect 26825 250 26877 294
rect 26825 242 26847 250
rect 26847 242 26877 250
rect 25692 175 25744 183
rect 25692 141 25699 175
rect 25699 141 25737 175
rect 25737 141 25744 175
rect 25692 131 25744 141
rect 27461 274 27513 282
rect 27461 240 27468 274
rect 27468 240 27506 274
rect 27506 240 27513 274
rect 27461 230 27513 240
rect 28941 250 28993 294
rect 28941 242 28963 250
rect 28963 242 28993 250
rect 27808 175 27860 183
rect 27808 141 27815 175
rect 27815 141 27853 175
rect 27853 141 27860 175
rect 27808 131 27860 141
rect 29577 274 29629 282
rect 29577 240 29584 274
rect 29584 240 29622 274
rect 29622 240 29629 274
rect 29577 230 29629 240
rect 31057 250 31109 294
rect 31057 242 31079 250
rect 31079 242 31109 250
rect 29924 175 29976 183
rect 29924 141 29931 175
rect 29931 141 29969 175
rect 29969 141 29976 175
rect 29924 131 29976 141
rect 31693 274 31745 282
rect 31693 240 31700 274
rect 31700 240 31738 274
rect 31738 240 31745 274
rect 31693 230 31745 240
rect 33173 250 33225 294
rect 33173 242 33195 250
rect 33195 242 33225 250
rect 32040 175 32092 183
rect 32040 141 32047 175
rect 32047 141 32085 175
rect 32085 141 32092 175
rect 32040 131 32092 141
rect 33809 274 33861 282
rect 33809 240 33816 274
rect 33816 240 33854 274
rect 33854 240 33861 274
rect 33809 230 33861 240
rect 35289 250 35341 294
rect 35289 242 35311 250
rect 35311 242 35341 250
rect 34156 175 34208 183
rect 34156 141 34163 175
rect 34163 141 34201 175
rect 34201 141 34208 175
rect 34156 131 34208 141
rect 35925 274 35977 282
rect 35925 240 35932 274
rect 35932 240 35970 274
rect 35970 240 35977 274
rect 35925 230 35977 240
rect 37405 250 37457 294
rect 37405 242 37427 250
rect 37427 242 37457 250
rect 36272 175 36324 183
rect 36272 141 36279 175
rect 36279 141 36317 175
rect 36317 141 36324 175
rect 36272 131 36324 141
rect 38041 274 38093 282
rect 38041 240 38048 274
rect 38048 240 38086 274
rect 38086 240 38093 274
rect 38041 230 38093 240
rect 39521 250 39573 294
rect 39521 242 39543 250
rect 39543 242 39573 250
rect 38388 175 38440 183
rect 38388 141 38395 175
rect 38395 141 38433 175
rect 38433 141 38440 175
rect 38388 131 38440 141
rect 40157 274 40209 282
rect 40157 240 40164 274
rect 40164 240 40202 274
rect 40202 240 40209 274
rect 40157 230 40209 240
rect 41637 250 41689 294
rect 41637 242 41659 250
rect 41659 242 41689 250
rect 40504 175 40556 183
rect 40504 141 40511 175
rect 40511 141 40549 175
rect 40549 141 40556 175
rect 40504 131 40556 141
rect 42273 274 42325 282
rect 42273 240 42280 274
rect 42280 240 42318 274
rect 42318 240 42325 274
rect 42273 230 42325 240
<< metal2 >>
rect 1409 357 41733 426
rect 1409 294 1529 357
rect 1409 242 1433 294
rect 1485 242 1529 294
rect 1409 220 1529 242
rect 2045 282 2138 325
rect 2045 230 2069 282
rect 2121 230 2138 282
rect 2045 191 2138 230
rect 3525 294 3645 357
rect 3525 242 3549 294
rect 3601 242 3645 294
rect 3525 220 3645 242
rect 4161 282 4254 325
rect 4161 230 4185 282
rect 4237 230 4254 282
rect 4161 191 4254 230
rect 5641 294 5761 357
rect 5641 242 5665 294
rect 5717 242 5761 294
rect 5641 220 5761 242
rect 6277 282 6370 325
rect 6277 230 6301 282
rect 6353 230 6370 282
rect 6277 191 6370 230
rect 7757 294 7877 357
rect 7757 242 7781 294
rect 7833 242 7877 294
rect 7757 220 7877 242
rect 8393 282 8486 325
rect 8393 230 8417 282
rect 8469 230 8486 282
rect 8393 191 8486 230
rect 9873 294 9993 357
rect 9873 242 9897 294
rect 9949 242 9993 294
rect 9873 220 9993 242
rect 10509 282 10602 325
rect 10509 230 10533 282
rect 10585 230 10602 282
rect 10509 191 10602 230
rect 11989 294 12109 357
rect 11989 242 12013 294
rect 12065 242 12109 294
rect 11989 220 12109 242
rect 12625 282 12718 325
rect 12625 230 12649 282
rect 12701 230 12718 282
rect 12625 191 12718 230
rect 14105 294 14225 357
rect 14105 242 14129 294
rect 14181 242 14225 294
rect 14105 220 14225 242
rect 14741 282 14834 325
rect 14741 230 14765 282
rect 14817 230 14834 282
rect 14741 191 14834 230
rect 16221 294 16341 357
rect 16221 242 16245 294
rect 16297 242 16341 294
rect 16221 220 16341 242
rect 16857 282 16950 325
rect 16857 230 16881 282
rect 16933 230 16950 282
rect 16857 191 16950 230
rect 18337 294 18457 357
rect 18337 242 18361 294
rect 18413 242 18457 294
rect 18337 220 18457 242
rect 18973 282 19066 325
rect 18973 230 18997 282
rect 19049 230 19066 282
rect 18973 191 19066 230
rect 20453 294 20573 357
rect 20453 242 20477 294
rect 20529 242 20573 294
rect 20453 220 20573 242
rect 21089 282 21182 325
rect 21089 230 21113 282
rect 21165 230 21182 282
rect 21089 191 21182 230
rect 22569 294 22689 357
rect 22569 242 22593 294
rect 22645 242 22689 294
rect 22569 220 22689 242
rect 23205 282 23298 325
rect 23205 230 23229 282
rect 23281 230 23298 282
rect 23205 191 23298 230
rect 24685 294 24805 357
rect 24685 242 24709 294
rect 24761 242 24805 294
rect 24685 220 24805 242
rect 25321 282 25414 325
rect 25321 230 25345 282
rect 25397 230 25414 282
rect 25321 191 25414 230
rect 26801 294 26921 357
rect 26801 242 26825 294
rect 26877 242 26921 294
rect 26801 220 26921 242
rect 27437 282 27530 325
rect 27437 230 27461 282
rect 27513 230 27530 282
rect 27437 191 27530 230
rect 28917 294 29037 357
rect 28917 242 28941 294
rect 28993 242 29037 294
rect 28917 220 29037 242
rect 29553 282 29646 325
rect 29553 230 29577 282
rect 29629 230 29646 282
rect 29553 191 29646 230
rect 31033 294 31153 357
rect 31033 242 31057 294
rect 31109 242 31153 294
rect 31033 220 31153 242
rect 31669 282 31762 325
rect 31669 230 31693 282
rect 31745 230 31762 282
rect 31669 191 31762 230
rect 33149 294 33269 357
rect 33149 242 33173 294
rect 33225 242 33269 294
rect 33149 220 33269 242
rect 33785 282 33878 325
rect 33785 230 33809 282
rect 33861 230 33878 282
rect 33785 191 33878 230
rect 35265 294 35385 357
rect 35265 242 35289 294
rect 35341 242 35385 294
rect 35265 220 35385 242
rect 35901 282 35994 325
rect 35901 230 35925 282
rect 35977 230 35994 282
rect 35901 191 35994 230
rect 37381 294 37501 357
rect 37381 242 37405 294
rect 37457 242 37501 294
rect 37381 220 37501 242
rect 38017 282 38110 325
rect 38017 230 38041 282
rect 38093 230 38110 282
rect 38017 191 38110 230
rect 39497 294 39617 357
rect 39497 242 39521 294
rect 39573 242 39617 294
rect 39497 220 39617 242
rect 40133 282 40226 325
rect 40133 230 40157 282
rect 40209 230 40226 282
rect 40133 191 40226 230
rect 41613 294 41733 357
rect 41613 242 41637 294
rect 41689 242 41733 294
rect 41613 220 41733 242
rect 42249 282 42342 325
rect 42249 230 42273 282
rect 42325 230 42342 282
rect 42249 191 42342 230
rect 249 183 2138 191
rect 249 131 300 183
rect 352 131 2138 183
rect 249 122 2138 131
rect 2365 183 4254 191
rect 2365 131 2416 183
rect 2468 131 4254 183
rect 2365 122 4254 131
rect 4481 183 6370 191
rect 4481 131 4532 183
rect 4584 131 6370 183
rect 4481 122 6370 131
rect 6597 183 8486 191
rect 6597 131 6648 183
rect 6700 131 8486 183
rect 6597 122 8486 131
rect 8713 183 10602 191
rect 8713 131 8764 183
rect 8816 131 10602 183
rect 8713 122 10602 131
rect 10829 183 12718 191
rect 10829 131 10880 183
rect 10932 131 12718 183
rect 10829 122 12718 131
rect 12945 183 14834 191
rect 12945 131 12996 183
rect 13048 131 14834 183
rect 12945 122 14834 131
rect 15061 183 16950 191
rect 15061 131 15112 183
rect 15164 131 16950 183
rect 15061 122 16950 131
rect 17177 183 19066 191
rect 17177 131 17228 183
rect 17280 131 19066 183
rect 17177 122 19066 131
rect 19293 183 21182 191
rect 19293 131 19344 183
rect 19396 131 21182 183
rect 19293 122 21182 131
rect 21409 183 23298 191
rect 21409 131 21460 183
rect 21512 131 23298 183
rect 21409 122 23298 131
rect 23525 183 25414 191
rect 23525 131 23576 183
rect 23628 131 25414 183
rect 23525 122 25414 131
rect 25641 183 27530 191
rect 25641 131 25692 183
rect 25744 131 27530 183
rect 25641 122 27530 131
rect 27757 183 29646 191
rect 27757 131 27808 183
rect 27860 131 29646 183
rect 27757 122 29646 131
rect 29873 183 31762 191
rect 29873 131 29924 183
rect 29976 131 31762 183
rect 29873 122 31762 131
rect 31989 183 33878 191
rect 31989 131 32040 183
rect 32092 131 33878 183
rect 31989 122 33878 131
rect 34105 183 35994 191
rect 34105 131 34156 183
rect 34208 131 35994 183
rect 34105 122 35994 131
rect 36221 183 38110 191
rect 36221 131 36272 183
rect 36324 131 38110 183
rect 36221 122 38110 131
rect 38337 183 40226 191
rect 38337 131 38388 183
rect 38440 131 40226 183
rect 38337 122 40226 131
rect 40453 183 42342 191
rect 40453 131 40504 183
rect 40556 131 42342 183
rect 40453 122 42342 131
<< labels >>
flabel locali 1481 153 1515 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
flabel locali 30 221 64 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK
rlabel viali 1481 153 1515 187 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel locali 1481 127 1529 207 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel locali 1421 207 1529 281 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 1469 147 1527 156 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 1409 193 1467 256 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 1409 184 1527 193 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 749 184 879 193 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 749 156 1527 184 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 749 147 879 156 1 sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
flabel locali 1754 218 1783 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/Q
flabel locali 2056 221 2078 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/Q_N
flabel locali 30 289 64 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK
flabel locali 305 289 339 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[0]/D
rlabel viali 29 527 63 561 3 sky130_fd_sc_hd__dfrbp_1_0[0]/VPWR
rlabel viali 121 527 155 561 3 sky130_fd_sc_hd__dfrbp_1_0[0]/VPB
rlabel viali 29 -17 63 17 3 sky130_fd_sc_hd__dfrbp_1_0[0]/VGND
rlabel viali 121 -17 155 17 3 sky130_fd_sc_hd__dfrbp_1_0[0]/VNB
flabel locali 3597 153 3631 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
flabel locali 2146 221 2180 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/CLK
rlabel viali 3597 153 3631 187 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel locali 3597 127 3645 207 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel locali 3537 207 3645 281 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 3585 147 3643 156 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 3525 193 3583 256 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 3525 184 3643 193 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 2865 184 2995 193 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 2865 156 3643 184 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 2865 147 2995 156 1 sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
flabel locali 3870 218 3899 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/Q
flabel locali 4172 221 4194 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/Q_N
flabel locali 2146 289 2180 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/CLK
flabel locali 2421 289 2455 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[1]/D
rlabel viali 2145 527 2179 561 3 sky130_fd_sc_hd__dfrbp_1_0[1]/VPWR
rlabel viali 2237 527 2271 561 3 sky130_fd_sc_hd__dfrbp_1_0[1]/VPB
rlabel viali 2145 -17 2179 17 3 sky130_fd_sc_hd__dfrbp_1_0[1]/VGND
rlabel viali 2237 -17 2271 17 3 sky130_fd_sc_hd__dfrbp_1_0[1]/VNB
flabel locali 5713 153 5747 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
flabel locali 4262 221 4296 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/CLK
rlabel viali 5713 153 5747 187 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel locali 5713 127 5761 207 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel locali 5653 207 5761 281 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 5701 147 5759 156 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 5641 193 5699 256 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 5641 184 5759 193 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 4981 184 5111 193 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 4981 156 5759 184 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 4981 147 5111 156 1 sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
flabel locali 5986 218 6015 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/Q
flabel locali 6288 221 6310 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/Q_N
flabel locali 4262 289 4296 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/CLK
flabel locali 4537 289 4571 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[2]/D
rlabel viali 4261 527 4295 561 3 sky130_fd_sc_hd__dfrbp_1_0[2]/VPWR
rlabel viali 4353 527 4387 561 3 sky130_fd_sc_hd__dfrbp_1_0[2]/VPB
rlabel viali 4261 -17 4295 17 3 sky130_fd_sc_hd__dfrbp_1_0[2]/VGND
rlabel viali 4353 -17 4387 17 3 sky130_fd_sc_hd__dfrbp_1_0[2]/VNB
flabel locali 7829 153 7863 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
flabel locali 6378 221 6412 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/CLK
rlabel viali 7829 153 7863 187 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel locali 7829 127 7877 207 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel locali 7769 207 7877 281 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7817 147 7875 156 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7757 193 7815 256 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7757 184 7875 193 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7097 184 7227 193 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7097 156 7875 184 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 7097 147 7227 156 1 sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
flabel locali 8102 218 8131 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/Q
flabel locali 8404 221 8426 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/Q_N
flabel locali 6378 289 6412 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/CLK
flabel locali 6653 289 6687 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[3]/D
rlabel viali 6377 527 6411 561 3 sky130_fd_sc_hd__dfrbp_1_0[3]/VPWR
rlabel viali 6469 527 6503 561 3 sky130_fd_sc_hd__dfrbp_1_0[3]/VPB
rlabel viali 6377 -17 6411 17 3 sky130_fd_sc_hd__dfrbp_1_0[3]/VGND
rlabel viali 6469 -17 6503 17 3 sky130_fd_sc_hd__dfrbp_1_0[3]/VNB
flabel locali 9945 153 9979 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
flabel locali 8494 221 8528 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/CLK
rlabel viali 9945 153 9979 187 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel locali 9945 127 9993 207 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel locali 9885 207 9993 281 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9933 147 9991 156 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9873 193 9931 256 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9873 184 9991 193 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9213 184 9343 193 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9213 156 9991 184 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 9213 147 9343 156 1 sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
flabel locali 10218 218 10247 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/Q
flabel locali 10520 221 10542 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/Q_N
flabel locali 8494 289 8528 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/CLK
flabel locali 8769 289 8803 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[4]/D
rlabel viali 8493 527 8527 561 3 sky130_fd_sc_hd__dfrbp_1_0[4]/VPWR
rlabel viali 8585 527 8619 561 3 sky130_fd_sc_hd__dfrbp_1_0[4]/VPB
rlabel viali 8493 -17 8527 17 3 sky130_fd_sc_hd__dfrbp_1_0[4]/VGND
rlabel viali 8585 -17 8619 17 3 sky130_fd_sc_hd__dfrbp_1_0[4]/VNB
flabel locali 12061 153 12095 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
flabel locali 10610 221 10644 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/CLK
rlabel viali 12061 153 12095 187 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel locali 12061 127 12109 207 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel locali 12001 207 12109 281 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 12049 147 12107 156 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 11989 193 12047 256 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 11989 184 12107 193 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 11329 184 11459 193 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 11329 156 12107 184 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 11329 147 11459 156 1 sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
flabel locali 12334 218 12363 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/Q
flabel locali 12636 221 12658 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/Q_N
flabel locali 10610 289 10644 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/CLK
flabel locali 10885 289 10919 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[5]/D
rlabel viali 10609 527 10643 561 3 sky130_fd_sc_hd__dfrbp_1_0[5]/VPWR
rlabel viali 10701 527 10735 561 3 sky130_fd_sc_hd__dfrbp_1_0[5]/VPB
rlabel viali 10609 -17 10643 17 3 sky130_fd_sc_hd__dfrbp_1_0[5]/VGND
rlabel viali 10701 -17 10735 17 3 sky130_fd_sc_hd__dfrbp_1_0[5]/VNB
flabel locali 14177 153 14211 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
flabel locali 12726 221 12760 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/CLK
rlabel viali 14177 153 14211 187 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel locali 14177 127 14225 207 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel locali 14117 207 14225 281 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 14165 147 14223 156 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 14105 193 14163 256 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 14105 184 14223 193 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 13445 184 13575 193 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 13445 156 14223 184 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 13445 147 13575 156 1 sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
flabel locali 14450 218 14479 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/Q
flabel locali 14752 221 14774 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/Q_N
flabel locali 12726 289 12760 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/CLK
flabel locali 13001 289 13035 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[6]/D
rlabel viali 12725 527 12759 561 3 sky130_fd_sc_hd__dfrbp_1_0[6]/VPWR
rlabel viali 12817 527 12851 561 3 sky130_fd_sc_hd__dfrbp_1_0[6]/VPB
rlabel viali 12725 -17 12759 17 3 sky130_fd_sc_hd__dfrbp_1_0[6]/VGND
rlabel viali 12817 -17 12851 17 3 sky130_fd_sc_hd__dfrbp_1_0[6]/VNB
flabel locali 16293 153 16327 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
flabel locali 14842 221 14876 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/CLK
rlabel viali 16293 153 16327 187 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel locali 16293 127 16341 207 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel locali 16233 207 16341 281 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 16281 147 16339 156 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 16221 193 16279 256 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 16221 184 16339 193 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 15561 184 15691 193 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 15561 156 16339 184 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 15561 147 15691 156 1 sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
flabel locali 16566 218 16595 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/Q
flabel locali 16868 221 16890 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/Q_N
flabel locali 14842 289 14876 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/CLK
flabel locali 15117 289 15151 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[7]/D
rlabel viali 14841 527 14875 561 3 sky130_fd_sc_hd__dfrbp_1_0[7]/VPWR
rlabel viali 14933 527 14967 561 3 sky130_fd_sc_hd__dfrbp_1_0[7]/VPB
rlabel viali 14841 -17 14875 17 3 sky130_fd_sc_hd__dfrbp_1_0[7]/VGND
rlabel viali 14933 -17 14967 17 3 sky130_fd_sc_hd__dfrbp_1_0[7]/VNB
flabel locali 18409 153 18443 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
flabel locali 16958 221 16992 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/CLK
rlabel viali 18409 153 18443 187 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel locali 18409 127 18457 207 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel locali 18349 207 18457 281 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 18397 147 18455 156 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 18337 193 18395 256 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 18337 184 18455 193 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 17677 184 17807 193 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 17677 156 18455 184 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 17677 147 17807 156 1 sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
flabel locali 18682 218 18711 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/Q
flabel locali 18984 221 19006 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/Q_N
flabel locali 16958 289 16992 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/CLK
flabel locali 17233 289 17267 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[8]/D
rlabel viali 16957 527 16991 561 3 sky130_fd_sc_hd__dfrbp_1_0[8]/VPWR
rlabel viali 17049 527 17083 561 3 sky130_fd_sc_hd__dfrbp_1_0[8]/VPB
rlabel viali 16957 -17 16991 17 3 sky130_fd_sc_hd__dfrbp_1_0[8]/VGND
rlabel viali 17049 -17 17083 17 3 sky130_fd_sc_hd__dfrbp_1_0[8]/VNB
flabel locali 20525 153 20559 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
flabel locali 19074 221 19108 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/CLK
rlabel viali 20525 153 20559 187 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel locali 20525 127 20573 207 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel locali 20465 207 20573 281 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 20513 147 20571 156 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 20453 193 20511 256 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 20453 184 20571 193 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 19793 184 19923 193 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 19793 156 20571 184 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 19793 147 19923 156 1 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
flabel locali 20798 218 20827 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/Q
flabel locali 21100 221 21122 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/Q_N
flabel locali 19074 289 19108 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/CLK
flabel locali 19349 289 19383 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[9]/D
rlabel viali 19073 527 19107 561 3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPWR
rlabel viali 19165 527 19199 561 3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB
rlabel viali 19073 -17 19107 17 3 sky130_fd_sc_hd__dfrbp_1_0[9]/VGND
rlabel viali 19165 -17 19199 17 3 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB
flabel locali 22641 153 22675 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
flabel locali 21190 221 21224 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/CLK
rlabel viali 22641 153 22675 187 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel locali 22641 127 22689 207 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel locali 22581 207 22689 281 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 22629 147 22687 156 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 22569 193 22627 256 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 22569 184 22687 193 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 21909 184 22039 193 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 21909 156 22687 184 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 21909 147 22039 156 1 sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
flabel locali 22914 218 22943 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/Q
flabel locali 23216 221 23238 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/Q_N
flabel locali 21190 289 21224 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/CLK
flabel locali 21465 289 21499 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[10]/D
rlabel viali 21189 527 21223 561 3 sky130_fd_sc_hd__dfrbp_1_0[10]/VPWR
rlabel viali 21281 527 21315 561 3 sky130_fd_sc_hd__dfrbp_1_0[10]/VPB
rlabel viali 21189 -17 21223 17 3 sky130_fd_sc_hd__dfrbp_1_0[10]/VGND
rlabel viali 21281 -17 21315 17 3 sky130_fd_sc_hd__dfrbp_1_0[10]/VNB
flabel locali 24757 153 24791 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
flabel locali 23306 221 23340 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/CLK
rlabel viali 24757 153 24791 187 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel locali 24757 127 24805 207 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel locali 24697 207 24805 281 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24745 147 24803 156 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24685 193 24743 256 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24685 184 24803 193 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24025 184 24155 193 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24025 156 24803 184 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 24025 147 24155 156 1 sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
flabel locali 25030 218 25059 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/Q
flabel locali 25332 221 25354 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/Q_N
flabel locali 23306 289 23340 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/CLK
flabel locali 23581 289 23615 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[11]/D
rlabel viali 23305 527 23339 561 3 sky130_fd_sc_hd__dfrbp_1_0[11]/VPWR
rlabel viali 23397 527 23431 561 3 sky130_fd_sc_hd__dfrbp_1_0[11]/VPB
rlabel viali 23305 -17 23339 17 3 sky130_fd_sc_hd__dfrbp_1_0[11]/VGND
rlabel viali 23397 -17 23431 17 3 sky130_fd_sc_hd__dfrbp_1_0[11]/VNB
flabel locali 26873 153 26907 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
flabel locali 25422 221 25456 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/CLK
rlabel viali 26873 153 26907 187 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel locali 26873 127 26921 207 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel locali 26813 207 26921 281 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26861 147 26919 156 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26801 193 26859 256 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26801 184 26919 193 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26141 184 26271 193 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26141 156 26919 184 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 26141 147 26271 156 1 sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
flabel locali 27146 218 27175 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/Q
flabel locali 27448 221 27470 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/Q_N
flabel locali 25422 289 25456 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/CLK
flabel locali 25697 289 25731 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[12]/D
rlabel viali 25421 527 25455 561 3 sky130_fd_sc_hd__dfrbp_1_0[12]/VPWR
rlabel viali 25513 527 25547 561 3 sky130_fd_sc_hd__dfrbp_1_0[12]/VPB
rlabel viali 25421 -17 25455 17 3 sky130_fd_sc_hd__dfrbp_1_0[12]/VGND
rlabel viali 25513 -17 25547 17 3 sky130_fd_sc_hd__dfrbp_1_0[12]/VNB
flabel locali 28989 153 29023 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
flabel locali 27538 221 27572 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/CLK
rlabel viali 28989 153 29023 187 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel locali 28989 127 29037 207 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel locali 28929 207 29037 281 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28977 147 29035 156 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28917 193 28975 256 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28917 184 29035 193 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28257 184 28387 193 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28257 156 29035 184 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 28257 147 28387 156 1 sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
flabel locali 29262 218 29291 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/Q
flabel locali 29564 221 29586 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/Q_N
flabel locali 27538 289 27572 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/CLK
flabel locali 27813 289 27847 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[13]/D
rlabel viali 27537 527 27571 561 3 sky130_fd_sc_hd__dfrbp_1_0[13]/VPWR
rlabel viali 27629 527 27663 561 3 sky130_fd_sc_hd__dfrbp_1_0[13]/VPB
rlabel viali 27537 -17 27571 17 3 sky130_fd_sc_hd__dfrbp_1_0[13]/VGND
rlabel viali 27629 -17 27663 17 3 sky130_fd_sc_hd__dfrbp_1_0[13]/VNB
flabel locali 31105 153 31139 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
flabel locali 29654 221 29688 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/CLK
rlabel viali 31105 153 31139 187 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel locali 31105 127 31153 207 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel locali 31045 207 31153 281 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 31093 147 31151 156 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 31033 193 31091 256 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 31033 184 31151 193 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 30373 184 30503 193 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 30373 156 31151 184 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 30373 147 30503 156 1 sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
flabel locali 31378 218 31407 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/Q
flabel locali 31680 221 31702 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/Q_N
flabel locali 29654 289 29688 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/CLK
flabel locali 29929 289 29963 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[14]/D
rlabel viali 29653 527 29687 561 3 sky130_fd_sc_hd__dfrbp_1_0[14]/VPWR
rlabel viali 29745 527 29779 561 3 sky130_fd_sc_hd__dfrbp_1_0[14]/VPB
rlabel viali 29653 -17 29687 17 3 sky130_fd_sc_hd__dfrbp_1_0[14]/VGND
rlabel viali 29745 -17 29779 17 3 sky130_fd_sc_hd__dfrbp_1_0[14]/VNB
flabel locali 33221 153 33255 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
flabel locali 31770 221 31804 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/CLK
rlabel viali 33221 153 33255 187 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel locali 33221 127 33269 207 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel locali 33161 207 33269 281 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 33209 147 33267 156 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 33149 193 33207 256 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 33149 184 33267 193 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 32489 184 32619 193 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 32489 156 33267 184 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 32489 147 32619 156 1 sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
flabel locali 33494 218 33523 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/Q
flabel locali 33796 221 33818 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/Q_N
flabel locali 31770 289 31804 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/CLK
flabel locali 32045 289 32079 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[15]/D
rlabel viali 31769 527 31803 561 3 sky130_fd_sc_hd__dfrbp_1_0[15]/VPWR
rlabel viali 31861 527 31895 561 3 sky130_fd_sc_hd__dfrbp_1_0[15]/VPB
rlabel viali 31769 -17 31803 17 3 sky130_fd_sc_hd__dfrbp_1_0[15]/VGND
rlabel viali 31861 -17 31895 17 3 sky130_fd_sc_hd__dfrbp_1_0[15]/VNB
flabel locali 35337 153 35371 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
flabel locali 33886 221 33920 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/CLK
rlabel viali 35337 153 35371 187 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel locali 35337 127 35385 207 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel locali 35277 207 35385 281 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 35325 147 35383 156 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 35265 193 35323 256 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 35265 184 35383 193 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 34605 184 34735 193 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 34605 156 35383 184 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 34605 147 34735 156 1 sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
flabel locali 35610 218 35639 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/Q
flabel locali 35912 221 35934 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/Q_N
flabel locali 33886 289 33920 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/CLK
flabel locali 34161 289 34195 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[16]/D
rlabel viali 33885 527 33919 561 3 sky130_fd_sc_hd__dfrbp_1_0[16]/VPWR
rlabel viali 33977 527 34011 561 3 sky130_fd_sc_hd__dfrbp_1_0[16]/VPB
rlabel viali 33885 -17 33919 17 3 sky130_fd_sc_hd__dfrbp_1_0[16]/VGND
rlabel viali 33977 -17 34011 17 3 sky130_fd_sc_hd__dfrbp_1_0[16]/VNB
flabel locali 37453 153 37487 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
flabel locali 36002 221 36036 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/CLK
rlabel viali 37453 153 37487 187 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel locali 37453 127 37501 207 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel locali 37393 207 37501 281 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 37441 147 37499 156 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 37381 193 37439 256 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 37381 184 37499 193 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 36721 184 36851 193 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 36721 156 37499 184 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 36721 147 36851 156 1 sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
flabel locali 37726 218 37755 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/Q
flabel locali 38028 221 38050 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/Q_N
flabel locali 36002 289 36036 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/CLK
flabel locali 36277 289 36311 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[17]/D
rlabel viali 36001 527 36035 561 3 sky130_fd_sc_hd__dfrbp_1_0[17]/VPWR
rlabel viali 36093 527 36127 561 3 sky130_fd_sc_hd__dfrbp_1_0[17]/VPB
rlabel viali 36001 -17 36035 17 3 sky130_fd_sc_hd__dfrbp_1_0[17]/VGND
rlabel viali 36093 -17 36127 17 3 sky130_fd_sc_hd__dfrbp_1_0[17]/VNB
flabel locali 39569 153 39603 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
flabel locali 38118 221 38152 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/CLK
rlabel viali 39569 153 39603 187 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel locali 39569 127 39617 207 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel locali 39509 207 39617 281 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 39557 147 39615 156 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 39497 193 39555 256 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 39497 184 39615 193 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 38837 184 38967 193 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 38837 156 39615 184 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 38837 147 38967 156 1 sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
flabel locali 39842 218 39871 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/Q
flabel locali 40144 221 40166 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/Q_N
flabel locali 38118 289 38152 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/CLK
flabel locali 38393 289 38427 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[18]/D
rlabel viali 38117 527 38151 561 3 sky130_fd_sc_hd__dfrbp_1_0[18]/VPWR
rlabel viali 38209 527 38243 561 3 sky130_fd_sc_hd__dfrbp_1_0[18]/VPB
rlabel viali 38117 -17 38151 17 3 sky130_fd_sc_hd__dfrbp_1_0[18]/VGND
rlabel viali 38209 -17 38243 17 3 sky130_fd_sc_hd__dfrbp_1_0[18]/VNB
flabel locali 41685 153 41719 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
flabel locali 40234 221 40268 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/CLK
rlabel viali 41685 153 41719 187 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel locali 41685 127 41733 207 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel locali 41625 207 41733 281 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 41673 147 41731 156 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 41613 193 41671 256 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 41613 184 41731 193 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 40953 184 41083 193 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 40953 156 41731 184 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 40953 147 41083 156 1 sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
flabel locali 41958 218 41987 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/Q
flabel locali 42260 221 42282 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/Q_N
flabel locali 40234 289 40268 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/CLK
flabel locali 40509 289 40543 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0[19]/D
rlabel viali 40233 527 40267 561 3 sky130_fd_sc_hd__dfrbp_1_0[19]/VPWR
rlabel viali 40325 527 40359 561 3 sky130_fd_sc_hd__dfrbp_1_0[19]/VPB
rlabel viali 40233 -17 40267 17 3 sky130_fd_sc_hd__dfrbp_1_0[19]/VGND
rlabel viali 40325 -17 40359 17 3 sky130_fd_sc_hd__dfrbp_1_0[19]/VNB
<< end >>
