magic
tech sky130A
magscale 1 2
timestamp 1634912350
<< nwell >>
rect 4452 657 4621 750
rect -38 261 2154 656
rect 2428 582 4621 657
rect 2428 261 4620 582
rect 1382 -186 1730 -181
rect 1380 -541 1732 -186
rect 2428 -541 4620 -174
<< pwell >>
rect 903 157 1089 201
rect 1633 157 2104 203
rect 3369 157 3555 201
rect 4099 157 4570 203
rect 1 21 2104 157
rect 2467 21 4570 157
rect 29 -17 63 21
rect 2495 -17 2529 21
rect 1421 -781 1691 -599
rect 3369 -645 3555 -601
rect 4099 -645 4570 -599
rect 2467 -781 4570 -645
rect 1447 -819 1481 -781
rect 2495 -819 2529 -781
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 418 47 448 131
rect 513 47 543 119
rect 609 47 639 119
rect 775 47 805 131
rect 847 47 877 131
rect 979 47 1009 175
rect 1078 47 1108 119
rect 1187 47 1217 119
rect 1283 47 1313 131
rect 1432 47 1462 131
rect 1523 47 1553 131
rect 1711 47 1741 177
rect 1899 47 1929 131
rect 1996 47 2026 177
rect 2545 47 2575 131
rect 2629 47 2659 131
rect 2884 47 2914 131
rect 2979 47 3009 119
rect 3075 47 3105 119
rect 3241 47 3271 131
rect 3313 47 3343 131
rect 3445 47 3475 175
rect 3544 47 3574 119
rect 3653 47 3683 119
rect 3749 47 3779 131
rect 3898 47 3928 131
rect 3989 47 4019 131
rect 4177 47 4207 177
rect 4365 47 4395 131
rect 4462 47 4492 177
rect 1499 -755 1529 -625
rect 1583 -755 1613 -625
rect 2545 -755 2575 -671
rect 2629 -755 2659 -671
rect 2884 -755 2914 -671
rect 2979 -755 3009 -683
rect 3075 -755 3105 -683
rect 3241 -755 3271 -671
rect 3313 -755 3343 -671
rect 3445 -755 3475 -627
rect 3544 -755 3574 -683
rect 3653 -755 3683 -683
rect 3749 -755 3779 -671
rect 3898 -755 3928 -671
rect 3989 -755 4019 -671
rect 4177 -755 4207 -625
rect 4365 -755 4395 -671
rect 4462 -755 4492 -625
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 430 413 460 497
rect 522 413 552 497
rect 621 413 651 497
rect 761 413 791 497
rect 858 413 888 497
rect 1055 329 1085 497
rect 1154 413 1184 497
rect 1240 413 1270 497
rect 1324 413 1354 497
rect 1432 413 1462 497
rect 1516 413 1546 497
rect 1680 297 1710 497
rect 1899 369 1929 497
rect 1996 297 2026 497
rect 2545 363 2575 491
rect 2629 363 2659 491
rect 2896 413 2926 497
rect 2988 413 3018 497
rect 3087 413 3117 497
rect 3227 413 3257 497
rect 3324 413 3354 497
rect 3521 329 3551 497
rect 3620 413 3650 497
rect 3706 413 3736 497
rect 3790 413 3820 497
rect 3898 413 3928 497
rect 3982 413 4012 497
rect 4146 297 4176 497
rect 4365 369 4395 497
rect 4462 297 4492 497
rect 1499 -505 1529 -305
rect 1583 -505 1613 -305
rect 2545 -439 2575 -311
rect 2629 -439 2659 -311
rect 2896 -389 2926 -305
rect 2988 -389 3018 -305
rect 3087 -389 3117 -305
rect 3227 -389 3257 -305
rect 3324 -389 3354 -305
rect 3521 -473 3551 -305
rect 3620 -389 3650 -305
rect 3706 -389 3736 -305
rect 3790 -389 3820 -305
rect 3898 -389 3928 -305
rect 3982 -389 4012 -305
rect 4146 -505 4176 -305
rect 4365 -433 4395 -305
rect 4462 -505 4492 -305
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 313 89 418 131
rect 313 55 325 89
rect 359 55 418 89
rect 313 47 418 55
rect 448 119 498 131
rect 929 131 979 175
rect 657 119 775 131
rect 448 95 513 119
rect 448 61 458 95
rect 492 61 513 95
rect 448 47 513 61
rect 543 95 609 119
rect 543 61 565 95
rect 599 61 609 95
rect 543 47 609 61
rect 639 47 775 119
rect 805 47 847 131
rect 877 93 979 131
rect 877 59 911 93
rect 945 59 979 93
rect 877 47 979 59
rect 1009 119 1063 175
rect 1659 132 1711 177
rect 1233 119 1283 131
rect 1009 89 1078 119
rect 1009 55 1023 89
rect 1057 55 1078 89
rect 1009 47 1078 55
rect 1108 93 1187 119
rect 1108 59 1133 93
rect 1167 59 1187 93
rect 1108 47 1187 59
rect 1217 47 1283 119
rect 1313 89 1432 131
rect 1313 55 1345 89
rect 1379 55 1432 89
rect 1313 47 1432 55
rect 1462 47 1523 131
rect 1553 109 1605 131
rect 1553 75 1563 109
rect 1597 75 1605 109
rect 1553 47 1605 75
rect 1659 98 1667 132
rect 1701 98 1711 132
rect 1659 47 1711 98
rect 1741 165 1793 177
rect 1741 131 1751 165
rect 1785 131 1793 165
rect 1944 131 1996 177
rect 1741 97 1793 131
rect 1741 63 1751 97
rect 1785 63 1793 97
rect 1741 47 1793 63
rect 1847 119 1899 131
rect 1847 85 1855 119
rect 1889 85 1899 119
rect 1847 47 1899 85
rect 1929 113 1996 131
rect 1929 79 1952 113
rect 1986 79 1996 113
rect 1929 47 1996 79
rect 2026 143 2078 177
rect 2026 109 2036 143
rect 2070 109 2078 143
rect 2026 47 2078 109
rect 2493 119 2545 131
rect 2493 85 2501 119
rect 2535 85 2545 119
rect 2493 47 2545 85
rect 2575 93 2629 131
rect 2575 59 2585 93
rect 2619 59 2629 93
rect 2575 47 2629 59
rect 2659 119 2711 131
rect 2659 85 2669 119
rect 2703 85 2711 119
rect 2659 47 2711 85
rect 2779 89 2884 131
rect 2779 55 2791 89
rect 2825 55 2884 89
rect 2779 47 2884 55
rect 2914 119 2964 131
rect 3395 131 3445 175
rect 3123 119 3241 131
rect 2914 95 2979 119
rect 2914 61 2924 95
rect 2958 61 2979 95
rect 2914 47 2979 61
rect 3009 95 3075 119
rect 3009 61 3031 95
rect 3065 61 3075 95
rect 3009 47 3075 61
rect 3105 47 3241 119
rect 3271 47 3313 131
rect 3343 93 3445 131
rect 3343 59 3377 93
rect 3411 59 3445 93
rect 3343 47 3445 59
rect 3475 119 3529 175
rect 4125 132 4177 177
rect 3699 119 3749 131
rect 3475 89 3544 119
rect 3475 55 3489 89
rect 3523 55 3544 89
rect 3475 47 3544 55
rect 3574 93 3653 119
rect 3574 59 3599 93
rect 3633 59 3653 93
rect 3574 47 3653 59
rect 3683 47 3749 119
rect 3779 89 3898 131
rect 3779 55 3811 89
rect 3845 55 3898 89
rect 3779 47 3898 55
rect 3928 47 3989 131
rect 4019 109 4071 131
rect 4019 75 4029 109
rect 4063 75 4071 109
rect 4019 47 4071 75
rect 4125 98 4133 132
rect 4167 98 4177 132
rect 4125 47 4177 98
rect 4207 165 4259 177
rect 4207 131 4217 165
rect 4251 131 4259 165
rect 4410 131 4462 177
rect 4207 97 4259 131
rect 4207 63 4217 97
rect 4251 63 4259 97
rect 4207 47 4259 63
rect 4313 119 4365 131
rect 4313 85 4321 119
rect 4355 85 4365 119
rect 4313 47 4365 85
rect 4395 113 4462 131
rect 4395 79 4418 113
rect 4452 79 4462 113
rect 4395 47 4462 79
rect 4492 143 4544 177
rect 4492 109 4502 143
rect 4536 109 4544 143
rect 4492 47 4544 109
rect 1447 -637 1499 -625
rect 1447 -671 1455 -637
rect 1489 -671 1499 -637
rect 1447 -709 1499 -671
rect 1447 -743 1455 -709
rect 1489 -743 1499 -709
rect 1447 -755 1499 -743
rect 1529 -637 1583 -625
rect 1529 -671 1539 -637
rect 1573 -671 1583 -637
rect 1529 -709 1583 -671
rect 1529 -743 1539 -709
rect 1573 -743 1583 -709
rect 1529 -755 1583 -743
rect 1613 -637 1665 -625
rect 1613 -671 1623 -637
rect 1657 -671 1665 -637
rect 1613 -709 1665 -671
rect 1613 -743 1623 -709
rect 1657 -743 1665 -709
rect 1613 -755 1665 -743
rect 2493 -683 2545 -671
rect 2493 -717 2501 -683
rect 2535 -717 2545 -683
rect 2493 -755 2545 -717
rect 2575 -709 2629 -671
rect 2575 -743 2585 -709
rect 2619 -743 2629 -709
rect 2575 -755 2629 -743
rect 2659 -683 2711 -671
rect 2659 -717 2669 -683
rect 2703 -717 2711 -683
rect 2659 -755 2711 -717
rect 2779 -713 2884 -671
rect 2779 -747 2791 -713
rect 2825 -747 2884 -713
rect 2779 -755 2884 -747
rect 2914 -683 2964 -671
rect 3395 -671 3445 -627
rect 3123 -683 3241 -671
rect 2914 -707 2979 -683
rect 2914 -741 2924 -707
rect 2958 -741 2979 -707
rect 2914 -755 2979 -741
rect 3009 -707 3075 -683
rect 3009 -741 3031 -707
rect 3065 -741 3075 -707
rect 3009 -755 3075 -741
rect 3105 -755 3241 -683
rect 3271 -755 3313 -671
rect 3343 -709 3445 -671
rect 3343 -743 3377 -709
rect 3411 -743 3445 -709
rect 3343 -755 3445 -743
rect 3475 -683 3529 -627
rect 4125 -670 4177 -625
rect 3699 -683 3749 -671
rect 3475 -713 3544 -683
rect 3475 -747 3489 -713
rect 3523 -747 3544 -713
rect 3475 -755 3544 -747
rect 3574 -709 3653 -683
rect 3574 -743 3599 -709
rect 3633 -743 3653 -709
rect 3574 -755 3653 -743
rect 3683 -755 3749 -683
rect 3779 -713 3898 -671
rect 3779 -747 3811 -713
rect 3845 -747 3898 -713
rect 3779 -755 3898 -747
rect 3928 -755 3989 -671
rect 4019 -693 4071 -671
rect 4019 -727 4029 -693
rect 4063 -727 4071 -693
rect 4019 -755 4071 -727
rect 4125 -704 4133 -670
rect 4167 -704 4177 -670
rect 4125 -755 4177 -704
rect 4207 -637 4259 -625
rect 4207 -671 4217 -637
rect 4251 -671 4259 -637
rect 4410 -671 4462 -625
rect 4207 -705 4259 -671
rect 4207 -739 4217 -705
rect 4251 -739 4259 -705
rect 4207 -755 4259 -739
rect 4313 -683 4365 -671
rect 4313 -717 4321 -683
rect 4355 -717 4365 -683
rect 4313 -755 4365 -717
rect 4395 -689 4462 -671
rect 4395 -723 4418 -689
rect 4452 -723 4462 -689
rect 4395 -755 4462 -723
rect 4492 -659 4544 -625
rect 4492 -693 4502 -659
rect 4536 -693 4544 -659
rect 4492 -755 4544 -693
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 378 485 430 497
rect 378 451 386 485
rect 420 451 430 485
rect 378 413 430 451
rect 460 477 522 497
rect 460 443 470 477
rect 504 443 522 477
rect 460 413 522 443
rect 552 483 621 497
rect 552 449 563 483
rect 597 449 621 483
rect 552 413 621 449
rect 651 459 761 497
rect 651 425 717 459
rect 751 425 761 459
rect 651 413 761 425
rect 791 475 858 497
rect 791 441 814 475
rect 848 441 858 475
rect 791 413 858 441
rect 888 459 940 497
rect 888 425 898 459
rect 932 425 940 459
rect 888 413 940 425
rect 1003 485 1055 497
rect 1003 451 1011 485
rect 1045 451 1055 485
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 1003 329 1055 451
rect 1085 477 1154 497
rect 1085 443 1099 477
rect 1133 443 1154 477
rect 1085 413 1154 443
rect 1184 484 1240 497
rect 1184 450 1196 484
rect 1230 450 1240 484
rect 1184 413 1240 450
rect 1270 413 1324 497
rect 1354 485 1432 497
rect 1354 451 1388 485
rect 1422 451 1432 485
rect 1354 413 1432 451
rect 1462 459 1516 497
rect 1462 425 1472 459
rect 1506 425 1516 459
rect 1462 413 1516 425
rect 1546 485 1680 497
rect 1546 451 1558 485
rect 1592 451 1636 485
rect 1670 451 1680 485
rect 1546 413 1680 451
rect 1085 329 1139 413
rect 1630 297 1680 413
rect 1710 477 1766 497
rect 1710 443 1720 477
rect 1754 443 1766 477
rect 1710 409 1766 443
rect 1710 375 1720 409
rect 1754 375 1766 409
rect 1710 341 1766 375
rect 1847 485 1899 497
rect 1847 451 1855 485
rect 1889 451 1899 485
rect 1847 417 1899 451
rect 1847 383 1855 417
rect 1889 383 1899 417
rect 1847 369 1899 383
rect 1929 485 1996 497
rect 1929 451 1952 485
rect 1986 451 1996 485
rect 1929 417 1996 451
rect 1929 383 1952 417
rect 1986 383 1996 417
rect 1929 369 1996 383
rect 1710 307 1720 341
rect 1754 307 1766 341
rect 1710 297 1766 307
rect 1944 349 1996 369
rect 1944 315 1952 349
rect 1986 315 1996 349
rect 1944 297 1996 315
rect 2026 449 2078 497
rect 2026 415 2036 449
rect 2070 415 2078 449
rect 2026 381 2078 415
rect 2026 347 2036 381
rect 2070 347 2078 381
rect 2493 477 2545 491
rect 2493 443 2501 477
rect 2535 443 2545 477
rect 2493 409 2545 443
rect 2493 375 2501 409
rect 2535 375 2545 409
rect 2493 363 2545 375
rect 2575 461 2629 491
rect 2575 427 2585 461
rect 2619 427 2629 461
rect 2575 363 2629 427
rect 2659 477 2711 491
rect 2659 443 2669 477
rect 2703 443 2711 477
rect 2659 409 2711 443
rect 2844 485 2896 497
rect 2844 451 2852 485
rect 2886 451 2896 485
rect 2844 413 2896 451
rect 2926 477 2988 497
rect 2926 443 2936 477
rect 2970 443 2988 477
rect 2926 413 2988 443
rect 3018 483 3087 497
rect 3018 449 3029 483
rect 3063 449 3087 483
rect 3018 413 3087 449
rect 3117 459 3227 497
rect 3117 425 3183 459
rect 3217 425 3227 459
rect 3117 413 3227 425
rect 3257 475 3324 497
rect 3257 441 3280 475
rect 3314 441 3324 475
rect 3257 413 3324 441
rect 3354 459 3406 497
rect 3354 425 3364 459
rect 3398 425 3406 459
rect 3354 413 3406 425
rect 3469 485 3521 497
rect 3469 451 3477 485
rect 3511 451 3521 485
rect 2659 375 2669 409
rect 2703 375 2711 409
rect 2659 363 2711 375
rect 2026 297 2078 347
rect 3469 329 3521 451
rect 3551 477 3620 497
rect 3551 443 3565 477
rect 3599 443 3620 477
rect 3551 413 3620 443
rect 3650 484 3706 497
rect 3650 450 3662 484
rect 3696 450 3706 484
rect 3650 413 3706 450
rect 3736 413 3790 497
rect 3820 485 3898 497
rect 3820 451 3854 485
rect 3888 451 3898 485
rect 3820 413 3898 451
rect 3928 459 3982 497
rect 3928 425 3938 459
rect 3972 425 3982 459
rect 3928 413 3982 425
rect 4012 485 4146 497
rect 4012 451 4024 485
rect 4058 451 4102 485
rect 4136 451 4146 485
rect 4012 413 4146 451
rect 3551 329 3605 413
rect 4096 297 4146 413
rect 4176 477 4232 497
rect 4176 443 4186 477
rect 4220 443 4232 477
rect 4176 409 4232 443
rect 4176 375 4186 409
rect 4220 375 4232 409
rect 4176 341 4232 375
rect 4313 485 4365 497
rect 4313 451 4321 485
rect 4355 451 4365 485
rect 4313 417 4365 451
rect 4313 383 4321 417
rect 4355 383 4365 417
rect 4313 369 4365 383
rect 4395 485 4462 497
rect 4395 451 4418 485
rect 4452 451 4462 485
rect 4395 417 4462 451
rect 4395 383 4418 417
rect 4452 383 4462 417
rect 4395 369 4462 383
rect 4176 307 4186 341
rect 4220 307 4232 341
rect 4176 297 4232 307
rect 4410 349 4462 369
rect 4410 315 4418 349
rect 4452 315 4462 349
rect 4410 297 4462 315
rect 4492 449 4544 497
rect 4492 415 4502 449
rect 4536 415 4544 449
rect 4492 381 4544 415
rect 4492 347 4502 381
rect 4536 347 4544 381
rect 4492 297 4544 347
rect 1447 -317 1499 -305
rect 1447 -351 1455 -317
rect 1489 -351 1499 -317
rect 1447 -385 1499 -351
rect 1447 -419 1455 -385
rect 1489 -419 1499 -385
rect 1447 -453 1499 -419
rect 1447 -487 1455 -453
rect 1489 -487 1499 -453
rect 1447 -505 1499 -487
rect 1529 -317 1583 -305
rect 1529 -351 1539 -317
rect 1573 -351 1583 -317
rect 1529 -385 1583 -351
rect 1529 -419 1539 -385
rect 1573 -419 1583 -385
rect 1529 -453 1583 -419
rect 1529 -487 1539 -453
rect 1573 -487 1583 -453
rect 1529 -505 1583 -487
rect 1613 -317 1665 -305
rect 1613 -351 1623 -317
rect 1657 -351 1665 -317
rect 1613 -385 1665 -351
rect 1613 -419 1623 -385
rect 1657 -419 1665 -385
rect 1613 -453 1665 -419
rect 2493 -325 2545 -311
rect 2493 -359 2501 -325
rect 2535 -359 2545 -325
rect 2493 -393 2545 -359
rect 2493 -427 2501 -393
rect 2535 -427 2545 -393
rect 2493 -439 2545 -427
rect 2575 -341 2629 -311
rect 2575 -375 2585 -341
rect 2619 -375 2629 -341
rect 2575 -439 2629 -375
rect 2659 -325 2711 -311
rect 2659 -359 2669 -325
rect 2703 -359 2711 -325
rect 2659 -393 2711 -359
rect 2844 -317 2896 -305
rect 2844 -351 2852 -317
rect 2886 -351 2896 -317
rect 2844 -389 2896 -351
rect 2926 -325 2988 -305
rect 2926 -359 2936 -325
rect 2970 -359 2988 -325
rect 2926 -389 2988 -359
rect 3018 -319 3087 -305
rect 3018 -353 3029 -319
rect 3063 -353 3087 -319
rect 3018 -389 3087 -353
rect 3117 -343 3227 -305
rect 3117 -377 3183 -343
rect 3217 -377 3227 -343
rect 3117 -389 3227 -377
rect 3257 -327 3324 -305
rect 3257 -361 3280 -327
rect 3314 -361 3324 -327
rect 3257 -389 3324 -361
rect 3354 -343 3406 -305
rect 3354 -377 3364 -343
rect 3398 -377 3406 -343
rect 3354 -389 3406 -377
rect 3469 -317 3521 -305
rect 3469 -351 3477 -317
rect 3511 -351 3521 -317
rect 2659 -427 2669 -393
rect 2703 -427 2711 -393
rect 2659 -439 2711 -427
rect 1613 -487 1623 -453
rect 1657 -487 1665 -453
rect 1613 -505 1665 -487
rect 3469 -473 3521 -351
rect 3551 -325 3620 -305
rect 3551 -359 3565 -325
rect 3599 -359 3620 -325
rect 3551 -389 3620 -359
rect 3650 -318 3706 -305
rect 3650 -352 3662 -318
rect 3696 -352 3706 -318
rect 3650 -389 3706 -352
rect 3736 -389 3790 -305
rect 3820 -317 3898 -305
rect 3820 -351 3854 -317
rect 3888 -351 3898 -317
rect 3820 -389 3898 -351
rect 3928 -343 3982 -305
rect 3928 -377 3938 -343
rect 3972 -377 3982 -343
rect 3928 -389 3982 -377
rect 4012 -317 4146 -305
rect 4012 -351 4024 -317
rect 4058 -351 4102 -317
rect 4136 -351 4146 -317
rect 4012 -389 4146 -351
rect 3551 -473 3605 -389
rect 4096 -505 4146 -389
rect 4176 -325 4232 -305
rect 4176 -359 4186 -325
rect 4220 -359 4232 -325
rect 4176 -393 4232 -359
rect 4176 -427 4186 -393
rect 4220 -427 4232 -393
rect 4176 -461 4232 -427
rect 4313 -317 4365 -305
rect 4313 -351 4321 -317
rect 4355 -351 4365 -317
rect 4313 -385 4365 -351
rect 4313 -419 4321 -385
rect 4355 -419 4365 -385
rect 4313 -433 4365 -419
rect 4395 -317 4462 -305
rect 4395 -351 4418 -317
rect 4452 -351 4462 -317
rect 4395 -385 4462 -351
rect 4395 -419 4418 -385
rect 4452 -419 4462 -385
rect 4395 -433 4462 -419
rect 4176 -495 4186 -461
rect 4220 -495 4232 -461
rect 4176 -505 4232 -495
rect 4410 -453 4462 -433
rect 4410 -487 4418 -453
rect 4452 -487 4462 -453
rect 4410 -505 4462 -487
rect 4492 -353 4544 -305
rect 4492 -387 4502 -353
rect 4536 -387 4544 -353
rect 4492 -421 4544 -387
rect 4492 -455 4502 -421
rect 4536 -455 4544 -421
rect 4492 -505 4544 -455
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 325 55 359 89
rect 458 61 492 95
rect 565 61 599 95
rect 911 59 945 93
rect 1023 55 1057 89
rect 1133 59 1167 93
rect 1345 55 1379 89
rect 1563 75 1597 109
rect 1667 98 1701 132
rect 1751 131 1785 165
rect 1751 63 1785 97
rect 1855 85 1889 119
rect 1952 79 1986 113
rect 2036 109 2070 143
rect 2501 85 2535 119
rect 2585 59 2619 93
rect 2669 85 2703 119
rect 2791 55 2825 89
rect 2924 61 2958 95
rect 3031 61 3065 95
rect 3377 59 3411 93
rect 3489 55 3523 89
rect 3599 59 3633 93
rect 3811 55 3845 89
rect 4029 75 4063 109
rect 4133 98 4167 132
rect 4217 131 4251 165
rect 4217 63 4251 97
rect 4321 85 4355 119
rect 4418 79 4452 113
rect 4502 109 4536 143
rect 1455 -671 1489 -637
rect 1455 -743 1489 -709
rect 1539 -671 1573 -637
rect 1539 -743 1573 -709
rect 1623 -671 1657 -637
rect 1623 -743 1657 -709
rect 2501 -717 2535 -683
rect 2585 -743 2619 -709
rect 2669 -717 2703 -683
rect 2791 -747 2825 -713
rect 2924 -741 2958 -707
rect 3031 -741 3065 -707
rect 3377 -743 3411 -709
rect 3489 -747 3523 -713
rect 3599 -743 3633 -709
rect 3811 -747 3845 -713
rect 4029 -727 4063 -693
rect 4133 -704 4167 -670
rect 4217 -671 4251 -637
rect 4217 -739 4251 -705
rect 4321 -717 4355 -683
rect 4418 -723 4452 -689
rect 4502 -693 4536 -659
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 386 451 420 485
rect 470 443 504 477
rect 563 449 597 483
rect 717 425 751 459
rect 814 441 848 475
rect 898 425 932 459
rect 1011 451 1045 485
rect 203 375 237 409
rect 1099 443 1133 477
rect 1196 450 1230 484
rect 1388 451 1422 485
rect 1472 425 1506 459
rect 1558 451 1592 485
rect 1636 451 1670 485
rect 1720 443 1754 477
rect 1720 375 1754 409
rect 1855 451 1889 485
rect 1855 383 1889 417
rect 1952 451 1986 485
rect 1952 383 1986 417
rect 1720 307 1754 341
rect 1952 315 1986 349
rect 2036 415 2070 449
rect 2036 347 2070 381
rect 2501 443 2535 477
rect 2501 375 2535 409
rect 2585 427 2619 461
rect 2669 443 2703 477
rect 2852 451 2886 485
rect 2936 443 2970 477
rect 3029 449 3063 483
rect 3183 425 3217 459
rect 3280 441 3314 475
rect 3364 425 3398 459
rect 3477 451 3511 485
rect 2669 375 2703 409
rect 3565 443 3599 477
rect 3662 450 3696 484
rect 3854 451 3888 485
rect 3938 425 3972 459
rect 4024 451 4058 485
rect 4102 451 4136 485
rect 4186 443 4220 477
rect 4186 375 4220 409
rect 4321 451 4355 485
rect 4321 383 4355 417
rect 4418 451 4452 485
rect 4418 383 4452 417
rect 4186 307 4220 341
rect 4418 315 4452 349
rect 4502 415 4536 449
rect 4502 347 4536 381
rect 1455 -351 1489 -317
rect 1455 -419 1489 -385
rect 1455 -487 1489 -453
rect 1539 -351 1573 -317
rect 1539 -419 1573 -385
rect 1539 -487 1573 -453
rect 1623 -351 1657 -317
rect 1623 -419 1657 -385
rect 2501 -359 2535 -325
rect 2501 -427 2535 -393
rect 2585 -375 2619 -341
rect 2669 -359 2703 -325
rect 2852 -351 2886 -317
rect 2936 -359 2970 -325
rect 3029 -353 3063 -319
rect 3183 -377 3217 -343
rect 3280 -361 3314 -327
rect 3364 -377 3398 -343
rect 3477 -351 3511 -317
rect 2669 -427 2703 -393
rect 1623 -487 1657 -453
rect 3565 -359 3599 -325
rect 3662 -352 3696 -318
rect 3854 -351 3888 -317
rect 3938 -377 3972 -343
rect 4024 -351 4058 -317
rect 4102 -351 4136 -317
rect 4186 -359 4220 -325
rect 4186 -427 4220 -393
rect 4321 -351 4355 -317
rect 4321 -419 4355 -385
rect 4418 -351 4452 -317
rect 4418 -419 4452 -385
rect 4186 -495 4220 -461
rect 4418 -487 4452 -453
rect 4502 -387 4536 -353
rect 4502 -455 4536 -421
<< psubdiff >>
rect 0 -45 29 -11
rect 63 -45 121 -11
rect 155 -45 213 -11
rect 247 -45 305 -11
rect 339 -45 397 -11
rect 431 -45 489 -11
rect 523 -45 581 -11
rect 615 -45 673 -11
rect 707 -45 765 -11
rect 799 -45 857 -11
rect 891 -45 949 -11
rect 983 -45 1041 -11
rect 1075 -45 1133 -11
rect 1167 -45 1225 -11
rect 1259 -45 1317 -11
rect 1351 -45 1409 -11
rect 1443 -45 1501 -11
rect 1535 -45 1593 -11
rect 1627 -45 1685 -11
rect 1719 -45 1777 -11
rect 1811 -45 1869 -11
rect 1903 -45 1961 -11
rect 1995 -45 2053 -11
rect 2087 -45 2116 -11
rect 2466 -44 2495 -10
rect 2529 -44 2587 -10
rect 2621 -44 2679 -10
rect 2713 -44 2771 -10
rect 2805 -44 2863 -10
rect 2897 -44 2955 -10
rect 2989 -44 3047 -10
rect 3081 -44 3139 -10
rect 3173 -44 3231 -10
rect 3265 -44 3323 -10
rect 3357 -44 3415 -10
rect 3449 -44 3507 -10
rect 3541 -44 3599 -10
rect 3633 -44 3691 -10
rect 3725 -44 3783 -10
rect 3817 -44 3875 -10
rect 3909 -44 3967 -10
rect 4001 -44 4059 -10
rect 4093 -44 4151 -10
rect 4185 -44 4243 -10
rect 4277 -44 4335 -10
rect 4369 -44 4427 -10
rect 4461 -44 4519 -10
rect 4553 -44 4582 -10
rect 1418 -845 1447 -811
rect 1481 -845 1539 -811
rect 1573 -845 1631 -811
rect 1665 -845 1694 -811
rect 2465 -847 2495 -813
rect 2529 -847 2587 -813
rect 2621 -847 2679 -813
rect 2713 -847 2771 -813
rect 2805 -847 2863 -813
rect 2897 -847 2955 -813
rect 2989 -847 3047 -813
rect 3081 -847 3139 -813
rect 3173 -847 3231 -813
rect 3265 -847 3323 -813
rect 3357 -847 3415 -813
rect 3449 -847 3507 -813
rect 3541 -847 3599 -813
rect 3633 -847 3691 -813
rect 3725 -847 3783 -813
rect 3817 -847 3875 -813
rect 3909 -847 3967 -813
rect 4001 -847 4059 -813
rect 4093 -847 4151 -813
rect 4185 -847 4243 -813
rect 4277 -847 4335 -813
rect 4369 -847 4427 -813
rect 4461 -847 4519 -813
rect 4553 -847 4582 -813
<< nsubdiff >>
rect 0 551 29 585
rect 63 551 121 585
rect 155 551 213 585
rect 247 551 305 585
rect 339 551 397 585
rect 431 551 489 585
rect 523 551 581 585
rect 615 551 673 585
rect 707 551 765 585
rect 799 551 857 585
rect 891 551 949 585
rect 983 551 1041 585
rect 1075 551 1133 585
rect 1167 551 1225 585
rect 1259 551 1317 585
rect 1351 551 1409 585
rect 1443 551 1501 585
rect 1535 551 1593 585
rect 1627 551 1685 585
rect 1719 551 1777 585
rect 1811 551 1869 585
rect 1903 551 1961 585
rect 1995 551 2053 585
rect 2087 551 2117 585
rect 2466 551 2495 585
rect 2529 551 2587 585
rect 2621 551 2679 585
rect 2713 551 2771 585
rect 2805 551 2863 585
rect 2897 551 2955 585
rect 2989 551 3047 585
rect 3081 551 3139 585
rect 3173 551 3231 585
rect 3265 551 3323 585
rect 3357 551 3415 585
rect 3449 551 3507 585
rect 3541 551 3599 585
rect 3633 551 3691 585
rect 3725 551 3783 585
rect 3817 551 3875 585
rect 3909 551 3967 585
rect 4001 551 4059 585
rect 4093 551 4151 585
rect 4185 551 4243 585
rect 4277 551 4335 585
rect 4369 551 4427 585
rect 4461 551 4519 585
rect 4553 551 4583 585
rect 1418 -251 1447 -217
rect 1481 -251 1539 -217
rect 1573 -251 1631 -217
rect 1665 -251 1694 -217
rect 2466 -250 2495 -216
rect 2529 -250 2587 -216
rect 2621 -250 2679 -216
rect 2713 -250 2771 -216
rect 2805 -250 2863 -216
rect 2897 -250 2955 -216
rect 2989 -250 3047 -216
rect 3081 -250 3139 -216
rect 3173 -250 3231 -216
rect 3265 -250 3323 -216
rect 3357 -250 3415 -216
rect 3449 -250 3507 -216
rect 3541 -250 3599 -216
rect 3633 -250 3691 -216
rect 3725 -250 3783 -216
rect 3817 -250 3875 -216
rect 3909 -250 3967 -216
rect 4001 -250 4059 -216
rect 4093 -250 4151 -216
rect 4185 -250 4243 -216
rect 4277 -250 4335 -216
rect 4369 -250 4427 -216
rect 4461 -250 4519 -216
rect 4553 -250 4582 -216
<< psubdiffcont >>
rect 29 -45 63 -11
rect 121 -45 155 -11
rect 213 -45 247 -11
rect 305 -45 339 -11
rect 397 -45 431 -11
rect 489 -45 523 -11
rect 581 -45 615 -11
rect 673 -45 707 -11
rect 765 -45 799 -11
rect 857 -45 891 -11
rect 949 -45 983 -11
rect 1041 -45 1075 -11
rect 1133 -45 1167 -11
rect 1225 -45 1259 -11
rect 1317 -45 1351 -11
rect 1409 -45 1443 -11
rect 1501 -45 1535 -11
rect 1593 -45 1627 -11
rect 1685 -45 1719 -11
rect 1777 -45 1811 -11
rect 1869 -45 1903 -11
rect 1961 -45 1995 -11
rect 2053 -45 2087 -11
rect 2495 -44 2529 -10
rect 2587 -44 2621 -10
rect 2679 -44 2713 -10
rect 2771 -44 2805 -10
rect 2863 -44 2897 -10
rect 2955 -44 2989 -10
rect 3047 -44 3081 -10
rect 3139 -44 3173 -10
rect 3231 -44 3265 -10
rect 3323 -44 3357 -10
rect 3415 -44 3449 -10
rect 3507 -44 3541 -10
rect 3599 -44 3633 -10
rect 3691 -44 3725 -10
rect 3783 -44 3817 -10
rect 3875 -44 3909 -10
rect 3967 -44 4001 -10
rect 4059 -44 4093 -10
rect 4151 -44 4185 -10
rect 4243 -44 4277 -10
rect 4335 -44 4369 -10
rect 4427 -44 4461 -10
rect 4519 -44 4553 -10
rect 1447 -845 1481 -811
rect 1539 -845 1573 -811
rect 1631 -845 1665 -811
rect 2495 -847 2529 -813
rect 2587 -847 2621 -813
rect 2679 -847 2713 -813
rect 2771 -847 2805 -813
rect 2863 -847 2897 -813
rect 2955 -847 2989 -813
rect 3047 -847 3081 -813
rect 3139 -847 3173 -813
rect 3231 -847 3265 -813
rect 3323 -847 3357 -813
rect 3415 -847 3449 -813
rect 3507 -847 3541 -813
rect 3599 -847 3633 -813
rect 3691 -847 3725 -813
rect 3783 -847 3817 -813
rect 3875 -847 3909 -813
rect 3967 -847 4001 -813
rect 4059 -847 4093 -813
rect 4151 -847 4185 -813
rect 4243 -847 4277 -813
rect 4335 -847 4369 -813
rect 4427 -847 4461 -813
rect 4519 -847 4553 -813
<< nsubdiffcont >>
rect 29 551 63 585
rect 121 551 155 585
rect 213 551 247 585
rect 305 551 339 585
rect 397 551 431 585
rect 489 551 523 585
rect 581 551 615 585
rect 673 551 707 585
rect 765 551 799 585
rect 857 551 891 585
rect 949 551 983 585
rect 1041 551 1075 585
rect 1133 551 1167 585
rect 1225 551 1259 585
rect 1317 551 1351 585
rect 1409 551 1443 585
rect 1501 551 1535 585
rect 1593 551 1627 585
rect 1685 551 1719 585
rect 1777 551 1811 585
rect 1869 551 1903 585
rect 1961 551 1995 585
rect 2053 551 2087 585
rect 2495 551 2529 585
rect 2587 551 2621 585
rect 2679 551 2713 585
rect 2771 551 2805 585
rect 2863 551 2897 585
rect 2955 551 2989 585
rect 3047 551 3081 585
rect 3139 551 3173 585
rect 3231 551 3265 585
rect 3323 551 3357 585
rect 3415 551 3449 585
rect 3507 551 3541 585
rect 3599 551 3633 585
rect 3691 551 3725 585
rect 3783 551 3817 585
rect 3875 551 3909 585
rect 3967 551 4001 585
rect 4059 551 4093 585
rect 4151 551 4185 585
rect 4243 551 4277 585
rect 4335 551 4369 585
rect 4427 551 4461 585
rect 4519 551 4553 585
rect 1447 -251 1481 -217
rect 1539 -251 1573 -217
rect 1631 -251 1665 -217
rect 2495 -250 2529 -216
rect 2587 -250 2621 -216
rect 2679 -250 2713 -216
rect 2771 -250 2805 -216
rect 2863 -250 2897 -216
rect 2955 -250 2989 -216
rect 3047 -250 3081 -216
rect 3139 -250 3173 -216
rect 3231 -250 3265 -216
rect 3323 -250 3357 -216
rect 3415 -250 3449 -216
rect 3507 -250 3541 -216
rect 3599 -250 3633 -216
rect 3691 -250 3725 -216
rect 3783 -250 3817 -216
rect 3875 -250 3909 -216
rect 3967 -250 4001 -216
rect 4059 -250 4093 -216
rect 4151 -250 4185 -216
rect 4243 -250 4277 -216
rect 4335 -250 4369 -216
rect 4427 -250 4461 -216
rect 4519 -250 4553 -216
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 430 497 460 523
rect 522 497 552 523
rect 621 497 651 523
rect 761 497 791 523
rect 858 497 888 523
rect 1055 497 1085 523
rect 1154 497 1184 523
rect 1240 497 1270 523
rect 1324 497 1354 523
rect 1432 497 1462 523
rect 1516 497 1546 523
rect 1680 497 1710 523
rect 1899 497 1929 523
rect 1996 497 2026 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 265 76 318
rect 163 274 193 363
rect 430 326 460 413
rect 522 375 552 413
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 331 310 460 326
rect 506 365 572 375
rect 506 331 522 365
rect 556 331 572 365
rect 506 321 572 331
rect 331 276 341 310
rect 375 296 460 310
rect 375 276 448 296
rect 621 279 651 413
rect 761 355 791 413
rect 761 339 816 355
rect 761 305 771 339
rect 805 305 816 339
rect 761 289 816 305
rect 331 260 448 276
rect 118 220 193 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 418 131 448 260
rect 513 249 651 279
rect 513 219 544 249
rect 490 203 544 219
rect 490 169 500 203
rect 534 169 544 203
rect 490 153 544 169
rect 586 197 652 207
rect 586 163 602 197
rect 636 163 652 197
rect 586 153 652 163
rect 513 119 543 153
rect 609 119 639 153
rect 775 131 805 289
rect 858 219 888 413
rect 1055 314 1085 329
rect 979 284 1085 314
rect 979 267 1009 284
rect 943 251 1009 267
rect 847 203 901 219
rect 847 169 857 203
rect 891 169 901 203
rect 943 217 953 251
rect 987 217 1009 251
rect 1154 279 1184 413
rect 1240 381 1270 413
rect 1226 365 1280 381
rect 1226 331 1236 365
rect 1270 331 1280 365
rect 1226 315 1280 331
rect 1154 267 1204 279
rect 1154 255 1217 267
rect 1154 249 1241 255
rect 1175 239 1241 249
rect 1175 237 1197 239
rect 943 201 1009 217
rect 979 175 1009 201
rect 1078 191 1145 207
rect 847 153 901 169
rect 847 131 877 153
rect 1078 157 1101 191
rect 1135 157 1145 191
rect 1078 141 1145 157
rect 1187 205 1197 237
rect 1231 205 1241 239
rect 1187 189 1241 205
rect 1324 229 1354 413
rect 1432 257 1462 413
rect 1516 365 1546 413
rect 1504 349 1558 365
rect 1504 315 1514 349
rect 1548 315 1558 349
rect 1504 299 1558 315
rect 1427 241 1481 257
rect 1324 213 1385 229
rect 1324 193 1341 213
rect 1078 119 1108 141
rect 1187 119 1217 189
rect 1283 179 1341 193
rect 1375 179 1385 213
rect 1427 207 1437 241
rect 1471 207 1481 241
rect 1427 191 1481 207
rect 1283 163 1385 179
rect 1283 131 1313 163
rect 1432 131 1462 191
rect 1523 131 1553 299
rect 1899 333 1929 369
rect 1888 303 1929 333
rect 1680 265 1710 297
rect 1888 265 1918 303
rect 2545 491 2575 517
rect 2629 491 2659 517
rect 2896 497 2926 523
rect 2988 497 3018 523
rect 3087 497 3117 523
rect 3227 497 3257 523
rect 3324 497 3354 523
rect 3521 497 3551 523
rect 3620 497 3650 523
rect 3706 497 3736 523
rect 3790 497 3820 523
rect 3898 497 3928 523
rect 3982 497 4012 523
rect 4146 497 4176 523
rect 4365 497 4395 523
rect 4462 497 4492 523
rect 2545 348 2575 363
rect 2512 318 2575 348
rect 1996 265 2026 297
rect 2512 265 2542 318
rect 2629 274 2659 363
rect 2896 326 2926 413
rect 2988 375 3018 413
rect 1609 249 1918 265
rect 1609 215 1637 249
rect 1671 215 1918 249
rect 1609 199 1918 215
rect 1967 249 2026 265
rect 1967 215 1977 249
rect 2011 215 2026 249
rect 1967 199 2026 215
rect 2488 249 2542 265
rect 2488 215 2498 249
rect 2532 215 2542 249
rect 2584 264 2659 274
rect 2584 230 2600 264
rect 2634 230 2659 264
rect 2797 310 2926 326
rect 2972 365 3038 375
rect 2972 331 2988 365
rect 3022 331 3038 365
rect 2972 321 3038 331
rect 2797 276 2807 310
rect 2841 296 2926 310
rect 2841 276 2914 296
rect 3087 279 3117 413
rect 3227 355 3257 413
rect 3227 339 3282 355
rect 3227 305 3237 339
rect 3271 305 3282 339
rect 3227 289 3282 305
rect 2797 260 2914 276
rect 2584 220 2659 230
rect 2488 199 2542 215
rect 1711 177 1741 199
rect 1888 176 1918 199
rect 1996 177 2026 199
rect 1888 146 1929 176
rect 1899 131 1929 146
rect 2512 176 2542 199
rect 2512 146 2575 176
rect 2545 131 2575 146
rect 2629 131 2659 220
rect 2884 131 2914 260
rect 2979 249 3117 279
rect 2979 219 3010 249
rect 2956 203 3010 219
rect 2956 169 2966 203
rect 3000 169 3010 203
rect 2956 153 3010 169
rect 3052 197 3118 207
rect 3052 163 3068 197
rect 3102 163 3118 197
rect 3052 153 3118 163
rect 2979 119 3009 153
rect 3075 119 3105 153
rect 3241 131 3271 289
rect 3324 219 3354 413
rect 3521 314 3551 329
rect 3445 284 3551 314
rect 3445 267 3475 284
rect 3409 251 3475 267
rect 3313 203 3367 219
rect 3313 169 3323 203
rect 3357 169 3367 203
rect 3409 217 3419 251
rect 3453 217 3475 251
rect 3620 279 3650 413
rect 3706 381 3736 413
rect 3692 365 3746 381
rect 3692 331 3702 365
rect 3736 331 3746 365
rect 3692 315 3746 331
rect 3620 267 3670 279
rect 3620 255 3683 267
rect 3620 249 3707 255
rect 3641 239 3707 249
rect 3641 237 3663 239
rect 3409 201 3475 217
rect 3445 175 3475 201
rect 3544 191 3611 207
rect 3313 153 3367 169
rect 3313 131 3343 153
rect 3544 157 3567 191
rect 3601 157 3611 191
rect 3544 141 3611 157
rect 3653 205 3663 237
rect 3697 205 3707 239
rect 3653 189 3707 205
rect 3790 229 3820 413
rect 3898 257 3928 413
rect 3982 365 4012 413
rect 3970 349 4024 365
rect 3970 315 3980 349
rect 4014 315 4024 349
rect 3970 299 4024 315
rect 3893 241 3947 257
rect 3790 213 3851 229
rect 3790 193 3807 213
rect 3544 119 3574 141
rect 3653 119 3683 189
rect 3749 179 3807 193
rect 3841 179 3851 213
rect 3893 207 3903 241
rect 3937 207 3947 241
rect 3893 191 3947 207
rect 3749 163 3851 179
rect 3749 131 3779 163
rect 3898 131 3928 191
rect 3989 131 4019 299
rect 4365 333 4395 369
rect 4354 303 4395 333
rect 4146 265 4176 297
rect 4354 265 4384 303
rect 4462 265 4492 297
rect 4075 249 4384 265
rect 4075 215 4103 249
rect 4137 215 4384 249
rect 4075 199 4384 215
rect 4433 249 4492 265
rect 4433 215 4443 249
rect 4477 215 4492 249
rect 4433 199 4492 215
rect 4177 177 4207 199
rect 4354 176 4384 199
rect 4462 177 4492 199
rect 4354 146 4395 176
rect 4365 131 4395 146
rect 79 21 109 47
rect 163 21 193 47
rect 418 21 448 47
rect 513 21 543 47
rect 609 21 639 47
rect 775 21 805 47
rect 847 21 877 47
rect 979 21 1009 47
rect 1078 21 1108 47
rect 1187 21 1217 47
rect 1283 21 1313 47
rect 1432 21 1462 47
rect 1523 21 1553 47
rect 1711 21 1741 47
rect 1899 21 1929 47
rect 1996 21 2026 47
rect 2545 21 2575 47
rect 2629 21 2659 47
rect 2884 21 2914 47
rect 2979 21 3009 47
rect 3075 21 3105 47
rect 3241 21 3271 47
rect 3313 21 3343 47
rect 3445 21 3475 47
rect 3544 21 3574 47
rect 3653 21 3683 47
rect 3749 21 3779 47
rect 3898 21 3928 47
rect 3989 21 4019 47
rect 4177 21 4207 47
rect 4365 21 4395 47
rect 4462 21 4492 47
rect 1499 -305 1529 -279
rect 1583 -305 1613 -279
rect 2545 -311 2575 -285
rect 2629 -311 2659 -285
rect 2896 -305 2926 -279
rect 2988 -305 3018 -279
rect 3087 -305 3117 -279
rect 3227 -305 3257 -279
rect 3324 -305 3354 -279
rect 3521 -305 3551 -279
rect 3620 -305 3650 -279
rect 3706 -305 3736 -279
rect 3790 -305 3820 -279
rect 3898 -305 3928 -279
rect 3982 -305 4012 -279
rect 4146 -305 4176 -279
rect 4365 -305 4395 -279
rect 4462 -305 4492 -279
rect 2545 -454 2575 -439
rect 2512 -484 2575 -454
rect 1499 -537 1529 -505
rect 1583 -537 1613 -505
rect 2512 -537 2542 -484
rect 2629 -528 2659 -439
rect 2896 -476 2926 -389
rect 2988 -427 3018 -389
rect 1439 -553 1613 -537
rect 1439 -587 1455 -553
rect 1489 -587 1613 -553
rect 1439 -603 1613 -587
rect 2488 -553 2542 -537
rect 2488 -587 2498 -553
rect 2532 -587 2542 -553
rect 2584 -538 2659 -528
rect 2584 -572 2600 -538
rect 2634 -572 2659 -538
rect 2797 -492 2926 -476
rect 2972 -437 3038 -427
rect 2972 -471 2988 -437
rect 3022 -471 3038 -437
rect 2972 -481 3038 -471
rect 2797 -526 2807 -492
rect 2841 -506 2926 -492
rect 2841 -526 2914 -506
rect 3087 -523 3117 -389
rect 3227 -447 3257 -389
rect 3227 -463 3282 -447
rect 3227 -497 3237 -463
rect 3271 -497 3282 -463
rect 3227 -513 3282 -497
rect 2797 -542 2914 -526
rect 2584 -582 2659 -572
rect 2488 -603 2542 -587
rect 1499 -625 1529 -603
rect 1583 -625 1613 -603
rect 2512 -626 2542 -603
rect 2512 -656 2575 -626
rect 2545 -671 2575 -656
rect 2629 -671 2659 -582
rect 2884 -671 2914 -542
rect 2979 -553 3117 -523
rect 2979 -583 3010 -553
rect 2956 -599 3010 -583
rect 2956 -633 2966 -599
rect 3000 -633 3010 -599
rect 2956 -649 3010 -633
rect 3052 -605 3118 -595
rect 3052 -639 3068 -605
rect 3102 -639 3118 -605
rect 3052 -649 3118 -639
rect 2979 -683 3009 -649
rect 3075 -683 3105 -649
rect 3241 -671 3271 -513
rect 3324 -583 3354 -389
rect 3521 -488 3551 -473
rect 3445 -518 3551 -488
rect 3445 -535 3475 -518
rect 3409 -551 3475 -535
rect 3313 -599 3367 -583
rect 3313 -633 3323 -599
rect 3357 -633 3367 -599
rect 3409 -585 3419 -551
rect 3453 -585 3475 -551
rect 3620 -523 3650 -389
rect 3706 -421 3736 -389
rect 3692 -437 3746 -421
rect 3692 -471 3702 -437
rect 3736 -471 3746 -437
rect 3692 -487 3746 -471
rect 3620 -535 3670 -523
rect 3620 -547 3683 -535
rect 3620 -553 3707 -547
rect 3641 -563 3707 -553
rect 3641 -565 3663 -563
rect 3409 -601 3475 -585
rect 3445 -627 3475 -601
rect 3544 -611 3611 -595
rect 3313 -649 3367 -633
rect 3313 -671 3343 -649
rect 3544 -645 3567 -611
rect 3601 -645 3611 -611
rect 3544 -661 3611 -645
rect 3653 -597 3663 -565
rect 3697 -597 3707 -563
rect 3653 -613 3707 -597
rect 3790 -573 3820 -389
rect 3898 -545 3928 -389
rect 3982 -437 4012 -389
rect 3970 -453 4024 -437
rect 3970 -487 3980 -453
rect 4014 -487 4024 -453
rect 3970 -503 4024 -487
rect 3893 -561 3947 -545
rect 3790 -589 3851 -573
rect 3790 -609 3807 -589
rect 3544 -683 3574 -661
rect 3653 -683 3683 -613
rect 3749 -623 3807 -609
rect 3841 -623 3851 -589
rect 3893 -595 3903 -561
rect 3937 -595 3947 -561
rect 3893 -611 3947 -595
rect 3749 -639 3851 -623
rect 3749 -671 3779 -639
rect 3898 -671 3928 -611
rect 3989 -671 4019 -503
rect 4365 -469 4395 -433
rect 4354 -499 4395 -469
rect 4146 -537 4176 -505
rect 4354 -537 4384 -499
rect 4462 -537 4492 -505
rect 4075 -553 4384 -537
rect 4075 -587 4103 -553
rect 4137 -587 4384 -553
rect 4075 -603 4384 -587
rect 4433 -553 4492 -537
rect 4433 -587 4443 -553
rect 4477 -587 4492 -553
rect 4433 -603 4492 -587
rect 4177 -625 4207 -603
rect 4354 -626 4384 -603
rect 4462 -625 4492 -603
rect 4354 -656 4395 -626
rect 4365 -671 4395 -656
rect 1499 -781 1529 -755
rect 1583 -781 1613 -755
rect 2545 -781 2575 -755
rect 2629 -781 2659 -755
rect 2884 -781 2914 -755
rect 2979 -781 3009 -755
rect 3075 -781 3105 -755
rect 3241 -781 3271 -755
rect 3313 -781 3343 -755
rect 3445 -781 3475 -755
rect 3544 -781 3574 -755
rect 3653 -781 3683 -755
rect 3749 -781 3779 -755
rect 3898 -781 3928 -755
rect 3989 -781 4019 -755
rect 4177 -781 4207 -755
rect 4365 -781 4395 -755
rect 4462 -781 4492 -755
<< polycont >>
rect 32 215 66 249
rect 134 230 168 264
rect 522 331 556 365
rect 341 276 375 310
rect 771 305 805 339
rect 500 169 534 203
rect 602 163 636 197
rect 857 169 891 203
rect 953 217 987 251
rect 1236 331 1270 365
rect 1101 157 1135 191
rect 1197 205 1231 239
rect 1514 315 1548 349
rect 1341 179 1375 213
rect 1437 207 1471 241
rect 1637 215 1671 249
rect 1977 215 2011 249
rect 2498 215 2532 249
rect 2600 230 2634 264
rect 2988 331 3022 365
rect 2807 276 2841 310
rect 3237 305 3271 339
rect 2966 169 3000 203
rect 3068 163 3102 197
rect 3323 169 3357 203
rect 3419 217 3453 251
rect 3702 331 3736 365
rect 3567 157 3601 191
rect 3663 205 3697 239
rect 3980 315 4014 349
rect 3807 179 3841 213
rect 3903 207 3937 241
rect 4103 215 4137 249
rect 4443 215 4477 249
rect 1455 -587 1489 -553
rect 2498 -587 2532 -553
rect 2600 -572 2634 -538
rect 2988 -471 3022 -437
rect 2807 -526 2841 -492
rect 3237 -497 3271 -463
rect 2966 -633 3000 -599
rect 3068 -639 3102 -605
rect 3323 -633 3357 -599
rect 3419 -585 3453 -551
rect 3702 -471 3736 -437
rect 3567 -645 3601 -611
rect 3663 -597 3697 -563
rect 3980 -487 4014 -453
rect 3807 -623 3841 -589
rect 3903 -595 3937 -561
rect 4103 -587 4137 -553
rect 4443 -587 4477 -553
<< locali >>
rect 0 585 2116 597
rect 0 527 29 585
rect 63 527 121 585
rect 155 527 213 585
rect 247 527 305 585
rect 339 527 397 585
rect 431 527 489 585
rect 523 527 581 585
rect 615 527 673 585
rect 707 527 765 585
rect 799 527 857 585
rect 891 527 949 585
rect 983 527 1041 585
rect 1075 527 1133 585
rect 1167 527 1225 585
rect 1259 527 1317 585
rect 1351 527 1409 585
rect 1443 527 1501 585
rect 1535 527 1593 585
rect 1627 527 1685 585
rect 1719 527 1777 585
rect 1811 527 1869 585
rect 1903 527 1961 585
rect 1995 527 2053 585
rect 2087 527 2116 585
rect 2466 585 4582 599
rect 2466 527 2495 585
rect 2529 527 2587 585
rect 2621 527 2679 585
rect 2713 527 2771 585
rect 2805 527 2863 585
rect 2897 527 2955 585
rect 2989 527 3047 585
rect 3081 527 3139 585
rect 3173 527 3231 585
rect 3265 527 3323 585
rect 3357 527 3415 585
rect 3449 527 3507 585
rect 3541 527 3599 585
rect 3633 527 3691 585
rect 3725 527 3783 585
rect 3817 527 3875 585
rect 3909 527 3967 585
rect 4001 527 4059 585
rect 4093 527 4151 585
rect 4185 527 4243 585
rect 4277 527 4335 585
rect 4369 527 4427 585
rect 4461 527 4519 585
rect 4553 527 4582 585
rect 18 477 69 493
rect 18 443 35 477
rect 18 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 18 375 35 409
rect 203 409 237 443
rect 69 375 168 393
rect 18 359 168 375
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 122 264 168 359
rect 122 255 134 264
rect 156 221 168 230
rect 122 161 168 221
rect 18 127 168 161
rect 18 119 69 127
rect 18 85 35 119
rect 203 119 237 357
rect 271 333 336 490
rect 370 485 420 527
rect 370 451 386 485
rect 370 435 420 451
rect 454 477 504 493
rect 454 443 470 477
rect 454 427 504 443
rect 547 483 683 493
rect 547 449 563 483
rect 597 449 683 483
rect 798 475 864 527
rect 991 485 1065 527
rect 547 427 683 449
rect 454 401 488 427
rect 409 367 488 401
rect 522 391 615 393
rect 283 323 375 333
rect 283 289 305 323
rect 339 310 375 323
rect 339 289 341 310
rect 283 276 341 289
rect 283 123 375 276
rect 18 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 409 95 443 367
rect 522 365 581 391
rect 556 357 581 365
rect 556 331 615 357
rect 522 315 615 331
rect 477 255 547 277
rect 477 221 489 255
rect 523 221 547 255
rect 477 203 547 221
rect 477 169 500 203
rect 534 169 547 203
rect 477 153 547 169
rect 581 197 615 315
rect 649 271 683 427
rect 717 459 751 475
rect 798 441 814 475
rect 848 441 864 475
rect 898 459 932 475
rect 717 407 751 425
rect 991 451 1011 485
rect 1045 451 1065 485
rect 991 435 1065 451
rect 1099 477 1133 493
rect 898 407 932 425
rect 717 373 932 407
rect 1099 401 1133 443
rect 1180 484 1354 493
rect 1180 450 1196 484
rect 1230 450 1354 484
rect 1180 425 1354 450
rect 1388 485 1438 527
rect 1422 451 1438 485
rect 1542 485 1686 527
rect 1388 435 1438 451
rect 1472 459 1506 475
rect 1021 367 1133 401
rect 1021 339 1055 367
rect 755 305 771 339
rect 805 305 1055 339
rect 1194 357 1205 391
rect 1239 365 1286 391
rect 1194 333 1236 357
rect 649 251 987 271
rect 649 237 953 251
rect 581 163 602 197
rect 636 163 652 197
rect 581 153 652 163
rect 686 95 720 237
rect 761 187 857 203
rect 795 153 833 187
rect 891 169 919 203
rect 953 201 987 217
rect 867 153 919 169
rect 1021 167 1055 305
rect 203 69 237 85
rect 103 17 169 59
rect 309 55 325 89
rect 359 55 375 89
rect 409 61 458 95
rect 492 61 508 95
rect 549 61 565 95
rect 599 61 720 95
rect 895 93 961 109
rect 309 17 375 55
rect 895 59 911 93
rect 945 59 961 93
rect 895 17 961 59
rect 1003 89 1055 167
rect 1093 331 1236 333
rect 1270 331 1286 365
rect 1320 349 1354 425
rect 1542 451 1558 485
rect 1592 451 1636 485
rect 1670 451 1686 485
rect 1720 477 1801 493
rect 1952 485 1986 527
rect 1472 417 1506 425
rect 1754 443 1801 477
rect 1472 383 1632 417
rect 1093 299 1228 331
rect 1320 315 1514 349
rect 1548 315 1564 349
rect 1093 191 1135 299
rect 1320 297 1354 315
rect 1093 157 1101 191
rect 1093 141 1135 157
rect 1169 255 1239 265
rect 1169 239 1205 255
rect 1169 205 1197 239
rect 1231 205 1239 221
rect 1169 141 1239 205
rect 1273 263 1354 297
rect 1273 107 1307 263
rect 1421 250 1529 281
rect 1598 265 1632 383
rect 1720 409 1801 443
rect 1754 375 1801 409
rect 1720 341 1801 375
rect 1754 307 1801 341
rect 1720 291 1801 307
rect 1598 259 1687 265
rect 1455 241 1529 250
rect 1341 213 1385 229
rect 1375 179 1385 213
rect 1421 207 1437 216
rect 1471 207 1529 241
rect 1341 173 1385 179
rect 1481 187 1529 207
rect 1341 139 1447 173
rect 1117 93 1307 107
rect 1003 55 1023 89
rect 1057 55 1073 89
rect 1117 59 1133 93
rect 1167 59 1307 93
rect 1117 51 1307 59
rect 1341 89 1379 105
rect 1341 55 1345 89
rect 1413 93 1447 139
rect 1515 153 1529 187
rect 1481 127 1529 153
rect 1563 249 1687 259
rect 1563 215 1637 249
rect 1671 215 1687 249
rect 1563 199 1687 215
rect 1735 253 1801 291
rect 1735 218 1754 253
rect 1788 218 1801 253
rect 1563 164 1628 199
rect 1735 165 1801 218
rect 1563 109 1627 164
rect 1413 75 1563 93
rect 1597 75 1627 109
rect 1413 59 1627 75
rect 1667 132 1701 154
rect 1341 17 1379 55
rect 1667 17 1701 98
rect 1735 131 1751 165
rect 1785 131 1801 165
rect 1735 97 1801 131
rect 1735 63 1751 97
rect 1785 63 1801 97
rect 1839 451 1855 485
rect 1889 451 1905 485
rect 1839 417 1905 451
rect 1839 383 1855 417
rect 1889 383 1905 417
rect 1839 265 1905 383
rect 2484 477 2535 493
rect 1952 417 1986 451
rect 1952 349 1986 383
rect 1952 299 1986 315
rect 2036 449 2087 465
rect 2070 415 2087 449
rect 2036 381 2087 415
rect 2070 347 2087 381
rect 2484 443 2501 477
rect 2484 409 2535 443
rect 2569 461 2635 527
rect 2569 427 2585 461
rect 2619 427 2635 461
rect 2669 477 2703 493
rect 2484 375 2501 409
rect 2669 409 2703 443
rect 2535 375 2634 393
rect 2484 359 2634 375
rect 2036 289 2087 347
rect 1839 249 2011 265
rect 1839 215 1977 249
rect 1839 199 2011 215
rect 2045 254 2087 289
rect 2045 220 2049 254
rect 2083 220 2087 254
rect 1839 119 1889 199
rect 2045 159 2087 220
rect 2484 255 2554 325
rect 2484 221 2496 255
rect 2530 249 2554 255
rect 2484 215 2498 221
rect 2532 215 2554 249
rect 2484 195 2554 215
rect 2588 264 2634 359
rect 2588 255 2600 264
rect 2622 221 2634 230
rect 2588 161 2634 221
rect 2036 143 2087 159
rect 1839 85 1855 119
rect 1839 69 1889 85
rect 1952 113 1986 136
rect 1735 55 1801 63
rect 1952 17 1986 79
rect 2070 109 2087 143
rect 2036 53 2087 109
rect 2484 127 2634 161
rect 2484 119 2535 127
rect 2484 85 2501 119
rect 2669 119 2703 357
rect 2737 333 2802 490
rect 2836 485 2886 527
rect 2836 451 2852 485
rect 2836 435 2886 451
rect 2920 477 2970 493
rect 2920 443 2936 477
rect 2920 427 2970 443
rect 3013 483 3149 493
rect 3013 449 3029 483
rect 3063 449 3149 483
rect 3264 475 3330 527
rect 3457 485 3531 527
rect 3013 427 3149 449
rect 2920 401 2954 427
rect 2875 367 2954 401
rect 2988 391 3081 393
rect 2749 323 2841 333
rect 2749 289 2771 323
rect 2805 310 2841 323
rect 2805 289 2807 310
rect 2749 276 2807 289
rect 2749 123 2841 276
rect 2484 69 2535 85
rect 2569 59 2585 93
rect 2619 59 2635 93
rect 2875 95 2909 367
rect 2988 365 3047 391
rect 3022 357 3047 365
rect 3022 331 3081 357
rect 2988 315 3081 331
rect 2943 255 3013 277
rect 2943 221 2955 255
rect 2989 221 3013 255
rect 2943 203 3013 221
rect 2943 169 2966 203
rect 3000 169 3013 203
rect 2943 153 3013 169
rect 3047 197 3081 315
rect 3115 271 3149 427
rect 3183 459 3217 475
rect 3264 441 3280 475
rect 3314 441 3330 475
rect 3364 459 3398 475
rect 3183 407 3217 425
rect 3457 451 3477 485
rect 3511 451 3531 485
rect 3457 435 3531 451
rect 3565 477 3599 493
rect 3364 407 3398 425
rect 3183 373 3398 407
rect 3565 401 3599 443
rect 3646 484 3820 493
rect 3646 450 3662 484
rect 3696 450 3820 484
rect 3646 425 3820 450
rect 3854 485 3904 527
rect 3888 451 3904 485
rect 4008 485 4152 527
rect 3854 435 3904 451
rect 3938 459 3972 475
rect 3487 367 3599 401
rect 3487 339 3521 367
rect 3221 305 3237 339
rect 3271 305 3521 339
rect 3660 357 3671 391
rect 3705 365 3752 391
rect 3660 333 3702 357
rect 3115 251 3453 271
rect 3115 237 3419 251
rect 3047 163 3068 197
rect 3102 163 3118 197
rect 3047 153 3118 163
rect 3152 95 3186 237
rect 3227 187 3323 203
rect 3261 153 3299 187
rect 3357 169 3385 203
rect 3419 201 3453 217
rect 3333 153 3385 169
rect 3487 167 3521 305
rect 2669 69 2703 85
rect 2569 17 2635 59
rect 2775 55 2791 89
rect 2825 55 2841 89
rect 2875 61 2924 95
rect 2958 61 2974 95
rect 3015 61 3031 95
rect 3065 61 3186 95
rect 3361 93 3427 109
rect 2775 17 2841 55
rect 3361 59 3377 93
rect 3411 59 3427 93
rect 3361 17 3427 59
rect 3469 89 3521 167
rect 3559 331 3702 333
rect 3736 331 3752 365
rect 3786 349 3820 425
rect 4008 451 4024 485
rect 4058 451 4102 485
rect 4136 451 4152 485
rect 4186 477 4267 493
rect 4418 485 4452 527
rect 3938 417 3972 425
rect 4220 443 4267 477
rect 3938 383 4098 417
rect 3559 299 3694 331
rect 3786 315 3980 349
rect 4014 315 4030 349
rect 3559 191 3601 299
rect 3786 297 3820 315
rect 3559 157 3567 191
rect 3559 141 3601 157
rect 3635 255 3705 265
rect 3635 239 3671 255
rect 3635 205 3663 239
rect 3697 205 3705 221
rect 3635 141 3705 205
rect 3739 263 3820 297
rect 3739 107 3773 263
rect 3887 250 3995 281
rect 4064 265 4098 383
rect 4186 409 4267 443
rect 4220 375 4267 409
rect 4186 341 4267 375
rect 4220 307 4267 341
rect 4186 291 4267 307
rect 4064 259 4153 265
rect 3921 241 3995 250
rect 3807 213 3851 229
rect 3841 179 3851 213
rect 3887 207 3903 216
rect 3937 207 3995 241
rect 3807 173 3851 179
rect 3947 187 3995 207
rect 3807 139 3913 173
rect 3583 93 3773 107
rect 3469 55 3489 89
rect 3523 55 3539 89
rect 3583 59 3599 93
rect 3633 59 3773 93
rect 3583 51 3773 59
rect 3807 89 3845 105
rect 3807 55 3811 89
rect 3879 93 3913 139
rect 3981 153 3995 187
rect 3947 127 3995 153
rect 4029 249 4153 259
rect 4029 215 4103 249
rect 4137 215 4153 249
rect 4029 199 4153 215
rect 4029 164 4094 199
rect 4201 165 4267 291
rect 4029 109 4093 164
rect 3879 75 4029 93
rect 4063 75 4093 109
rect 3879 59 4093 75
rect 4133 132 4167 154
rect 3807 17 3845 55
rect 4133 17 4167 98
rect 4201 131 4217 165
rect 4251 131 4267 165
rect 4201 97 4267 131
rect 4201 63 4217 97
rect 4251 63 4267 97
rect 4305 451 4321 485
rect 4355 451 4371 485
rect 4305 417 4371 451
rect 4305 383 4321 417
rect 4355 383 4371 417
rect 4305 265 4371 383
rect 4418 417 4452 451
rect 4418 349 4452 383
rect 4418 299 4452 315
rect 4502 449 4553 465
rect 4536 415 4553 449
rect 4502 381 4553 415
rect 4536 347 4553 381
rect 4502 289 4553 347
rect 4305 249 4477 265
rect 4305 215 4443 249
rect 4305 199 4477 215
rect 4511 255 4553 289
rect 4511 221 4517 255
rect 4551 221 4553 255
rect 4305 119 4355 199
rect 4511 159 4553 221
rect 4502 143 4553 159
rect 4305 85 4321 119
rect 4305 69 4355 85
rect 4418 113 4452 136
rect 4201 55 4267 63
rect 4418 17 4452 79
rect 4536 109 4553 143
rect 4502 53 4553 109
rect 0 -45 29 17
rect 63 -45 121 17
rect 155 -45 213 17
rect 247 -45 305 17
rect 339 -45 397 17
rect 431 -45 489 17
rect 523 -45 581 17
rect 615 -45 673 17
rect 707 -45 765 17
rect 799 -45 857 17
rect 891 -45 949 17
rect 983 -45 1041 17
rect 1075 -45 1133 17
rect 1167 -45 1225 17
rect 1259 -45 1317 17
rect 1351 -45 1409 17
rect 1443 -45 1501 17
rect 1535 -45 1593 17
rect 1627 -45 1685 17
rect 1719 -45 1777 17
rect 1811 -45 1869 17
rect 1903 -45 1961 17
rect 1995 -45 2053 17
rect 2087 -45 2116 17
rect 0 -88 2116 -45
rect 2466 -44 2495 17
rect 2529 -44 2587 17
rect 2621 -44 2679 17
rect 2713 -44 2771 17
rect 2805 -44 2863 17
rect 2897 -44 2955 17
rect 2989 -44 3047 17
rect 3081 -44 3139 17
rect 3173 -44 3231 17
rect 3265 -44 3323 17
rect 3357 -44 3415 17
rect 3449 -44 3507 17
rect 3541 -44 3599 17
rect 3633 -44 3691 17
rect 3725 -44 3783 17
rect 3817 -44 3875 17
rect 3909 -44 3967 17
rect 4001 -44 4059 17
rect 4093 -44 4151 17
rect 4185 -44 4243 17
rect 4277 -44 4335 17
rect 4369 -44 4427 17
rect 4461 -44 4519 17
rect 4553 -44 4582 17
rect 2466 -47 4582 -44
rect 1418 -217 1694 -213
rect 1418 -275 1447 -217
rect 1481 -275 1539 -217
rect 1573 -275 1631 -217
rect 1665 -275 1694 -217
rect 2466 -275 2495 -216
rect 2529 -275 2587 -216
rect 2621 -275 2679 -216
rect 2713 -275 2771 -216
rect 2805 -275 2863 -216
rect 2897 -275 2955 -216
rect 2989 -275 3047 -216
rect 3081 -275 3139 -216
rect 3173 -275 3231 -216
rect 3265 -275 3323 -216
rect 3357 -275 3415 -216
rect 3449 -275 3507 -216
rect 3541 -275 3599 -216
rect 3633 -275 3691 -216
rect 3725 -275 3783 -216
rect 3817 -275 3875 -216
rect 3909 -275 3967 -216
rect 4001 -275 4059 -216
rect 4093 -275 4151 -216
rect 4185 -275 4243 -216
rect 4277 -275 4335 -216
rect 4369 -275 4427 -216
rect 4461 -275 4519 -216
rect 4553 -275 4582 -216
rect 1443 -317 1489 -275
rect 1443 -351 1455 -317
rect 1443 -385 1489 -351
rect 1443 -419 1455 -385
rect 1443 -453 1489 -419
rect 1443 -487 1455 -453
rect 1443 -503 1489 -487
rect 1523 -317 1589 -309
rect 1523 -351 1539 -317
rect 1573 -351 1589 -317
rect 1523 -385 1589 -351
rect 1523 -419 1539 -385
rect 1573 -419 1589 -385
rect 1523 -453 1589 -419
rect 1523 -487 1539 -453
rect 1573 -487 1589 -453
rect 1523 -505 1589 -487
rect 1623 -317 1665 -275
rect 1657 -351 1665 -317
rect 1623 -385 1665 -351
rect 1657 -419 1665 -385
rect 1623 -453 1665 -419
rect 2484 -325 2535 -309
rect 2484 -359 2501 -325
rect 2484 -393 2535 -359
rect 2569 -341 2635 -275
rect 2569 -375 2585 -341
rect 2619 -375 2635 -341
rect 2669 -325 2703 -309
rect 2484 -427 2501 -393
rect 2669 -393 2703 -359
rect 2535 -427 2634 -409
rect 2484 -443 2634 -427
rect 1657 -487 1665 -453
rect 1623 -503 1665 -487
rect 1439 -547 1505 -537
rect 1439 -581 1447 -547
rect 1481 -553 1505 -547
rect 1439 -587 1455 -581
rect 1489 -587 1505 -553
rect 1539 -577 1589 -505
rect 1573 -611 1589 -577
rect 2484 -513 2554 -477
rect 2484 -547 2496 -513
rect 2531 -547 2554 -513
rect 2484 -553 2554 -547
rect 2484 -587 2498 -553
rect 2532 -587 2554 -553
rect 2484 -607 2554 -587
rect 2588 -538 2634 -443
rect 2588 -547 2600 -538
rect 2622 -581 2634 -572
rect 1443 -637 1489 -621
rect 1539 -625 1589 -611
rect 1443 -671 1455 -637
rect 1443 -709 1489 -671
rect 1443 -743 1455 -709
rect 1443 -785 1489 -743
rect 1523 -637 1589 -625
rect 1523 -671 1539 -637
rect 1573 -671 1589 -637
rect 1523 -709 1589 -671
rect 1523 -743 1539 -709
rect 1573 -743 1589 -709
rect 1523 -751 1589 -743
rect 1623 -637 1665 -621
rect 1657 -671 1665 -637
rect 2588 -641 2634 -581
rect 1623 -709 1665 -671
rect 1657 -743 1665 -709
rect 2484 -675 2634 -641
rect 2484 -683 2535 -675
rect 2484 -717 2501 -683
rect 2669 -683 2703 -445
rect 2737 -469 2802 -312
rect 2836 -317 2886 -275
rect 2836 -351 2852 -317
rect 2836 -367 2886 -351
rect 2920 -325 2970 -309
rect 2920 -359 2936 -325
rect 2920 -375 2970 -359
rect 3013 -319 3149 -309
rect 3013 -353 3029 -319
rect 3063 -353 3149 -319
rect 3264 -327 3330 -275
rect 3457 -317 3531 -275
rect 3013 -375 3149 -353
rect 2920 -401 2954 -375
rect 2875 -435 2954 -401
rect 2988 -411 3081 -409
rect 2749 -492 2841 -469
rect 2749 -509 2807 -492
rect 2749 -543 2771 -509
rect 2805 -526 2807 -509
rect 2805 -543 2841 -526
rect 2749 -679 2841 -543
rect 2484 -733 2535 -717
rect 1623 -785 1665 -743
rect 2569 -743 2585 -709
rect 2619 -743 2635 -709
rect 2875 -707 2909 -435
rect 2988 -437 3047 -411
rect 3022 -445 3047 -437
rect 3022 -471 3081 -445
rect 2988 -487 3081 -471
rect 2943 -547 3013 -525
rect 2943 -581 2955 -547
rect 2989 -581 3013 -547
rect 2943 -599 3013 -581
rect 2943 -633 2966 -599
rect 3000 -633 3013 -599
rect 2943 -649 3013 -633
rect 3047 -605 3081 -487
rect 3115 -531 3149 -375
rect 3183 -343 3217 -327
rect 3264 -361 3280 -327
rect 3314 -361 3330 -327
rect 3364 -343 3398 -327
rect 3183 -395 3217 -377
rect 3457 -351 3477 -317
rect 3511 -351 3531 -317
rect 3457 -367 3531 -351
rect 3565 -325 3599 -309
rect 3364 -395 3398 -377
rect 3183 -429 3398 -395
rect 3565 -401 3599 -359
rect 3646 -318 3820 -309
rect 3646 -352 3662 -318
rect 3696 -352 3820 -318
rect 3646 -377 3820 -352
rect 3854 -317 3904 -275
rect 3888 -351 3904 -317
rect 4008 -317 4152 -275
rect 3854 -367 3904 -351
rect 3938 -343 3972 -327
rect 3487 -435 3599 -401
rect 3487 -463 3521 -435
rect 3221 -497 3237 -463
rect 3271 -497 3521 -463
rect 3660 -445 3671 -411
rect 3705 -437 3752 -411
rect 3660 -469 3702 -445
rect 3115 -551 3453 -531
rect 3115 -565 3419 -551
rect 3047 -639 3068 -605
rect 3102 -639 3118 -605
rect 3047 -649 3118 -639
rect 3152 -707 3186 -565
rect 3227 -615 3323 -599
rect 3261 -649 3299 -615
rect 3357 -633 3385 -599
rect 3419 -601 3453 -585
rect 3333 -649 3385 -633
rect 3487 -635 3521 -497
rect 2669 -733 2703 -717
rect 2569 -785 2635 -743
rect 2775 -747 2791 -713
rect 2825 -747 2841 -713
rect 2875 -741 2924 -707
rect 2958 -741 2974 -707
rect 3015 -741 3031 -707
rect 3065 -741 3186 -707
rect 3361 -709 3427 -693
rect 2775 -785 2841 -747
rect 3361 -743 3377 -709
rect 3411 -743 3427 -709
rect 3361 -785 3427 -743
rect 3469 -713 3521 -635
rect 3559 -471 3702 -469
rect 3736 -471 3752 -437
rect 3786 -453 3820 -377
rect 4008 -351 4024 -317
rect 4058 -351 4102 -317
rect 4136 -351 4152 -317
rect 4186 -325 4267 -309
rect 4418 -317 4452 -275
rect 3938 -385 3972 -377
rect 4220 -359 4267 -325
rect 3938 -419 4098 -385
rect 3559 -503 3694 -471
rect 3786 -487 3980 -453
rect 4014 -487 4030 -453
rect 3559 -611 3601 -503
rect 3786 -505 3820 -487
rect 3559 -645 3567 -611
rect 3559 -661 3601 -645
rect 3635 -547 3705 -537
rect 3635 -563 3671 -547
rect 3635 -597 3663 -563
rect 3697 -597 3705 -581
rect 3635 -661 3705 -597
rect 3739 -539 3820 -505
rect 3739 -695 3773 -539
rect 3887 -552 3995 -521
rect 4064 -537 4098 -419
rect 4186 -393 4267 -359
rect 4220 -427 4267 -393
rect 4186 -461 4267 -427
rect 4220 -495 4267 -461
rect 4186 -511 4267 -495
rect 4064 -543 4153 -537
rect 3921 -561 3995 -552
rect 3807 -589 3851 -573
rect 3841 -623 3851 -589
rect 3887 -595 3903 -586
rect 3937 -595 3995 -561
rect 3807 -629 3851 -623
rect 3947 -615 3995 -595
rect 3807 -663 3913 -629
rect 3583 -709 3773 -695
rect 3469 -747 3489 -713
rect 3523 -747 3539 -713
rect 3583 -743 3599 -709
rect 3633 -743 3773 -709
rect 3583 -751 3773 -743
rect 3807 -713 3845 -697
rect 3807 -747 3811 -713
rect 3879 -709 3913 -663
rect 3981 -649 3995 -615
rect 3947 -675 3995 -649
rect 4029 -553 4153 -543
rect 4029 -587 4103 -553
rect 4137 -587 4153 -553
rect 4029 -603 4153 -587
rect 4029 -638 4094 -603
rect 4201 -637 4267 -511
rect 4029 -693 4093 -638
rect 3879 -727 4029 -709
rect 4063 -727 4093 -693
rect 3879 -743 4093 -727
rect 4133 -670 4167 -648
rect 3807 -785 3845 -747
rect 4133 -785 4167 -704
rect 4201 -671 4217 -637
rect 4251 -671 4267 -637
rect 4201 -705 4267 -671
rect 4201 -739 4217 -705
rect 4251 -739 4267 -705
rect 4305 -351 4321 -317
rect 4355 -351 4371 -317
rect 4305 -385 4371 -351
rect 4305 -419 4321 -385
rect 4355 -419 4371 -385
rect 4305 -537 4371 -419
rect 4418 -385 4452 -351
rect 4418 -453 4452 -419
rect 4418 -503 4452 -487
rect 4502 -353 4553 -337
rect 4536 -387 4553 -353
rect 4502 -421 4553 -387
rect 4536 -455 4553 -421
rect 4502 -513 4553 -455
rect 4305 -553 4477 -537
rect 4305 -587 4443 -553
rect 4305 -603 4477 -587
rect 4511 -578 4553 -513
rect 4305 -683 4355 -603
rect 4511 -612 4515 -578
rect 4549 -612 4553 -578
rect 4511 -643 4553 -612
rect 4502 -659 4553 -643
rect 4305 -717 4321 -683
rect 4305 -733 4355 -717
rect 4418 -689 4452 -666
rect 4201 -747 4267 -739
rect 4418 -785 4452 -723
rect 4536 -693 4553 -659
rect 4502 -749 4553 -693
rect 1418 -845 1447 -785
rect 1481 -845 1539 -785
rect 1573 -845 1631 -785
rect 1665 -845 1694 -785
rect 1418 -847 1694 -845
rect 2466 -847 2495 -785
rect 2529 -847 2587 -785
rect 2621 -847 2679 -785
rect 2713 -847 2771 -785
rect 2805 -847 2863 -785
rect 2897 -847 2955 -785
rect 2989 -847 3047 -785
rect 3081 -847 3139 -785
rect 3173 -847 3231 -785
rect 3265 -847 3323 -785
rect 3357 -847 3415 -785
rect 3449 -847 3507 -785
rect 3541 -847 3599 -785
rect 3633 -847 3691 -785
rect 3725 -847 3783 -785
rect 3817 -847 3875 -785
rect 3909 -847 3967 -785
rect 4001 -847 4059 -785
rect 4093 -847 4151 -785
rect 4185 -847 4243 -785
rect 4277 -847 4335 -785
rect 4369 -847 4427 -785
rect 4461 -847 4519 -785
rect 4553 -847 4582 -785
rect 2466 -848 4582 -847
<< viali >>
rect 29 551 63 561
rect 29 527 63 551
rect 121 551 155 561
rect 121 527 155 551
rect 213 551 247 561
rect 213 527 247 551
rect 305 551 339 561
rect 305 527 339 551
rect 397 551 431 561
rect 397 527 431 551
rect 489 551 523 561
rect 489 527 523 551
rect 581 551 615 561
rect 581 527 615 551
rect 673 551 707 561
rect 673 527 707 551
rect 765 551 799 561
rect 765 527 799 551
rect 857 551 891 561
rect 857 527 891 551
rect 949 551 983 561
rect 949 527 983 551
rect 1041 551 1075 561
rect 1041 527 1075 551
rect 1133 551 1167 561
rect 1133 527 1167 551
rect 1225 551 1259 561
rect 1225 527 1259 551
rect 1317 551 1351 561
rect 1317 527 1351 551
rect 1409 551 1443 561
rect 1409 527 1443 551
rect 1501 551 1535 561
rect 1501 527 1535 551
rect 1593 551 1627 561
rect 1593 527 1627 551
rect 1685 551 1719 561
rect 1685 527 1719 551
rect 1777 551 1811 561
rect 1777 527 1811 551
rect 1869 551 1903 561
rect 1869 527 1903 551
rect 1961 551 1995 561
rect 1961 527 1995 551
rect 2053 551 2087 561
rect 2053 527 2087 551
rect 2495 551 2529 561
rect 2495 527 2529 551
rect 2587 551 2621 561
rect 2587 527 2621 551
rect 2679 551 2713 561
rect 2679 527 2713 551
rect 2771 551 2805 561
rect 2771 527 2805 551
rect 2863 551 2897 561
rect 2863 527 2897 551
rect 2955 551 2989 561
rect 2955 527 2989 551
rect 3047 551 3081 561
rect 3047 527 3081 551
rect 3139 551 3173 561
rect 3139 527 3173 551
rect 3231 551 3265 561
rect 3231 527 3265 551
rect 3323 551 3357 561
rect 3323 527 3357 551
rect 3415 551 3449 561
rect 3415 527 3449 551
rect 3507 551 3541 561
rect 3507 527 3541 551
rect 3599 551 3633 561
rect 3599 527 3633 551
rect 3691 551 3725 561
rect 3691 527 3725 551
rect 3783 551 3817 561
rect 3783 527 3817 551
rect 3875 551 3909 561
rect 3875 527 3909 551
rect 3967 551 4001 561
rect 3967 527 4001 551
rect 4059 551 4093 561
rect 4059 527 4093 551
rect 4151 551 4185 561
rect 4151 527 4185 551
rect 4243 551 4277 561
rect 4243 527 4277 551
rect 4335 551 4369 561
rect 4335 527 4369 551
rect 4427 551 4461 561
rect 4427 527 4461 551
rect 4519 551 4553 561
rect 4519 527 4553 551
rect 122 230 134 255
rect 134 230 156 255
rect 122 221 156 230
rect 203 375 237 391
rect 203 357 237 375
rect 305 289 339 323
rect 581 357 615 391
rect 489 221 523 255
rect 1205 365 1239 391
rect 1205 357 1236 365
rect 1236 357 1239 365
rect 761 153 795 187
rect 833 169 857 187
rect 857 169 867 187
rect 833 153 867 169
rect 1205 239 1239 255
rect 1205 221 1231 239
rect 1231 221 1239 239
rect 1421 241 1455 250
rect 1421 216 1437 241
rect 1437 216 1455 241
rect 1481 153 1515 187
rect 1754 218 1788 253
rect 2049 220 2083 254
rect 2496 249 2530 255
rect 2496 221 2498 249
rect 2498 221 2530 249
rect 2588 230 2600 255
rect 2600 230 2622 255
rect 2588 221 2622 230
rect 2669 375 2703 391
rect 2669 357 2703 375
rect 2771 289 2805 323
rect 3047 357 3081 391
rect 2955 221 2989 255
rect 3671 365 3705 391
rect 3671 357 3702 365
rect 3702 357 3705 365
rect 3227 153 3261 187
rect 3299 169 3323 187
rect 3323 169 3333 187
rect 3299 153 3333 169
rect 3671 239 3705 255
rect 3671 221 3697 239
rect 3697 221 3705 239
rect 3887 241 3921 250
rect 3887 216 3903 241
rect 3903 216 3921 241
rect 3947 153 3981 187
rect 4517 221 4551 255
rect 29 -11 63 17
rect 29 -17 63 -11
rect 121 -11 155 17
rect 121 -17 155 -11
rect 213 -11 247 17
rect 213 -17 247 -11
rect 305 -11 339 17
rect 305 -17 339 -11
rect 397 -11 431 17
rect 397 -17 431 -11
rect 489 -11 523 17
rect 489 -17 523 -11
rect 581 -11 615 17
rect 581 -17 615 -11
rect 673 -11 707 17
rect 673 -17 707 -11
rect 765 -11 799 17
rect 765 -17 799 -11
rect 857 -11 891 17
rect 857 -17 891 -11
rect 949 -11 983 17
rect 949 -17 983 -11
rect 1041 -11 1075 17
rect 1041 -17 1075 -11
rect 1133 -11 1167 17
rect 1133 -17 1167 -11
rect 1225 -11 1259 17
rect 1225 -17 1259 -11
rect 1317 -11 1351 17
rect 1317 -17 1351 -11
rect 1409 -11 1443 17
rect 1409 -17 1443 -11
rect 1501 -11 1535 17
rect 1501 -17 1535 -11
rect 1593 -11 1627 17
rect 1593 -17 1627 -11
rect 1685 -11 1719 17
rect 1685 -17 1719 -11
rect 1777 -11 1811 17
rect 1777 -17 1811 -11
rect 1869 -11 1903 17
rect 1869 -17 1903 -11
rect 1961 -11 1995 17
rect 1961 -17 1995 -11
rect 2053 -11 2087 17
rect 2053 -17 2087 -11
rect 2495 -10 2529 17
rect 2495 -17 2529 -10
rect 2587 -10 2621 17
rect 2587 -17 2621 -10
rect 2679 -10 2713 17
rect 2679 -17 2713 -10
rect 2771 -10 2805 17
rect 2771 -17 2805 -10
rect 2863 -10 2897 17
rect 2863 -17 2897 -10
rect 2955 -10 2989 17
rect 2955 -17 2989 -10
rect 3047 -10 3081 17
rect 3047 -17 3081 -10
rect 3139 -10 3173 17
rect 3139 -17 3173 -10
rect 3231 -10 3265 17
rect 3231 -17 3265 -10
rect 3323 -10 3357 17
rect 3323 -17 3357 -10
rect 3415 -10 3449 17
rect 3415 -17 3449 -10
rect 3507 -10 3541 17
rect 3507 -17 3541 -10
rect 3599 -10 3633 17
rect 3599 -17 3633 -10
rect 3691 -10 3725 17
rect 3691 -17 3725 -10
rect 3783 -10 3817 17
rect 3783 -17 3817 -10
rect 3875 -10 3909 17
rect 3875 -17 3909 -10
rect 3967 -10 4001 17
rect 3967 -17 4001 -10
rect 4059 -10 4093 17
rect 4059 -17 4093 -10
rect 4151 -10 4185 17
rect 4151 -17 4185 -10
rect 4243 -10 4277 17
rect 4243 -17 4277 -10
rect 4335 -10 4369 17
rect 4335 -17 4369 -10
rect 4427 -10 4461 17
rect 4427 -17 4461 -10
rect 4519 -10 4553 17
rect 4519 -17 4553 -10
rect 1447 -251 1481 -241
rect 1447 -275 1481 -251
rect 1539 -251 1573 -241
rect 1539 -275 1573 -251
rect 1631 -251 1665 -241
rect 1631 -275 1665 -251
rect 2495 -250 2529 -241
rect 2495 -275 2529 -250
rect 2587 -250 2621 -241
rect 2587 -275 2621 -250
rect 2679 -250 2713 -241
rect 2679 -275 2713 -250
rect 2771 -250 2805 -241
rect 2771 -275 2805 -250
rect 2863 -250 2897 -241
rect 2863 -275 2897 -250
rect 2955 -250 2989 -241
rect 2955 -275 2989 -250
rect 3047 -250 3081 -241
rect 3047 -275 3081 -250
rect 3139 -250 3173 -241
rect 3139 -275 3173 -250
rect 3231 -250 3265 -241
rect 3231 -275 3265 -250
rect 3323 -250 3357 -241
rect 3323 -275 3357 -250
rect 3415 -250 3449 -241
rect 3415 -275 3449 -250
rect 3507 -250 3541 -241
rect 3507 -275 3541 -250
rect 3599 -250 3633 -241
rect 3599 -275 3633 -250
rect 3691 -250 3725 -241
rect 3691 -275 3725 -250
rect 3783 -250 3817 -241
rect 3783 -275 3817 -250
rect 3875 -250 3909 -241
rect 3875 -275 3909 -250
rect 3967 -250 4001 -241
rect 3967 -275 4001 -250
rect 4059 -250 4093 -241
rect 4059 -275 4093 -250
rect 4151 -250 4185 -241
rect 4151 -275 4185 -250
rect 4243 -250 4277 -241
rect 4243 -275 4277 -250
rect 4335 -250 4369 -241
rect 4335 -275 4369 -250
rect 4427 -250 4461 -241
rect 4427 -275 4461 -250
rect 4519 -250 4553 -241
rect 4519 -275 4553 -250
rect 1447 -553 1481 -547
rect 1447 -581 1455 -553
rect 1455 -581 1481 -553
rect 1539 -611 1573 -577
rect 2496 -547 2531 -513
rect 2588 -572 2600 -547
rect 2600 -572 2622 -547
rect 2588 -581 2622 -572
rect 2669 -427 2703 -411
rect 2669 -445 2703 -427
rect 2771 -543 2805 -509
rect 3047 -445 3081 -411
rect 2955 -581 2989 -547
rect 3671 -437 3705 -411
rect 3671 -445 3702 -437
rect 3702 -445 3705 -437
rect 3227 -649 3261 -615
rect 3299 -633 3323 -615
rect 3323 -633 3333 -615
rect 3299 -649 3333 -633
rect 3671 -563 3705 -547
rect 3671 -581 3697 -563
rect 3697 -581 3705 -563
rect 3887 -561 3921 -552
rect 3887 -586 3903 -561
rect 3903 -586 3921 -561
rect 3947 -649 3981 -615
rect 4515 -612 4549 -578
rect 1447 -811 1481 -785
rect 1447 -819 1481 -811
rect 1539 -811 1573 -785
rect 1539 -819 1573 -811
rect 1631 -811 1665 -785
rect 1631 -819 1665 -811
rect 2495 -813 2529 -785
rect 2495 -819 2529 -813
rect 2587 -813 2621 -785
rect 2587 -819 2621 -813
rect 2679 -813 2713 -785
rect 2679 -819 2713 -813
rect 2771 -813 2805 -785
rect 2771 -819 2805 -813
rect 2863 -813 2897 -785
rect 2863 -819 2897 -813
rect 2955 -813 2989 -785
rect 2955 -819 2989 -813
rect 3047 -813 3081 -785
rect 3047 -819 3081 -813
rect 3139 -813 3173 -785
rect 3139 -819 3173 -813
rect 3231 -813 3265 -785
rect 3231 -819 3265 -813
rect 3323 -813 3357 -785
rect 3323 -819 3357 -813
rect 3415 -813 3449 -785
rect 3415 -819 3449 -813
rect 3507 -813 3541 -785
rect 3507 -819 3541 -813
rect 3599 -813 3633 -785
rect 3599 -819 3633 -813
rect 3691 -813 3725 -785
rect 3691 -819 3725 -813
rect 3783 -813 3817 -785
rect 3783 -819 3817 -813
rect 3875 -813 3909 -785
rect 3875 -819 3909 -813
rect 3967 -813 4001 -785
rect 3967 -819 4001 -813
rect 4059 -813 4093 -785
rect 4059 -819 4093 -813
rect 4151 -813 4185 -785
rect 4151 -819 4185 -813
rect 4243 -813 4277 -785
rect 4243 -819 4277 -813
rect 4335 -813 4369 -785
rect 4335 -819 4369 -813
rect 4427 -813 4461 -785
rect 4427 -819 4461 -813
rect 4519 -813 4553 -785
rect 4519 -819 4553 -813
<< metal1 >>
rect 291 672 2223 715
rect 4674 714 4713 715
rect 291 660 2156 672
rect 291 627 355 660
rect 0 561 2116 627
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 496 2116 527
rect 191 391 249 397
rect 191 357 203 391
rect 237 388 249 391
rect 291 388 355 496
rect 569 391 627 397
rect 569 388 581 391
rect 237 360 581 388
rect 237 357 249 360
rect 191 351 249 357
rect 291 335 355 360
rect 569 357 581 360
rect 615 388 627 391
rect 1193 391 1251 397
rect 1193 388 1205 391
rect 615 360 1205 388
rect 615 357 627 360
rect 569 351 627 357
rect 1193 357 1205 360
rect 1239 357 1251 391
rect 1193 351 1251 357
rect 291 283 297 335
rect 349 283 355 335
rect 291 280 355 283
rect 1726 263 1812 285
rect 2185 268 2221 672
rect 2757 664 4713 714
rect 2757 627 2822 664
rect 2466 561 4582 627
rect 2466 527 2495 561
rect 2529 527 2587 561
rect 2621 527 2679 561
rect 2713 527 2771 561
rect 2805 527 2863 561
rect 2897 527 2955 561
rect 2989 527 3047 561
rect 3081 527 3139 561
rect 3173 527 3231 561
rect 3265 527 3323 561
rect 3357 527 3415 561
rect 3449 527 3507 561
rect 3541 527 3599 561
rect 3633 527 3691 561
rect 3725 527 3783 561
rect 3817 527 3875 561
rect 3909 527 3967 561
rect 4001 527 4059 561
rect 4093 527 4151 561
rect 4185 527 4243 561
rect 4277 527 4335 561
rect 4369 527 4427 561
rect 4461 527 4519 561
rect 4553 527 4582 561
rect 2466 496 4582 527
rect 2657 391 2715 397
rect 2657 357 2669 391
rect 2703 388 2715 391
rect 2757 388 2822 496
rect 3035 391 3093 397
rect 3035 388 3047 391
rect 2703 360 3047 388
rect 2703 357 2715 360
rect 2657 351 2715 357
rect 2757 336 2822 360
rect 3035 357 3047 360
rect 3081 388 3093 391
rect 3659 391 3717 397
rect 3659 388 3671 391
rect 3081 360 3671 388
rect 3081 357 3093 360
rect 3035 351 3093 357
rect 3659 357 3671 360
rect 3705 357 3717 391
rect 3659 351 3717 357
rect 2757 284 2763 336
rect 2815 284 2822 336
rect 2757 280 2822 284
rect 110 255 168 261
rect 110 221 122 255
rect 156 252 168 255
rect 477 255 535 261
rect 477 252 489 255
rect 156 224 489 252
rect 156 221 168 224
rect 110 215 168 221
rect 477 221 489 224
rect 523 252 535 255
rect 1193 255 1251 261
rect 1193 252 1205 255
rect 523 224 1205 252
rect 523 221 535 224
rect 477 215 535 221
rect 1193 221 1205 224
rect 1239 221 1251 255
rect 1193 215 1251 221
rect 1409 250 1467 256
rect 1409 216 1421 250
rect 1455 216 1467 250
rect 1409 197 1467 216
rect 1726 211 1744 263
rect 1796 211 1812 263
rect 1409 194 1531 197
rect 749 187 879 193
rect 749 153 761 187
rect 795 153 833 187
rect 867 184 879 187
rect 1409 184 1471 194
rect 867 156 1471 184
rect 867 153 879 156
rect 749 147 879 153
rect 1107 146 1471 156
rect 1107 48 1160 146
rect 1463 142 1471 146
rect 1523 142 1531 194
rect 1463 48 1531 142
rect 1726 142 1812 211
rect 2035 262 2221 268
rect 2035 210 2041 262
rect 2093 210 2221 262
rect 2035 204 2221 210
rect 2327 265 2548 271
rect 4674 270 4713 664
rect 2327 233 2486 265
rect 2327 142 2357 233
rect 2406 213 2486 233
rect 2538 213 2548 265
rect 4498 265 4713 270
rect 2576 255 2634 261
rect 2576 221 2588 255
rect 2622 252 2634 255
rect 2943 255 3001 261
rect 2943 252 2955 255
rect 2622 224 2955 252
rect 2622 221 2634 224
rect 2576 215 2634 221
rect 2943 221 2955 224
rect 2989 252 3001 255
rect 3659 255 3717 261
rect 3659 252 3671 255
rect 2989 224 3671 252
rect 2989 221 3001 224
rect 2943 215 3001 221
rect 3659 221 3671 224
rect 3705 221 3717 255
rect 3659 215 3717 221
rect 3875 250 3933 256
rect 3875 216 3887 250
rect 3921 216 3933 250
rect 2406 206 2548 213
rect 3875 196 3933 216
rect 4498 213 4510 265
rect 4562 213 4713 265
rect 4498 206 4713 213
rect 3215 187 3345 193
rect 3215 153 3227 187
rect 3261 153 3299 187
rect 3333 184 3345 187
rect 3875 192 4004 196
rect 3875 184 3940 192
rect 3333 156 3940 184
rect 3333 153 3345 156
rect 3215 147 3345 153
rect 1726 104 2357 142
rect 2136 100 2357 104
rect 3930 140 3940 156
rect 3992 140 4004 192
rect 2136 75 2172 100
rect 0 17 2116 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 -48 2116 -17
rect -1 -95 2116 -48
rect 1107 -580 1160 -95
rect 2144 -132 2172 75
rect 3930 87 4004 140
rect 3930 48 4929 87
rect 2466 31 4929 48
rect 2466 17 4582 31
rect 2466 -17 2495 17
rect 2529 -17 2587 17
rect 2621 -17 2679 17
rect 2713 -17 2771 17
rect 2805 -17 2863 17
rect 2897 -17 2955 17
rect 2989 -17 3047 17
rect 3081 -17 3139 17
rect 3173 -17 3231 17
rect 3265 -17 3323 17
rect 3357 -17 3415 17
rect 3449 -17 3507 17
rect 3541 -17 3599 17
rect 3633 -17 3691 17
rect 3725 -17 3783 17
rect 3817 -17 3875 17
rect 3909 -17 3967 17
rect 4001 -17 4059 17
rect 4093 -17 4151 17
rect 4185 -17 4243 17
rect 4277 -17 4335 17
rect 4369 -17 4427 17
rect 4461 -17 4519 17
rect 4553 -17 4582 17
rect 2466 -48 4582 -17
rect 2467 -87 4583 -48
rect 1108 -924 1160 -580
rect 1341 -161 2172 -132
rect 1341 -165 1390 -161
rect 1722 -165 2172 -161
rect 1341 -531 1369 -165
rect 2756 -180 4713 -151
rect 2756 -210 2827 -180
rect 1418 -241 1694 -210
rect 1418 -275 1447 -241
rect 1481 -275 1539 -241
rect 1573 -275 1631 -241
rect 1665 -275 1694 -241
rect 1418 -306 1694 -275
rect 2466 -241 4582 -210
rect 2466 -275 2495 -241
rect 2529 -275 2587 -241
rect 2621 -275 2679 -241
rect 2713 -275 2771 -241
rect 2805 -275 2863 -241
rect 2897 -275 2955 -241
rect 2989 -275 3047 -241
rect 3081 -275 3139 -241
rect 3173 -275 3231 -241
rect 3265 -275 3323 -241
rect 3357 -275 3415 -241
rect 3449 -275 3507 -241
rect 3541 -275 3599 -241
rect 3633 -275 3691 -241
rect 3725 -275 3783 -241
rect 3817 -275 3875 -241
rect 3909 -275 3967 -241
rect 4001 -275 4059 -241
rect 4093 -275 4151 -241
rect 4185 -275 4243 -241
rect 4277 -275 4335 -241
rect 4369 -275 4427 -241
rect 4461 -275 4519 -241
rect 4553 -275 4582 -241
rect 2466 -306 4582 -275
rect 2657 -411 2715 -405
rect 2657 -445 2669 -411
rect 2703 -414 2715 -411
rect 2756 -414 2827 -306
rect 3035 -411 3093 -405
rect 3035 -414 3047 -411
rect 2703 -442 3047 -414
rect 2703 -445 2715 -442
rect 2657 -451 2715 -445
rect 2756 -497 2827 -442
rect 3035 -445 3047 -442
rect 3081 -414 3093 -411
rect 3659 -411 3717 -405
rect 3659 -414 3671 -411
rect 3081 -442 3671 -414
rect 3081 -445 3093 -442
rect 3035 -451 3093 -445
rect 3659 -445 3671 -442
rect 3705 -445 3717 -411
rect 3659 -451 3717 -445
rect 2025 -500 2173 -499
rect 2025 -506 2545 -500
rect 1341 -547 1487 -531
rect 1341 -567 1447 -547
rect 1481 -567 1487 -547
rect 2025 -558 2487 -506
rect 2539 -558 2545 -506
rect 2025 -563 2545 -558
rect 1341 -619 1432 -567
rect 1484 -619 1487 -567
rect 1341 -631 1487 -619
rect 1524 -564 2545 -563
rect 2576 -547 2634 -541
rect 1524 -569 2077 -564
rect 1524 -621 1530 -569
rect 1582 -621 2077 -569
rect 2576 -581 2588 -547
rect 2622 -550 2634 -547
rect 2756 -549 2766 -497
rect 2818 -549 2827 -497
rect 2756 -550 2827 -549
rect 2943 -547 3001 -541
rect 2943 -550 2955 -547
rect 2622 -578 2955 -550
rect 2622 -581 2634 -578
rect 2576 -587 2634 -581
rect 2943 -581 2955 -578
rect 2989 -550 3001 -547
rect 3659 -547 3717 -541
rect 3659 -550 3671 -547
rect 2989 -578 3671 -550
rect 2989 -581 3001 -578
rect 2943 -587 3001 -581
rect 3659 -581 3671 -578
rect 3705 -581 3717 -547
rect 3659 -587 3717 -581
rect 3875 -552 3933 -546
rect 3875 -586 3887 -552
rect 3921 -586 3933 -552
rect 4668 -567 4713 -180
rect 3875 -604 3933 -586
rect 4502 -571 4713 -567
rect 3875 -609 4005 -604
rect 1524 -627 2077 -621
rect 3215 -615 3345 -609
rect 3215 -649 3227 -615
rect 3261 -649 3299 -615
rect 3333 -618 3345 -615
rect 3875 -618 3940 -609
rect 3333 -646 3940 -618
rect 3333 -649 3345 -646
rect 3215 -655 3345 -649
rect 3930 -661 3940 -646
rect 3992 -661 4005 -609
rect 4502 -623 4508 -571
rect 4560 -623 4713 -571
rect 4502 -627 4713 -623
rect 4668 -628 4713 -627
rect 3930 -754 4005 -661
rect 1418 -785 1694 -754
rect 1418 -819 1447 -785
rect 1481 -819 1539 -785
rect 1573 -819 1631 -785
rect 1665 -819 1694 -785
rect 1418 -876 1694 -819
rect 2466 -785 4582 -754
rect 2466 -819 2495 -785
rect 2529 -819 2587 -785
rect 2621 -819 2679 -785
rect 2713 -819 2771 -785
rect 2805 -819 2863 -785
rect 2897 -819 2955 -785
rect 2989 -819 3047 -785
rect 3081 -819 3139 -785
rect 3173 -819 3231 -785
rect 3265 -819 3323 -785
rect 3357 -819 3415 -785
rect 3449 -819 3507 -785
rect 3541 -819 3599 -785
rect 3633 -819 3691 -785
rect 3725 -819 3783 -785
rect 3817 -819 3875 -785
rect 3909 -819 3967 -785
rect 4001 -819 4059 -785
rect 4093 -819 4151 -785
rect 4185 -819 4243 -785
rect 4277 -819 4335 -785
rect 4369 -819 4427 -785
rect 4461 -819 4519 -785
rect 4553 -819 4582 -785
rect 2466 -868 4582 -819
rect 3930 -924 4005 -868
rect 4869 -924 4929 31
rect 1108 -961 4931 -924
rect 1108 -963 3943 -961
rect 4004 -962 4931 -961
<< via1 >>
rect 297 323 349 335
rect 297 289 305 323
rect 305 289 339 323
rect 339 289 349 323
rect 297 283 349 289
rect 2763 323 2815 336
rect 2763 289 2771 323
rect 2771 289 2805 323
rect 2805 289 2815 323
rect 2763 284 2815 289
rect 1744 253 1796 263
rect 1744 218 1754 253
rect 1754 218 1788 253
rect 1788 218 1796 253
rect 1744 211 1796 218
rect 1471 187 1523 194
rect 1471 153 1481 187
rect 1481 153 1515 187
rect 1515 153 1523 187
rect 1471 142 1523 153
rect 2041 254 2093 262
rect 2041 220 2049 254
rect 2049 220 2083 254
rect 2083 220 2093 254
rect 2041 210 2093 220
rect 2486 255 2538 265
rect 2486 221 2496 255
rect 2496 221 2530 255
rect 2530 221 2538 255
rect 2486 213 2538 221
rect 4510 255 4562 265
rect 4510 221 4517 255
rect 4517 221 4551 255
rect 4551 221 4562 255
rect 4510 213 4562 221
rect 3940 187 3992 192
rect 3940 153 3947 187
rect 3947 153 3981 187
rect 3981 153 3992 187
rect 3940 140 3992 153
rect 2487 -513 2539 -506
rect 2487 -547 2496 -513
rect 2496 -547 2531 -513
rect 2531 -547 2539 -513
rect 2487 -558 2539 -547
rect 1432 -581 1447 -567
rect 1447 -581 1481 -567
rect 1481 -581 1484 -567
rect 1432 -619 1484 -581
rect 1530 -577 1582 -569
rect 1530 -611 1539 -577
rect 1539 -611 1573 -577
rect 1573 -611 1582 -577
rect 1530 -621 1582 -611
rect 2766 -509 2818 -497
rect 2766 -543 2771 -509
rect 2771 -543 2805 -509
rect 2805 -543 2818 -509
rect 2766 -549 2818 -543
rect 3940 -615 3992 -609
rect 3940 -649 3947 -615
rect 3947 -649 3981 -615
rect 3981 -649 3992 -615
rect 3940 -661 3992 -649
rect 4508 -578 4560 -571
rect 4508 -612 4515 -578
rect 4515 -612 4549 -578
rect 4549 -612 4560 -578
rect 4508 -623 4560 -612
<< metal2 >>
rect 291 672 2223 715
rect 4674 714 4713 715
rect 291 660 2156 672
rect 291 335 355 660
rect 291 283 297 335
rect 349 283 355 335
rect 291 280 355 283
rect 1727 263 1812 285
rect 2185 268 2221 672
rect 2757 664 4713 714
rect 2757 336 2822 664
rect 2757 284 2763 336
rect 2815 284 2822 336
rect 2757 280 2822 284
rect 1727 211 1744 263
rect 1796 211 1812 263
rect 1463 194 1531 196
rect 1463 183 1471 194
rect 1107 146 1471 183
rect 1107 -580 1160 146
rect 1463 142 1471 146
rect 1523 142 1531 194
rect 1463 135 1531 142
rect 1727 142 1812 211
rect 2035 262 2221 268
rect 2035 210 2041 262
rect 2093 210 2221 262
rect 2035 204 2221 210
rect 2327 265 2548 271
rect 4674 270 4713 664
rect 2327 233 2486 265
rect 2327 142 2357 233
rect 2406 213 2486 233
rect 2538 213 2548 265
rect 2406 205 2548 213
rect 4498 265 4713 270
rect 4498 213 4510 265
rect 4562 213 4713 265
rect 4498 206 4713 213
rect 1727 104 2357 142
rect 2136 100 2357 104
rect 3930 192 4004 196
rect 3930 140 3940 192
rect 3992 140 4004 192
rect 2136 75 2172 100
rect 2144 -132 2172 75
rect 3930 87 4004 140
rect 3930 31 4929 87
rect 1108 -924 1160 -580
rect 1341 -161 2172 -132
rect 1341 -165 1390 -161
rect 1722 -165 2172 -161
rect 1341 -531 1369 -165
rect 2756 -180 4713 -151
rect 2756 -497 2827 -180
rect 2025 -500 2173 -499
rect 2025 -506 2545 -500
rect 1341 -567 1487 -531
rect 2025 -558 2487 -506
rect 2539 -558 2545 -506
rect 2756 -549 2766 -497
rect 2818 -549 2827 -497
rect 2756 -551 2827 -549
rect 2025 -563 2545 -558
rect 1341 -619 1432 -567
rect 1484 -619 1487 -567
rect 1341 -631 1487 -619
rect 1524 -564 2545 -563
rect 1524 -569 2077 -564
rect 4668 -567 4713 -180
rect 1524 -621 1530 -569
rect 1582 -621 2077 -569
rect 4502 -571 4713 -567
rect 1524 -627 2077 -621
rect 3930 -609 4005 -604
rect 3930 -661 3940 -609
rect 3992 -661 4005 -609
rect 4502 -623 4508 -571
rect 4560 -623 4713 -571
rect 4502 -627 4713 -623
rect 4668 -628 4713 -627
rect 3930 -924 4005 -661
rect 4869 -924 4929 31
rect 1108 -961 4931 -924
rect 1108 -963 3943 -961
rect 4004 -962 4931 -961
<< labels >>
flabel locali 1447 -581 1481 -547 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0/A
flabel locali 1539 -649 1573 -615 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0/Y
flabel locali 1539 -513 1573 -479 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0/Y
flabel locali 1539 -581 1573 -547 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0/Y
flabel nwell 1447 -275 1481 -241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0/VPB
flabel pwell 1447 -819 1481 -785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0/VNB
flabel metal1 1447 -275 1481 -241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0/VPWR
flabel metal1 1447 -819 1481 -785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0/VGND
rlabel comment 1418 -802 1418 -802 4 sky130_fd_sc_hd__inv_2_0/inv_2
flabel locali 4220 218 4249 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/Q
flabel locali 4522 221 4544 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/Q_N
flabel locali 3947 153 3981 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 2771 289 2805 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/D
flabel locali 2496 289 2530 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 2496 221 2530 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 3947 221 3981 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel metal1 2495 -17 2529 17 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VGND
flabel metal1 2495 527 2529 561 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VPWR
flabel nwell 2495 527 2529 561 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VPB
flabel pwell 2495 -17 2529 17 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_1/VNB
rlabel comment 2466 0 2466 0 4 sky130_fd_sc_hd__dfrbp_1_1/dfrbp_1
rlabel viali 3947 153 3981 187 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel viali 3887 216 3921 250 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 3947 127 3995 207 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 3887 207 3995 281 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3935 147 3993 156 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3875 193 3933 256 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3875 184 3993 193 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3215 184 3345 193 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3215 156 3993 184 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 3215 147 3345 156 1 sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 1754 218 1783 253 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q
flabel locali 2056 221 2078 254 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/Q_N
flabel locali 1481 153 1515 187 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 305 289 339 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/D
flabel locali 30 289 64 323 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 30 221 64 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 1481 221 1515 255 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 29 -17 63 17 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VGND
flabel metal1 29 527 63 561 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPWR
flabel nwell 29 527 63 561 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VPB
flabel pwell 29 -17 63 17 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_0/VNB
rlabel comment 0 0 0 0 4 sky130_fd_sc_hd__dfrbp_1_0/dfrbp_1
rlabel viali 1481 153 1515 187 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel viali 1421 216 1455 250 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1481 127 1529 207 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 1421 207 1529 281 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1469 147 1527 156 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1409 193 1467 256 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 1409 184 1527 193 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 749 184 879 193 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 749 156 1527 184 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 749 147 879 156 1 sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 4220 -584 4249 -549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/Q
flabel locali 4522 -581 4544 -548 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/Q_N
flabel locali 3947 -649 3981 -615 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
flabel locali 2771 -513 2805 -479 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/D
flabel locali 2496 -513 2530 -479 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/CLK
flabel locali 2496 -581 2530 -547 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/CLK
flabel locali 3947 -581 3981 -547 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
flabel metal1 2495 -819 2529 -785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/VGND
flabel metal1 2495 -275 2529 -241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/VPWR
flabel nwell 2495 -275 2529 -241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/VPB
flabel pwell 2495 -819 2529 -785 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfrbp_1_2/VNB
rlabel comment 2466 -802 2466 -802 4 sky130_fd_sc_hd__dfrbp_1_2/dfrbp_1
rlabel viali 3947 -649 3981 -615 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel viali 3887 -586 3921 -552 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel locali 3947 -675 3995 -595 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel locali 3887 -595 3995 -521 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3935 -655 3993 -646 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3875 -609 3933 -546 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3875 -618 3993 -609 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3215 -618 3345 -609 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3215 -646 3993 -618 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 3215 -655 3345 -646 1 sky130_fd_sc_hd__dfrbp_1_2/RESET_B
<< end >>
