* SPICE3 file created from extract1.ext - technology: sky130A

X0 out clkb_in net2 GND sky130_fd_pr__nfet_01v8 ad=3.012e+11p pd=2.62e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X1 net2 cl_in in GND sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=4.588e+11p ps=1.3325e+06u w=1e+06u l=150000u
X2 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X3 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X4 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X5 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X6 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X7 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X8 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X9 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X10 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X11 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X12 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X13 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X14 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X15 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X16 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X17 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X18 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X19 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X20 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X21 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X22 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X23 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X24 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X25 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X26 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X27 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X28 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X29 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X30 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X31 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X32 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X33 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X34 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X35 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X36 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X37 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X38 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X39 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X40 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X41 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X42 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X43 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X44 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X45 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X46 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X47 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X48 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X49 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X50 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X51 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X52 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X53 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X54 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X55 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X56 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X57 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X58 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X59 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X60 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X61 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X62 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X63 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X64 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X65 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X66 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X67 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X68 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X69 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X70 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X71 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X72 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X73 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X74 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X75 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X76 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X77 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X78 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X79 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X80 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X81 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X82 out clkb_in net1 VDD sky130_fd_pr__pfet_01v8 ad=6.6085e+11p pd=1.8025e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X83 net1 cl_in in VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=6.012e+11p ps=4.62e+06u w=2e+06u l=150000u
X84 out cl_in net2 VDD sky130_fd_pr__pfet_01v8 ad=6.6085e+11p pd=1.8025e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X85 net2 clkb_in in VDD sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=6.012e+11p ps=4.62e+06u w=2e+06u l=150000u
X86 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X87 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X88 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X89 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X90 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X91 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X92 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X93 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X94 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X95 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X96 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X97 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X98 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X99 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X100 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X101 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X102 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X103 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X104 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X105 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X106 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X107 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X108 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X109 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X110 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X111 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X112 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X113 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X114 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X115 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X116 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X117 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X118 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X119 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X120 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X121 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X122 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X123 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X124 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X125 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X126 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X127 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X128 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X129 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X130 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X131 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X132 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X133 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X134 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X135 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X136 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X137 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X138 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X139 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X140 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X141 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X142 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X143 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X144 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X145 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X146 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X147 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X148 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X149 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X150 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X151 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X152 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X153 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X154 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X155 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X156 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X157 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X158 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X159 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X160 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X161 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X162 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X163 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X164 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X165 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X166 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X167 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X168 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X169 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X170 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X171 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X172 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X173 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X174 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X175 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X176 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X177 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X178 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X179 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X180 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X181 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X182 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X183 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X184 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X185 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X186 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X187 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X188 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X189 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X190 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X191 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X192 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X193 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X194 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X195 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X196 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X197 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X198 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X199 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X200 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X201 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X202 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X203 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X204 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X205 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X206 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X207 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X208 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X209 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X210 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X211 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X212 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X213 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X214 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X215 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X216 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X217 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X218 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X219 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X220 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X221 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X222 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X223 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X224 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X225 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X226 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X227 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X228 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X229 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X230 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X231 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X232 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X233 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X234 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X235 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X236 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X237 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X238 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X239 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X240 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X241 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X242 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X243 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X244 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X245 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X246 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X247 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X248 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X249 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X250 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X251 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X252 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X253 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X254 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X255 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X256 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X257 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X258 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X259 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X260 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X261 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X262 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X263 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X264 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X265 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X266 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X267 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X268 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X269 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X270 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X271 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X272 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X273 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X274 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X275 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X276 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X277 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X278 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X279 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X280 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X281 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X282 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X283 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X284 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X285 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X286 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X287 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X288 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X289 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X290 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X291 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X292 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X293 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X294 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X295 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X296 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X297 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X298 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X299 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X300 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X301 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X302 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X303 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X304 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X305 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X306 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X307 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X308 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X309 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X310 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X311 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X312 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X313 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X314 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X315 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X316 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X317 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X318 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X319 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X320 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X321 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X322 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X323 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X324 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X325 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X326 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X327 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X328 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X329 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X330 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X331 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X332 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X333 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X334 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X335 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X336 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X337 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X338 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X339 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X340 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X341 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X342 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X343 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X344 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X345 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X346 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X347 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X348 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X349 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X350 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X351 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X352 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X353 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X354 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X355 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X356 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X357 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X358 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X359 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X360 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X361 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X362 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X363 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X364 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X365 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X366 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X367 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X368 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X369 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X370 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X371 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X372 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X373 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X374 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X375 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X376 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X377 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X378 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X379 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X380 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X381 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X382 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X383 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X384 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X385 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X386 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X387 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X388 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X389 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X390 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X391 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X392 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X393 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X394 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X395 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X396 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X397 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X398 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X399 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X400 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X401 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X402 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X403 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X404 VDD net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X405 VDD net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.04037e+12p pd=7.47225e+06u as=1.04037e+12p ps=7.47225e+06u w=7e+06u l=8e+06u
X406 out cl_in net1 GND sky130_fd_pr__nfet_01v8 ad=3.012e+11p pd=2.62e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X407 net1 clkb_in in GND sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=4.588e+11p ps=1.3325e+06u w=1e+06u l=150000u

