**.subckt 20bitCounter
x1 CLK net1 RESET GND VDD out0 net1 sky130_fd_sc_hd__dfrbp_1
x2 net1 net2 RESET GND VDD out1 net2 sky130_fd_sc_hd__dfrbp_1
x3 net2 net3 RESET GND VDD out2 net3 sky130_fd_sc_hd__dfrbp_1
x4 net3 net4 RESET GND VDD out3 net4 sky130_fd_sc_hd__dfrbp_1
x5 net4 net5 RESET GND VDD out4 net5 sky130_fd_sc_hd__dfrbp_1
x6 net5 net6 RESET GND VDD out5 net6 sky130_fd_sc_hd__dfrbp_1
x7 net6 net7 RESET GND VDD out6 net7 sky130_fd_sc_hd__dfrbp_1
x8 net7 net8 RESET GND VDD out7 net8 sky130_fd_sc_hd__dfrbp_1
x9 net8 net9 RESET GND VDD out8 net9 sky130_fd_sc_hd__dfrbp_1
x10 net9 net10 RESET GND VDD out9 net10 sky130_fd_sc_hd__dfrbp_1
x11 net10 net11 RESET GND VDD out10 net11 sky130_fd_sc_hd__dfrbp_1
x12 net11 net12 RESET GND VDD out11 net12 sky130_fd_sc_hd__dfrbp_1
x13 net12 net13 RESET GND VDD out12 net13 sky130_fd_sc_hd__dfrbp_1
x14 net13 net14 RESET GND VDD out13 net14 sky130_fd_sc_hd__dfrbp_1
x15 net14 net15 RESET GND VDD out14 net15 sky130_fd_sc_hd__dfrbp_1
x16 net15 net16 RESET GND VDD out15 net16 sky130_fd_sc_hd__dfrbp_1
x17 net16 net17 RESET GND VDD out16 net17 sky130_fd_sc_hd__dfrbp_1
x18 net17 net18 RESET GND VDD out17 net18 sky130_fd_sc_hd__dfrbp_1
x19 net18 net19 RESET GND VDD out18 net19 sky130_fd_sc_hd__dfrbp_1
x20 net19 net20 RESET GND VDD out19 net20 sky130_fd_sc_hd__dfrbp_1
**** begin user architecture code
.lib ~/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ~/Documents/counter/layout/lvs_check/tempFix/poseEdge_Dff.spice
**** end user architecture code
**.ends
** flattened .save nodes
.end
