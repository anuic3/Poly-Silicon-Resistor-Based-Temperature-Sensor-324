magic
tech sky130A
magscale 1 2
timestamp 1634913479
<< nwell >>
rect -96394 4314 -26088 22510
rect 844 4522 18876 6254
rect 844 4518 9820 4522
rect 10122 4518 18876 4522
rect 13112 4412 16262 4518
rect 16924 4346 18024 4518
rect -96512 4182 -26088 4314
rect -96532 3980 -26088 4182
rect -96532 2872 -62316 3980
rect -62056 3950 -26096 3980
rect -62056 3916 -61162 3950
rect -61934 3758 -61162 3916
rect -61848 3380 -61162 3758
rect -61356 3378 -61162 3380
rect -60826 3184 -26096 3950
rect 25958 3872 28060 3874
rect -60826 2876 -26074 3184
rect -96396 2870 -62316 2872
rect 25958 2494 32912 3872
rect 26634 2450 32912 2494
rect 26634 2380 31924 2450
rect 32702 2448 32912 2450
rect 26634 2370 26856 2380
rect 27146 2378 31924 2380
rect 27156 2376 30882 2378
rect 31538 2376 31924 2378
rect 27156 2372 28128 2376
rect 28776 2374 30216 2376
rect 27156 2370 27824 2372
rect 29752 2370 30216 2374
rect 27694 1202 28914 1242
rect 27692 696 28914 1202
rect 27694 694 28914 696
rect 27694 692 28882 694
rect 27694 334 28852 692
rect 27694 -660 28850 334
rect 13186 -862 13355 -769
rect 8696 -1258 10888 -863
rect 11162 -937 13355 -862
rect 11162 -1258 13354 -937
rect 27694 -1020 28846 -660
rect 10116 -1705 10464 -1700
rect 10114 -2060 10466 -1705
rect 11162 -2060 13354 -1693
rect -9196 -4528 33200 -4168
rect 8858 -7215 16374 -7213
rect 8858 -7862 16786 -7215
rect 8858 -7885 16808 -7862
rect 8871 -9268 16808 -7885
rect 8872 -9331 16808 -9268
rect 16062 -9333 16808 -9331
rect 8844 -14941 16816 -13689
rect 16458 -19387 16920 -19385
rect 8619 -19416 9081 -19403
rect 16458 -19416 17340 -19387
rect 8619 -20181 17340 -19416
rect 8619 -20829 16490 -20181
rect 8866 -20832 16490 -20829
<< pwell >>
rect 9637 -1362 9823 -1318
rect 10367 -1362 10838 -1316
rect 12103 -1362 12289 -1318
rect 12833 -1362 13304 -1316
rect 8735 -1498 10838 -1362
rect 11201 -1498 13304 -1362
rect 8763 -1536 8797 -1498
rect 11229 -1536 11263 -1498
rect 10155 -2300 10425 -2118
rect 12103 -2164 12289 -2120
rect 12833 -2164 13304 -2118
rect 11201 -2300 13304 -2164
rect 10181 -2338 10215 -2300
rect 11229 -2338 11263 -2300
rect -8255 -4632 -8069 -4588
rect -7525 -4632 -7054 -4586
rect -6139 -4632 -5953 -4588
rect -5409 -4632 -4938 -4586
rect -4023 -4632 -3837 -4588
rect -3293 -4632 -2822 -4586
rect -1907 -4632 -1721 -4588
rect -1177 -4632 -706 -4586
rect 209 -4632 395 -4588
rect 939 -4632 1410 -4586
rect 2325 -4632 2511 -4588
rect 3055 -4632 3526 -4586
rect 4441 -4632 4627 -4588
rect 5171 -4632 5642 -4586
rect 6557 -4632 6743 -4588
rect 7287 -4632 7758 -4586
rect 8673 -4632 8859 -4588
rect 9403 -4632 9874 -4586
rect 10789 -4632 10975 -4588
rect 11519 -4632 11990 -4586
rect 12905 -4632 13091 -4588
rect 13635 -4632 14106 -4586
rect 15021 -4632 15207 -4588
rect 15751 -4632 16222 -4586
rect 17137 -4632 17323 -4588
rect 17867 -4632 18338 -4586
rect 19253 -4632 19439 -4588
rect 19983 -4632 20454 -4586
rect 21369 -4632 21555 -4588
rect 22099 -4632 22570 -4586
rect 23485 -4632 23671 -4588
rect 24215 -4632 24686 -4586
rect 25601 -4632 25787 -4588
rect 26331 -4632 26802 -4586
rect 27717 -4632 27903 -4588
rect 28447 -4632 28918 -4586
rect 29833 -4632 30019 -4588
rect 30563 -4632 31034 -4586
rect 31949 -4632 32135 -4588
rect 32679 -4632 33150 -4586
rect -9157 -4741 -7054 -4632
rect -7041 -4741 -4938 -4632
rect -4925 -4741 -2822 -4632
rect -2809 -4741 -706 -4632
rect -693 -4741 1410 -4632
rect 1423 -4741 3526 -4632
rect 3539 -4741 5642 -4632
rect 5655 -4741 7758 -4632
rect 7771 -4741 9874 -4632
rect 9887 -4741 11990 -4632
rect 12003 -4741 14106 -4632
rect 14119 -4741 16222 -4632
rect 16235 -4741 18338 -4632
rect 18351 -4741 20454 -4632
rect 20467 -4741 22570 -4632
rect 22583 -4741 24686 -4632
rect 24699 -4741 26802 -4632
rect 26815 -4741 28918 -4632
rect 28931 -4741 31034 -4632
rect 31047 -4741 33150 -4632
rect -9158 -4866 33162 -4741
rect 4219 -7520 4231 -7514
rect 4219 -25843 7869 -7520
rect 17840 -7519 17852 -7513
rect 16836 -20199 16922 -20181
rect 16508 -20677 17312 -20199
rect 16508 -20699 16922 -20677
rect 16508 -20703 17352 -20699
rect 17840 -25842 21490 -7519
<< nmos >>
rect 1144 4200 1174 4400
rect 1360 4202 1390 4402
rect 1578 4202 1608 4402
rect 1800 4200 1830 4400
rect 6330 4218 6360 4418
rect 6546 4220 6576 4420
rect 6764 4220 6794 4420
rect 6986 4218 7016 4418
rect 11506 4230 11536 4430
rect 11722 4232 11752 4432
rect 11940 4232 11970 4432
rect 12162 4230 12192 4430
rect 17162 4022 17192 4222
rect 17378 4024 17408 4224
rect 17596 4024 17626 4224
rect 17818 4022 17848 4222
rect -61768 3046 -61738 3246
rect -61672 3046 -61642 3246
rect -61576 3046 -61546 3246
rect -61480 3046 -61450 3246
rect 26936 2060 26966 2208
rect 27032 2060 27062 2208
rect 27548 2068 27578 2216
rect 27644 2068 27674 2216
rect 28126 2064 28156 2212
rect 28222 2064 28252 2212
rect 28700 2072 28730 2220
rect 28796 2072 28826 2220
rect 29278 2072 29308 2220
rect 29374 2072 29404 2220
rect 29856 2072 29886 2220
rect 29952 2072 29982 2220
rect 30438 2076 30468 2224
rect 30534 2076 30564 2224
rect 31014 2072 31044 2220
rect 31110 2072 31140 2220
rect 31584 2068 31614 2216
rect 31680 2068 31710 2216
rect 28994 -278 29024 370
rect 29090 -278 29120 370
rect 29186 -278 29216 370
rect 29282 -278 29312 370
rect 29378 -278 29408 370
rect 29474 -278 29504 370
rect 29570 -278 29600 370
rect 29666 -278 29696 370
rect 29762 -278 29792 370
rect 4415 -9023 6015 -7623
rect 6073 -9023 7673 -7623
rect 4415 -10533 6015 -9133
rect 6073 -10533 7673 -9133
rect 4415 -12043 6015 -10643
rect 6073 -12043 7673 -10643
rect 4415 -13553 6015 -12153
rect 6073 -13553 7673 -12153
rect 4415 -15063 6015 -13663
rect 6073 -15063 7673 -13663
rect 4415 -16573 6015 -15173
rect 6073 -16573 7673 -15173
rect 4415 -18083 6015 -16683
rect 6073 -18083 7673 -16683
rect 4415 -19593 6015 -18193
rect 6073 -19593 7673 -18193
rect 4415 -21103 6015 -19703
rect 6073 -21103 7673 -19703
rect 4415 -22613 6015 -21213
rect 6073 -22613 7673 -21213
rect 4415 -24123 6015 -22723
rect 6073 -24123 7673 -22723
rect 4415 -25633 6015 -24233
rect 6073 -25633 7673 -24233
rect 16704 -20493 16734 -20409
rect 17094 -20493 17124 -20409
rect 18036 -9022 19636 -7622
rect 19694 -9022 21294 -7622
rect 18036 -10532 19636 -9132
rect 19694 -10532 21294 -9132
rect 18036 -12042 19636 -10642
rect 19694 -12042 21294 -10642
rect 18036 -13552 19636 -12152
rect 19694 -13552 21294 -12152
rect 18036 -15062 19636 -13662
rect 19694 -15062 21294 -13662
rect 18036 -16572 19636 -15172
rect 19694 -16572 21294 -15172
rect 18036 -18082 19636 -16682
rect 19694 -18082 21294 -16682
rect 18036 -19592 19636 -18192
rect 19694 -19592 21294 -18192
rect 18036 -21102 19636 -19702
rect 19694 -21102 21294 -19702
rect 18036 -22612 19636 -21212
rect 19694 -22612 21294 -21212
rect 18036 -24122 19636 -22722
rect 19694 -24122 21294 -22722
rect 18036 -25632 19636 -24232
rect 19694 -25632 21294 -24232
<< scnmos >>
rect 8813 -1472 8843 -1388
rect 8897 -1472 8927 -1388
rect 9152 -1472 9182 -1388
rect 9247 -1472 9277 -1400
rect 9343 -1472 9373 -1400
rect 9509 -1472 9539 -1388
rect 9581 -1472 9611 -1388
rect 9713 -1472 9743 -1344
rect 9812 -1472 9842 -1400
rect 9921 -1472 9951 -1400
rect 10017 -1472 10047 -1388
rect 10166 -1472 10196 -1388
rect 10257 -1472 10287 -1388
rect 10445 -1472 10475 -1342
rect 10633 -1472 10663 -1388
rect 10730 -1472 10760 -1342
rect 11279 -1472 11309 -1388
rect 11363 -1472 11393 -1388
rect 11618 -1472 11648 -1388
rect 11713 -1472 11743 -1400
rect 11809 -1472 11839 -1400
rect 11975 -1472 12005 -1388
rect 12047 -1472 12077 -1388
rect 12179 -1472 12209 -1344
rect 12278 -1472 12308 -1400
rect 12387 -1472 12417 -1400
rect 12483 -1472 12513 -1388
rect 12632 -1472 12662 -1388
rect 12723 -1472 12753 -1388
rect 12911 -1472 12941 -1342
rect 13099 -1472 13129 -1388
rect 13196 -1472 13226 -1342
rect 10233 -2274 10263 -2144
rect 10317 -2274 10347 -2144
rect 11279 -2274 11309 -2190
rect 11363 -2274 11393 -2190
rect 11618 -2274 11648 -2190
rect 11713 -2274 11743 -2202
rect 11809 -2274 11839 -2202
rect 11975 -2274 12005 -2190
rect 12047 -2274 12077 -2190
rect 12179 -2274 12209 -2146
rect 12278 -2274 12308 -2202
rect 12387 -2274 12417 -2202
rect 12483 -2274 12513 -2190
rect 12632 -2274 12662 -2190
rect 12723 -2274 12753 -2190
rect 12911 -2274 12941 -2144
rect 13099 -2274 13129 -2190
rect 13196 -2274 13226 -2144
rect -9079 -4742 -9049 -4658
rect -8995 -4742 -8965 -4658
rect -8740 -4742 -8710 -4658
rect -8645 -4742 -8615 -4670
rect -8549 -4742 -8519 -4670
rect -8383 -4742 -8353 -4658
rect -8311 -4742 -8281 -4658
rect -8179 -4742 -8149 -4614
rect -8080 -4742 -8050 -4670
rect -7971 -4742 -7941 -4670
rect -7875 -4742 -7845 -4658
rect -7726 -4742 -7696 -4658
rect -7635 -4742 -7605 -4658
rect -7447 -4742 -7417 -4612
rect -7259 -4742 -7229 -4658
rect -7162 -4742 -7132 -4612
rect -6963 -4742 -6933 -4658
rect -6879 -4742 -6849 -4658
rect -6624 -4742 -6594 -4658
rect -6529 -4742 -6499 -4670
rect -6433 -4742 -6403 -4670
rect -6267 -4742 -6237 -4658
rect -6195 -4742 -6165 -4658
rect -6063 -4742 -6033 -4614
rect -5964 -4742 -5934 -4670
rect -5855 -4742 -5825 -4670
rect -5759 -4742 -5729 -4658
rect -5610 -4742 -5580 -4658
rect -5519 -4742 -5489 -4658
rect -5331 -4742 -5301 -4612
rect -5143 -4742 -5113 -4658
rect -5046 -4742 -5016 -4612
rect -4847 -4742 -4817 -4658
rect -4763 -4742 -4733 -4658
rect -4508 -4742 -4478 -4658
rect -4413 -4742 -4383 -4670
rect -4317 -4742 -4287 -4670
rect -4151 -4742 -4121 -4658
rect -4079 -4742 -4049 -4658
rect -3947 -4742 -3917 -4614
rect -3848 -4742 -3818 -4670
rect -3739 -4742 -3709 -4670
rect -3643 -4742 -3613 -4658
rect -3494 -4742 -3464 -4658
rect -3403 -4742 -3373 -4658
rect -3215 -4742 -3185 -4612
rect -3027 -4742 -2997 -4658
rect -2930 -4742 -2900 -4612
rect -2731 -4742 -2701 -4658
rect -2647 -4742 -2617 -4658
rect -2392 -4742 -2362 -4658
rect -2297 -4742 -2267 -4670
rect -2201 -4742 -2171 -4670
rect -2035 -4742 -2005 -4658
rect -1963 -4742 -1933 -4658
rect -1831 -4742 -1801 -4614
rect -1732 -4742 -1702 -4670
rect -1623 -4742 -1593 -4670
rect -1527 -4742 -1497 -4658
rect -1378 -4742 -1348 -4658
rect -1287 -4742 -1257 -4658
rect -1099 -4742 -1069 -4612
rect -911 -4742 -881 -4658
rect -814 -4742 -784 -4612
rect -615 -4742 -585 -4658
rect -531 -4742 -501 -4658
rect -276 -4742 -246 -4658
rect -181 -4742 -151 -4670
rect -85 -4742 -55 -4670
rect 81 -4742 111 -4658
rect 153 -4742 183 -4658
rect 285 -4742 315 -4614
rect 384 -4742 414 -4670
rect 493 -4742 523 -4670
rect 589 -4742 619 -4658
rect 738 -4742 768 -4658
rect 829 -4742 859 -4658
rect 1017 -4742 1047 -4612
rect 1205 -4742 1235 -4658
rect 1302 -4742 1332 -4612
rect 1501 -4742 1531 -4658
rect 1585 -4742 1615 -4658
rect 1840 -4742 1870 -4658
rect 1935 -4742 1965 -4670
rect 2031 -4742 2061 -4670
rect 2197 -4742 2227 -4658
rect 2269 -4742 2299 -4658
rect 2401 -4742 2431 -4614
rect 2500 -4742 2530 -4670
rect 2609 -4742 2639 -4670
rect 2705 -4742 2735 -4658
rect 2854 -4742 2884 -4658
rect 2945 -4742 2975 -4658
rect 3133 -4742 3163 -4612
rect 3321 -4742 3351 -4658
rect 3418 -4742 3448 -4612
rect 3617 -4742 3647 -4658
rect 3701 -4742 3731 -4658
rect 3956 -4742 3986 -4658
rect 4051 -4742 4081 -4670
rect 4147 -4742 4177 -4670
rect 4313 -4742 4343 -4658
rect 4385 -4742 4415 -4658
rect 4517 -4742 4547 -4614
rect 4616 -4742 4646 -4670
rect 4725 -4742 4755 -4670
rect 4821 -4742 4851 -4658
rect 4970 -4742 5000 -4658
rect 5061 -4742 5091 -4658
rect 5249 -4742 5279 -4612
rect 5437 -4742 5467 -4658
rect 5534 -4742 5564 -4612
rect 5733 -4742 5763 -4658
rect 5817 -4742 5847 -4658
rect 6072 -4742 6102 -4658
rect 6167 -4742 6197 -4670
rect 6263 -4742 6293 -4670
rect 6429 -4742 6459 -4658
rect 6501 -4742 6531 -4658
rect 6633 -4742 6663 -4614
rect 6732 -4742 6762 -4670
rect 6841 -4742 6871 -4670
rect 6937 -4742 6967 -4658
rect 7086 -4742 7116 -4658
rect 7177 -4742 7207 -4658
rect 7365 -4742 7395 -4612
rect 7553 -4742 7583 -4658
rect 7650 -4742 7680 -4612
rect 7849 -4742 7879 -4658
rect 7933 -4742 7963 -4658
rect 8188 -4742 8218 -4658
rect 8283 -4742 8313 -4670
rect 8379 -4742 8409 -4670
rect 8545 -4742 8575 -4658
rect 8617 -4742 8647 -4658
rect 8749 -4742 8779 -4614
rect 8848 -4742 8878 -4670
rect 8957 -4742 8987 -4670
rect 9053 -4742 9083 -4658
rect 9202 -4742 9232 -4658
rect 9293 -4742 9323 -4658
rect 9481 -4742 9511 -4612
rect 9669 -4742 9699 -4658
rect 9766 -4742 9796 -4612
rect 9965 -4742 9995 -4658
rect 10049 -4742 10079 -4658
rect 10304 -4742 10334 -4658
rect 10399 -4742 10429 -4670
rect 10495 -4742 10525 -4670
rect 10661 -4742 10691 -4658
rect 10733 -4742 10763 -4658
rect 10865 -4742 10895 -4614
rect 10964 -4742 10994 -4670
rect 11073 -4742 11103 -4670
rect 11169 -4742 11199 -4658
rect 11318 -4742 11348 -4658
rect 11409 -4742 11439 -4658
rect 11597 -4742 11627 -4612
rect 11785 -4742 11815 -4658
rect 11882 -4742 11912 -4612
rect 12081 -4742 12111 -4658
rect 12165 -4742 12195 -4658
rect 12420 -4742 12450 -4658
rect 12515 -4742 12545 -4670
rect 12611 -4742 12641 -4670
rect 12777 -4742 12807 -4658
rect 12849 -4742 12879 -4658
rect 12981 -4742 13011 -4614
rect 13080 -4742 13110 -4670
rect 13189 -4742 13219 -4670
rect 13285 -4742 13315 -4658
rect 13434 -4742 13464 -4658
rect 13525 -4742 13555 -4658
rect 13713 -4742 13743 -4612
rect 13901 -4742 13931 -4658
rect 13998 -4742 14028 -4612
rect 14197 -4742 14227 -4658
rect 14281 -4742 14311 -4658
rect 14536 -4742 14566 -4658
rect 14631 -4742 14661 -4670
rect 14727 -4742 14757 -4670
rect 14893 -4742 14923 -4658
rect 14965 -4742 14995 -4658
rect 15097 -4742 15127 -4614
rect 15196 -4742 15226 -4670
rect 15305 -4742 15335 -4670
rect 15401 -4742 15431 -4658
rect 15550 -4742 15580 -4658
rect 15641 -4742 15671 -4658
rect 15829 -4742 15859 -4612
rect 16017 -4742 16047 -4658
rect 16114 -4742 16144 -4612
rect 16313 -4742 16343 -4658
rect 16397 -4742 16427 -4658
rect 16652 -4742 16682 -4658
rect 16747 -4742 16777 -4670
rect 16843 -4742 16873 -4670
rect 17009 -4742 17039 -4658
rect 17081 -4742 17111 -4658
rect 17213 -4742 17243 -4614
rect 17312 -4742 17342 -4670
rect 17421 -4742 17451 -4670
rect 17517 -4742 17547 -4658
rect 17666 -4742 17696 -4658
rect 17757 -4742 17787 -4658
rect 17945 -4742 17975 -4612
rect 18133 -4742 18163 -4658
rect 18230 -4742 18260 -4612
rect 18429 -4742 18459 -4658
rect 18513 -4742 18543 -4658
rect 18768 -4742 18798 -4658
rect 18863 -4742 18893 -4670
rect 18959 -4742 18989 -4670
rect 19125 -4742 19155 -4658
rect 19197 -4742 19227 -4658
rect 19329 -4742 19359 -4614
rect 19428 -4742 19458 -4670
rect 19537 -4742 19567 -4670
rect 19633 -4742 19663 -4658
rect 19782 -4742 19812 -4658
rect 19873 -4742 19903 -4658
rect 20061 -4742 20091 -4612
rect 20249 -4742 20279 -4658
rect 20346 -4742 20376 -4612
rect 20545 -4742 20575 -4658
rect 20629 -4742 20659 -4658
rect 20884 -4742 20914 -4658
rect 20979 -4742 21009 -4670
rect 21075 -4742 21105 -4670
rect 21241 -4742 21271 -4658
rect 21313 -4742 21343 -4658
rect 21445 -4742 21475 -4614
rect 21544 -4742 21574 -4670
rect 21653 -4742 21683 -4670
rect 21749 -4742 21779 -4658
rect 21898 -4742 21928 -4658
rect 21989 -4742 22019 -4658
rect 22177 -4742 22207 -4612
rect 22365 -4742 22395 -4658
rect 22462 -4742 22492 -4612
rect 22661 -4742 22691 -4658
rect 22745 -4742 22775 -4658
rect 23000 -4742 23030 -4658
rect 23095 -4742 23125 -4670
rect 23191 -4742 23221 -4670
rect 23357 -4742 23387 -4658
rect 23429 -4742 23459 -4658
rect 23561 -4742 23591 -4614
rect 23660 -4742 23690 -4670
rect 23769 -4742 23799 -4670
rect 23865 -4742 23895 -4658
rect 24014 -4742 24044 -4658
rect 24105 -4742 24135 -4658
rect 24293 -4742 24323 -4612
rect 24481 -4742 24511 -4658
rect 24578 -4742 24608 -4612
rect 24777 -4742 24807 -4658
rect 24861 -4742 24891 -4658
rect 25116 -4742 25146 -4658
rect 25211 -4742 25241 -4670
rect 25307 -4742 25337 -4670
rect 25473 -4742 25503 -4658
rect 25545 -4742 25575 -4658
rect 25677 -4742 25707 -4614
rect 25776 -4742 25806 -4670
rect 25885 -4742 25915 -4670
rect 25981 -4742 26011 -4658
rect 26130 -4742 26160 -4658
rect 26221 -4742 26251 -4658
rect 26409 -4742 26439 -4612
rect 26597 -4742 26627 -4658
rect 26694 -4742 26724 -4612
rect 26893 -4742 26923 -4658
rect 26977 -4742 27007 -4658
rect 27232 -4742 27262 -4658
rect 27327 -4742 27357 -4670
rect 27423 -4742 27453 -4670
rect 27589 -4742 27619 -4658
rect 27661 -4742 27691 -4658
rect 27793 -4742 27823 -4614
rect 27892 -4742 27922 -4670
rect 28001 -4742 28031 -4670
rect 28097 -4742 28127 -4658
rect 28246 -4742 28276 -4658
rect 28337 -4742 28367 -4658
rect 28525 -4742 28555 -4612
rect 28713 -4742 28743 -4658
rect 28810 -4742 28840 -4612
rect 29009 -4742 29039 -4658
rect 29093 -4742 29123 -4658
rect 29348 -4742 29378 -4658
rect 29443 -4742 29473 -4670
rect 29539 -4742 29569 -4670
rect 29705 -4742 29735 -4658
rect 29777 -4742 29807 -4658
rect 29909 -4742 29939 -4614
rect 30008 -4742 30038 -4670
rect 30117 -4742 30147 -4670
rect 30213 -4742 30243 -4658
rect 30362 -4742 30392 -4658
rect 30453 -4742 30483 -4658
rect 30641 -4742 30671 -4612
rect 30829 -4742 30859 -4658
rect 30926 -4742 30956 -4612
rect 31125 -4742 31155 -4658
rect 31209 -4742 31239 -4658
rect 31464 -4742 31494 -4658
rect 31559 -4742 31589 -4670
rect 31655 -4742 31685 -4670
rect 31821 -4742 31851 -4658
rect 31893 -4742 31923 -4658
rect 32025 -4742 32055 -4614
rect 32124 -4742 32154 -4670
rect 32233 -4742 32263 -4670
rect 32329 -4742 32359 -4658
rect 32478 -4742 32508 -4658
rect 32569 -4742 32599 -4658
rect 32757 -4742 32787 -4612
rect 32945 -4742 32975 -4658
rect 33042 -4742 33072 -4612
<< pmos >>
rect -61720 3490 -61690 3890
rect -61624 3490 -61594 3890
rect -61528 3490 -61498 3890
rect -61432 3490 -61402 3890
rect 1120 4638 1150 5038
rect 1352 4636 1382 5036
rect 1580 4634 1610 5034
rect 1798 4636 1828 5036
rect 6306 4656 6336 5056
rect 6538 4654 6568 5054
rect 6766 4652 6796 5052
rect 6984 4654 7014 5054
rect 11482 4668 11512 5068
rect 11714 4666 11744 5066
rect 11942 4664 11972 5064
rect 12160 4666 12190 5066
rect 17138 4460 17168 4860
rect 17370 4458 17400 4858
rect 17598 4456 17628 4856
rect 17816 4458 17846 4858
rect 26932 2470 26962 2806
rect 27136 2508 27166 2844
rect 27544 2478 27574 2814
rect 27748 2516 27778 2852
rect 28122 2474 28152 2810
rect 28326 2512 28356 2848
rect 28696 2482 28726 2818
rect 28900 2520 28930 2856
rect 29274 2482 29304 2818
rect 29478 2520 29508 2856
rect 29852 2482 29882 2818
rect 30056 2520 30086 2856
rect 30434 2486 30464 2822
rect 30638 2524 30668 2860
rect 31010 2482 31040 2818
rect 31214 2520 31244 2856
rect 31580 2478 31610 2814
rect 31784 2516 31814 2852
rect 28326 416 28356 752
rect 28526 454 28556 790
rect 28728 414 28758 750
rect 28326 -90 28356 246
rect 28526 -52 28556 284
rect 28726 -90 28756 246
rect 28326 -598 28356 -262
rect 28526 -560 28556 -224
rect 28726 -598 28756 -262
rect 9384 -8759 9500 -8649
rect 10770 -8759 10886 -8649
rect 11140 -8759 11256 -8649
rect 11562 -8759 11678 -8649
rect 11984 -8759 12100 -8649
rect 13484 -8759 13600 -8649
rect 13854 -8759 13970 -8649
rect 14276 -8759 14392 -8649
rect 14698 -8759 14814 -8649
rect 16138 -8759 16254 -8649
rect 9384 -14441 9500 -14331
rect 10770 -14442 10886 -14332
rect 11140 -14442 11256 -14332
rect 11562 -14442 11678 -14332
rect 11984 -14442 12100 -14332
rect 13484 -14438 13600 -14328
rect 13854 -14438 13970 -14328
rect 14276 -14438 14392 -14328
rect 14698 -14438 14814 -14328
rect 16082 -14441 16198 -14331
rect 9429 -20365 9545 -20255
rect 10770 -20367 10886 -20257
rect 11140 -20367 11256 -20257
rect 11562 -20367 11678 -20257
rect 11984 -20367 12100 -20257
rect 13471 -20367 13587 -20257
rect 13841 -20367 13957 -20257
rect 14263 -20367 14379 -20257
rect 14685 -20367 14801 -20257
rect 16700 -19958 16730 -19622
rect 17090 -19960 17120 -19624
<< scpmoshvt >>
rect 8813 -1156 8843 -1028
rect 8897 -1156 8927 -1028
rect 9164 -1106 9194 -1022
rect 9256 -1106 9286 -1022
rect 9355 -1106 9385 -1022
rect 9495 -1106 9525 -1022
rect 9592 -1106 9622 -1022
rect 9789 -1190 9819 -1022
rect 9888 -1106 9918 -1022
rect 9974 -1106 10004 -1022
rect 10058 -1106 10088 -1022
rect 10166 -1106 10196 -1022
rect 10250 -1106 10280 -1022
rect 10414 -1222 10444 -1022
rect 10633 -1150 10663 -1022
rect 10730 -1222 10760 -1022
rect 11279 -1156 11309 -1028
rect 11363 -1156 11393 -1028
rect 11630 -1106 11660 -1022
rect 11722 -1106 11752 -1022
rect 11821 -1106 11851 -1022
rect 11961 -1106 11991 -1022
rect 12058 -1106 12088 -1022
rect 12255 -1190 12285 -1022
rect 12354 -1106 12384 -1022
rect 12440 -1106 12470 -1022
rect 12524 -1106 12554 -1022
rect 12632 -1106 12662 -1022
rect 12716 -1106 12746 -1022
rect 12880 -1222 12910 -1022
rect 13099 -1150 13129 -1022
rect 13196 -1222 13226 -1022
rect 10233 -2024 10263 -1824
rect 10317 -2024 10347 -1824
rect 11279 -1958 11309 -1830
rect 11363 -1958 11393 -1830
rect 11630 -1908 11660 -1824
rect 11722 -1908 11752 -1824
rect 11821 -1908 11851 -1824
rect 11961 -1908 11991 -1824
rect 12058 -1908 12088 -1824
rect 12255 -1992 12285 -1824
rect 12354 -1908 12384 -1824
rect 12440 -1908 12470 -1824
rect 12524 -1908 12554 -1824
rect 12632 -1908 12662 -1824
rect 12716 -1908 12746 -1824
rect 12880 -2024 12910 -1824
rect 13099 -1952 13129 -1824
rect 13196 -2024 13226 -1824
rect -9079 -4426 -9049 -4298
rect -8995 -4426 -8965 -4298
rect -8728 -4376 -8698 -4292
rect -8636 -4376 -8606 -4292
rect -8537 -4376 -8507 -4292
rect -8397 -4376 -8367 -4292
rect -8300 -4376 -8270 -4292
rect -8103 -4460 -8073 -4292
rect -8004 -4376 -7974 -4292
rect -7918 -4376 -7888 -4292
rect -7834 -4376 -7804 -4292
rect -7726 -4376 -7696 -4292
rect -7642 -4376 -7612 -4292
rect -7478 -4492 -7448 -4292
rect -7259 -4420 -7229 -4292
rect -7162 -4492 -7132 -4292
rect -6963 -4426 -6933 -4298
rect -6879 -4426 -6849 -4298
rect -6612 -4376 -6582 -4292
rect -6520 -4376 -6490 -4292
rect -6421 -4376 -6391 -4292
rect -6281 -4376 -6251 -4292
rect -6184 -4376 -6154 -4292
rect -5987 -4460 -5957 -4292
rect -5888 -4376 -5858 -4292
rect -5802 -4376 -5772 -4292
rect -5718 -4376 -5688 -4292
rect -5610 -4376 -5580 -4292
rect -5526 -4376 -5496 -4292
rect -5362 -4492 -5332 -4292
rect -5143 -4420 -5113 -4292
rect -5046 -4492 -5016 -4292
rect -4847 -4426 -4817 -4298
rect -4763 -4426 -4733 -4298
rect -4496 -4376 -4466 -4292
rect -4404 -4376 -4374 -4292
rect -4305 -4376 -4275 -4292
rect -4165 -4376 -4135 -4292
rect -4068 -4376 -4038 -4292
rect -3871 -4460 -3841 -4292
rect -3772 -4376 -3742 -4292
rect -3686 -4376 -3656 -4292
rect -3602 -4376 -3572 -4292
rect -3494 -4376 -3464 -4292
rect -3410 -4376 -3380 -4292
rect -3246 -4492 -3216 -4292
rect -3027 -4420 -2997 -4292
rect -2930 -4492 -2900 -4292
rect -2731 -4426 -2701 -4298
rect -2647 -4426 -2617 -4298
rect -2380 -4376 -2350 -4292
rect -2288 -4376 -2258 -4292
rect -2189 -4376 -2159 -4292
rect -2049 -4376 -2019 -4292
rect -1952 -4376 -1922 -4292
rect -1755 -4460 -1725 -4292
rect -1656 -4376 -1626 -4292
rect -1570 -4376 -1540 -4292
rect -1486 -4376 -1456 -4292
rect -1378 -4376 -1348 -4292
rect -1294 -4376 -1264 -4292
rect -1130 -4492 -1100 -4292
rect -911 -4420 -881 -4292
rect -814 -4492 -784 -4292
rect -615 -4426 -585 -4298
rect -531 -4426 -501 -4298
rect -264 -4376 -234 -4292
rect -172 -4376 -142 -4292
rect -73 -4376 -43 -4292
rect 67 -4376 97 -4292
rect 164 -4376 194 -4292
rect 361 -4460 391 -4292
rect 460 -4376 490 -4292
rect 546 -4376 576 -4292
rect 630 -4376 660 -4292
rect 738 -4376 768 -4292
rect 822 -4376 852 -4292
rect 986 -4492 1016 -4292
rect 1205 -4420 1235 -4292
rect 1302 -4492 1332 -4292
rect 1501 -4426 1531 -4298
rect 1585 -4426 1615 -4298
rect 1852 -4376 1882 -4292
rect 1944 -4376 1974 -4292
rect 2043 -4376 2073 -4292
rect 2183 -4376 2213 -4292
rect 2280 -4376 2310 -4292
rect 2477 -4460 2507 -4292
rect 2576 -4376 2606 -4292
rect 2662 -4376 2692 -4292
rect 2746 -4376 2776 -4292
rect 2854 -4376 2884 -4292
rect 2938 -4376 2968 -4292
rect 3102 -4492 3132 -4292
rect 3321 -4420 3351 -4292
rect 3418 -4492 3448 -4292
rect 3617 -4426 3647 -4298
rect 3701 -4426 3731 -4298
rect 3968 -4376 3998 -4292
rect 4060 -4376 4090 -4292
rect 4159 -4376 4189 -4292
rect 4299 -4376 4329 -4292
rect 4396 -4376 4426 -4292
rect 4593 -4460 4623 -4292
rect 4692 -4376 4722 -4292
rect 4778 -4376 4808 -4292
rect 4862 -4376 4892 -4292
rect 4970 -4376 5000 -4292
rect 5054 -4376 5084 -4292
rect 5218 -4492 5248 -4292
rect 5437 -4420 5467 -4292
rect 5534 -4492 5564 -4292
rect 5733 -4426 5763 -4298
rect 5817 -4426 5847 -4298
rect 6084 -4376 6114 -4292
rect 6176 -4376 6206 -4292
rect 6275 -4376 6305 -4292
rect 6415 -4376 6445 -4292
rect 6512 -4376 6542 -4292
rect 6709 -4460 6739 -4292
rect 6808 -4376 6838 -4292
rect 6894 -4376 6924 -4292
rect 6978 -4376 7008 -4292
rect 7086 -4376 7116 -4292
rect 7170 -4376 7200 -4292
rect 7334 -4492 7364 -4292
rect 7553 -4420 7583 -4292
rect 7650 -4492 7680 -4292
rect 7849 -4426 7879 -4298
rect 7933 -4426 7963 -4298
rect 8200 -4376 8230 -4292
rect 8292 -4376 8322 -4292
rect 8391 -4376 8421 -4292
rect 8531 -4376 8561 -4292
rect 8628 -4376 8658 -4292
rect 8825 -4460 8855 -4292
rect 8924 -4376 8954 -4292
rect 9010 -4376 9040 -4292
rect 9094 -4376 9124 -4292
rect 9202 -4376 9232 -4292
rect 9286 -4376 9316 -4292
rect 9450 -4492 9480 -4292
rect 9669 -4420 9699 -4292
rect 9766 -4492 9796 -4292
rect 9965 -4426 9995 -4298
rect 10049 -4426 10079 -4298
rect 10316 -4376 10346 -4292
rect 10408 -4376 10438 -4292
rect 10507 -4376 10537 -4292
rect 10647 -4376 10677 -4292
rect 10744 -4376 10774 -4292
rect 10941 -4460 10971 -4292
rect 11040 -4376 11070 -4292
rect 11126 -4376 11156 -4292
rect 11210 -4376 11240 -4292
rect 11318 -4376 11348 -4292
rect 11402 -4376 11432 -4292
rect 11566 -4492 11596 -4292
rect 11785 -4420 11815 -4292
rect 11882 -4492 11912 -4292
rect 12081 -4426 12111 -4298
rect 12165 -4426 12195 -4298
rect 12432 -4376 12462 -4292
rect 12524 -4376 12554 -4292
rect 12623 -4376 12653 -4292
rect 12763 -4376 12793 -4292
rect 12860 -4376 12890 -4292
rect 13057 -4460 13087 -4292
rect 13156 -4376 13186 -4292
rect 13242 -4376 13272 -4292
rect 13326 -4376 13356 -4292
rect 13434 -4376 13464 -4292
rect 13518 -4376 13548 -4292
rect 13682 -4492 13712 -4292
rect 13901 -4420 13931 -4292
rect 13998 -4492 14028 -4292
rect 14197 -4426 14227 -4298
rect 14281 -4426 14311 -4298
rect 14548 -4376 14578 -4292
rect 14640 -4376 14670 -4292
rect 14739 -4376 14769 -4292
rect 14879 -4376 14909 -4292
rect 14976 -4376 15006 -4292
rect 15173 -4460 15203 -4292
rect 15272 -4376 15302 -4292
rect 15358 -4376 15388 -4292
rect 15442 -4376 15472 -4292
rect 15550 -4376 15580 -4292
rect 15634 -4376 15664 -4292
rect 15798 -4492 15828 -4292
rect 16017 -4420 16047 -4292
rect 16114 -4492 16144 -4292
rect 16313 -4426 16343 -4298
rect 16397 -4426 16427 -4298
rect 16664 -4376 16694 -4292
rect 16756 -4376 16786 -4292
rect 16855 -4376 16885 -4292
rect 16995 -4376 17025 -4292
rect 17092 -4376 17122 -4292
rect 17289 -4460 17319 -4292
rect 17388 -4376 17418 -4292
rect 17474 -4376 17504 -4292
rect 17558 -4376 17588 -4292
rect 17666 -4376 17696 -4292
rect 17750 -4376 17780 -4292
rect 17914 -4492 17944 -4292
rect 18133 -4420 18163 -4292
rect 18230 -4492 18260 -4292
rect 18429 -4426 18459 -4298
rect 18513 -4426 18543 -4298
rect 18780 -4376 18810 -4292
rect 18872 -4376 18902 -4292
rect 18971 -4376 19001 -4292
rect 19111 -4376 19141 -4292
rect 19208 -4376 19238 -4292
rect 19405 -4460 19435 -4292
rect 19504 -4376 19534 -4292
rect 19590 -4376 19620 -4292
rect 19674 -4376 19704 -4292
rect 19782 -4376 19812 -4292
rect 19866 -4376 19896 -4292
rect 20030 -4492 20060 -4292
rect 20249 -4420 20279 -4292
rect 20346 -4492 20376 -4292
rect 20545 -4426 20575 -4298
rect 20629 -4426 20659 -4298
rect 20896 -4376 20926 -4292
rect 20988 -4376 21018 -4292
rect 21087 -4376 21117 -4292
rect 21227 -4376 21257 -4292
rect 21324 -4376 21354 -4292
rect 21521 -4460 21551 -4292
rect 21620 -4376 21650 -4292
rect 21706 -4376 21736 -4292
rect 21790 -4376 21820 -4292
rect 21898 -4376 21928 -4292
rect 21982 -4376 22012 -4292
rect 22146 -4492 22176 -4292
rect 22365 -4420 22395 -4292
rect 22462 -4492 22492 -4292
rect 22661 -4426 22691 -4298
rect 22745 -4426 22775 -4298
rect 23012 -4376 23042 -4292
rect 23104 -4376 23134 -4292
rect 23203 -4376 23233 -4292
rect 23343 -4376 23373 -4292
rect 23440 -4376 23470 -4292
rect 23637 -4460 23667 -4292
rect 23736 -4376 23766 -4292
rect 23822 -4376 23852 -4292
rect 23906 -4376 23936 -4292
rect 24014 -4376 24044 -4292
rect 24098 -4376 24128 -4292
rect 24262 -4492 24292 -4292
rect 24481 -4420 24511 -4292
rect 24578 -4492 24608 -4292
rect 24777 -4426 24807 -4298
rect 24861 -4426 24891 -4298
rect 25128 -4376 25158 -4292
rect 25220 -4376 25250 -4292
rect 25319 -4376 25349 -4292
rect 25459 -4376 25489 -4292
rect 25556 -4376 25586 -4292
rect 25753 -4460 25783 -4292
rect 25852 -4376 25882 -4292
rect 25938 -4376 25968 -4292
rect 26022 -4376 26052 -4292
rect 26130 -4376 26160 -4292
rect 26214 -4376 26244 -4292
rect 26378 -4492 26408 -4292
rect 26597 -4420 26627 -4292
rect 26694 -4492 26724 -4292
rect 26893 -4426 26923 -4298
rect 26977 -4426 27007 -4298
rect 27244 -4376 27274 -4292
rect 27336 -4376 27366 -4292
rect 27435 -4376 27465 -4292
rect 27575 -4376 27605 -4292
rect 27672 -4376 27702 -4292
rect 27869 -4460 27899 -4292
rect 27968 -4376 27998 -4292
rect 28054 -4376 28084 -4292
rect 28138 -4376 28168 -4292
rect 28246 -4376 28276 -4292
rect 28330 -4376 28360 -4292
rect 28494 -4492 28524 -4292
rect 28713 -4420 28743 -4292
rect 28810 -4492 28840 -4292
rect 29009 -4426 29039 -4298
rect 29093 -4426 29123 -4298
rect 29360 -4376 29390 -4292
rect 29452 -4376 29482 -4292
rect 29551 -4376 29581 -4292
rect 29691 -4376 29721 -4292
rect 29788 -4376 29818 -4292
rect 29985 -4460 30015 -4292
rect 30084 -4376 30114 -4292
rect 30170 -4376 30200 -4292
rect 30254 -4376 30284 -4292
rect 30362 -4376 30392 -4292
rect 30446 -4376 30476 -4292
rect 30610 -4492 30640 -4292
rect 30829 -4420 30859 -4292
rect 30926 -4492 30956 -4292
rect 31125 -4426 31155 -4298
rect 31209 -4426 31239 -4298
rect 31476 -4376 31506 -4292
rect 31568 -4376 31598 -4292
rect 31667 -4376 31697 -4292
rect 31807 -4376 31837 -4292
rect 31904 -4376 31934 -4292
rect 32101 -4460 32131 -4292
rect 32200 -4376 32230 -4292
rect 32286 -4376 32316 -4292
rect 32370 -4376 32400 -4292
rect 32478 -4376 32508 -4292
rect 32562 -4376 32592 -4292
rect 32726 -4492 32756 -4292
rect 32945 -4420 32975 -4292
rect 33042 -4492 33072 -4292
<< pmoslvt >>
rect -94564 19168 -92964 20568
rect -92906 19168 -91306 20568
rect -91248 19168 -89648 20568
rect -89590 19168 -87990 20568
rect -87932 19168 -86332 20568
rect -86274 19168 -84674 20568
rect -84616 19168 -83016 20568
rect -82958 19168 -81358 20568
rect -81300 19168 -79700 20568
rect -79642 19168 -78042 20568
rect -77984 19168 -76384 20568
rect -76326 19168 -74726 20568
rect -74668 19168 -73068 20568
rect -73010 19168 -71410 20568
rect -71352 19168 -69752 20568
rect -69694 19168 -68094 20568
rect -68036 19168 -66436 20568
rect -66378 19168 -64778 20568
rect -64720 19168 -63120 20568
rect -63062 19168 -61462 20568
rect -61404 19168 -59804 20568
rect -59746 19168 -58146 20568
rect -58088 19168 -56488 20568
rect -56430 19168 -54830 20568
rect -54772 19168 -53172 20568
rect -53114 19168 -51514 20568
rect -51456 19168 -49856 20568
rect -49798 19168 -48198 20568
rect -48140 19168 -46540 20568
rect -46482 19168 -44882 20568
rect -44824 19168 -43224 20568
rect -43166 19168 -41566 20568
rect -41508 19168 -39908 20568
rect -39850 19168 -38250 20568
rect -38192 19168 -36592 20568
rect -36534 19168 -34934 20568
rect -34876 19168 -33276 20568
rect -33218 19168 -31618 20568
rect -31560 19168 -29960 20568
rect -29902 19168 -28302 20568
rect -94564 17532 -92964 18932
rect -92906 17532 -91306 18932
rect -91248 17532 -89648 18932
rect -89590 17532 -87990 18932
rect -87932 17532 -86332 18932
rect -86274 17532 -84674 18932
rect -84616 17532 -83016 18932
rect -82958 17532 -81358 18932
rect -81300 17532 -79700 18932
rect -79642 17532 -78042 18932
rect -77984 17532 -76384 18932
rect -76326 17532 -74726 18932
rect -74668 17532 -73068 18932
rect -73010 17532 -71410 18932
rect -71352 17532 -69752 18932
rect -69694 17532 -68094 18932
rect -68036 17532 -66436 18932
rect -66378 17532 -64778 18932
rect -64720 17532 -63120 18932
rect -63062 17532 -61462 18932
rect -61404 17532 -59804 18932
rect -59746 17532 -58146 18932
rect -58088 17532 -56488 18932
rect -56430 17532 -54830 18932
rect -54772 17532 -53172 18932
rect -53114 17532 -51514 18932
rect -51456 17532 -49856 18932
rect -49798 17532 -48198 18932
rect -48140 17532 -46540 18932
rect -46482 17532 -44882 18932
rect -44824 17532 -43224 18932
rect -43166 17532 -41566 18932
rect -41508 17532 -39908 18932
rect -39850 17532 -38250 18932
rect -38192 17532 -36592 18932
rect -36534 17532 -34934 18932
rect -34876 17532 -33276 18932
rect -33218 17532 -31618 18932
rect -31560 17532 -29960 18932
rect -29902 17532 -28302 18932
rect -94562 15786 -92962 17186
rect -92904 15786 -91304 17186
rect -91246 15786 -89646 17186
rect -89588 15786 -87988 17186
rect -87930 15786 -86330 17186
rect -86272 15786 -84672 17186
rect -84614 15786 -83014 17186
rect -82956 15786 -81356 17186
rect -81298 15786 -79698 17186
rect -79640 15786 -78040 17186
rect -77982 15786 -76382 17186
rect -76324 15786 -74724 17186
rect -74666 15786 -73066 17186
rect -73008 15786 -71408 17186
rect -71350 15786 -69750 17186
rect -69692 15786 -68092 17186
rect -68034 15786 -66434 17186
rect -66376 15786 -64776 17186
rect -64718 15786 -63118 17186
rect -63060 15786 -61460 17186
rect -61402 15786 -59802 17186
rect -59744 15786 -58144 17186
rect -58086 15786 -56486 17186
rect -56428 15786 -54828 17186
rect -54770 15786 -53170 17186
rect -53112 15786 -51512 17186
rect -51454 15786 -49854 17186
rect -49796 15786 -48196 17186
rect -48138 15786 -46538 17186
rect -46480 15786 -44880 17186
rect -44822 15786 -43222 17186
rect -43164 15786 -41564 17186
rect -41506 15786 -39906 17186
rect -39848 15786 -38248 17186
rect -38190 15786 -36590 17186
rect -36532 15786 -34932 17186
rect -34874 15786 -33274 17186
rect -33216 15786 -31616 17186
rect -31558 15786 -29958 17186
rect -29900 15786 -28300 17186
rect -94562 14150 -92962 15550
rect -92904 14150 -91304 15550
rect -91246 14150 -89646 15550
rect -89588 14150 -87988 15550
rect -87930 14150 -86330 15550
rect -86272 14150 -84672 15550
rect -84614 14150 -83014 15550
rect -82956 14150 -81356 15550
rect -81298 14150 -79698 15550
rect -79640 14150 -78040 15550
rect -77982 14150 -76382 15550
rect -76324 14150 -74724 15550
rect -74666 14150 -73066 15550
rect -73008 14150 -71408 15550
rect -71350 14150 -69750 15550
rect -69692 14150 -68092 15550
rect -68034 14150 -66434 15550
rect -66376 14150 -64776 15550
rect -64718 14150 -63118 15550
rect -63060 14150 -61460 15550
rect -61402 14150 -59802 15550
rect -59744 14150 -58144 15550
rect -58086 14150 -56486 15550
rect -56428 14150 -54828 15550
rect -54770 14150 -53170 15550
rect -53112 14150 -51512 15550
rect -51454 14150 -49854 15550
rect -49796 14150 -48196 15550
rect -48138 14150 -46538 15550
rect -46480 14150 -44880 15550
rect -44822 14150 -43222 15550
rect -43164 14150 -41564 15550
rect -41506 14150 -39906 15550
rect -39848 14150 -38248 15550
rect -38190 14150 -36590 15550
rect -36532 14150 -34932 15550
rect -34874 14150 -33274 15550
rect -33216 14150 -31616 15550
rect -31558 14150 -29958 15550
rect -29900 14150 -28300 15550
rect -94562 12514 -92962 13914
rect -92904 12514 -91304 13914
rect -91246 12514 -89646 13914
rect -89588 12514 -87988 13914
rect -87930 12514 -86330 13914
rect -86272 12514 -84672 13914
rect -84614 12514 -83014 13914
rect -82956 12514 -81356 13914
rect -81298 12514 -79698 13914
rect -79640 12514 -78040 13914
rect -77982 12514 -76382 13914
rect -76324 12514 -74724 13914
rect -74666 12514 -73066 13914
rect -73008 12514 -71408 13914
rect -71350 12514 -69750 13914
rect -69692 12514 -68092 13914
rect -68034 12514 -66434 13914
rect -66376 12514 -64776 13914
rect -64718 12514 -63118 13914
rect -63060 12514 -61460 13914
rect -61402 12514 -59802 13914
rect -59744 12514 -58144 13914
rect -58086 12514 -56486 13914
rect -56428 12514 -54828 13914
rect -54770 12514 -53170 13914
rect -53112 12514 -51512 13914
rect -51454 12514 -49854 13914
rect -49796 12514 -48196 13914
rect -48138 12514 -46538 13914
rect -46480 12514 -44880 13914
rect -44822 12514 -43222 13914
rect -43164 12514 -41564 13914
rect -41506 12514 -39906 13914
rect -39848 12514 -38248 13914
rect -38190 12514 -36590 13914
rect -36532 12514 -34932 13914
rect -34874 12514 -33274 13914
rect -33216 12514 -31616 13914
rect -31558 12514 -29958 13914
rect -29900 12514 -28300 13914
rect -94562 10878 -92962 12278
rect -92904 10878 -91304 12278
rect -91246 10878 -89646 12278
rect -89588 10878 -87988 12278
rect -87930 10878 -86330 12278
rect -86272 10878 -84672 12278
rect -84614 10878 -83014 12278
rect -82956 10878 -81356 12278
rect -81298 10878 -79698 12278
rect -79640 10878 -78040 12278
rect -77982 10878 -76382 12278
rect -76324 10878 -74724 12278
rect -74666 10878 -73066 12278
rect -73008 10878 -71408 12278
rect -71350 10878 -69750 12278
rect -69692 10878 -68092 12278
rect -68034 10878 -66434 12278
rect -66376 10878 -64776 12278
rect -64718 10878 -63118 12278
rect -63060 10878 -61460 12278
rect -61402 10878 -59802 12278
rect -59744 10878 -58144 12278
rect -58086 10878 -56486 12278
rect -56428 10878 -54828 12278
rect -54770 10878 -53170 12278
rect -53112 10878 -51512 12278
rect -51454 10878 -49854 12278
rect -49796 10878 -48196 12278
rect -48138 10878 -46538 12278
rect -46480 10878 -44880 12278
rect -44822 10878 -43222 12278
rect -43164 10878 -41564 12278
rect -41506 10878 -39906 12278
rect -39848 10878 -38248 12278
rect -38190 10878 -36590 12278
rect -36532 10878 -34932 12278
rect -34874 10878 -33274 12278
rect -33216 10878 -31616 12278
rect -31558 10878 -29958 12278
rect -29900 10878 -28300 12278
rect -94562 9240 -92962 10640
rect -92904 9240 -91304 10640
rect -91246 9240 -89646 10640
rect -89588 9240 -87988 10640
rect -87930 9240 -86330 10640
rect -86272 9240 -84672 10640
rect -84614 9240 -83014 10640
rect -82956 9240 -81356 10640
rect -81298 9240 -79698 10640
rect -79640 9240 -78040 10640
rect -77982 9240 -76382 10640
rect -76324 9240 -74724 10640
rect -74666 9240 -73066 10640
rect -73008 9240 -71408 10640
rect -71350 9240 -69750 10640
rect -69692 9240 -68092 10640
rect -68034 9240 -66434 10640
rect -66376 9240 -64776 10640
rect -64718 9240 -63118 10640
rect -63060 9240 -61460 10640
rect -61402 9240 -59802 10640
rect -59744 9240 -58144 10640
rect -58086 9240 -56486 10640
rect -56428 9240 -54828 10640
rect -54770 9240 -53170 10640
rect -53112 9240 -51512 10640
rect -51454 9240 -49854 10640
rect -49796 9240 -48196 10640
rect -48138 9240 -46538 10640
rect -46480 9240 -44880 10640
rect -44822 9240 -43222 10640
rect -43164 9240 -41564 10640
rect -41506 9240 -39906 10640
rect -39848 9240 -38248 10640
rect -38190 9240 -36590 10640
rect -36532 9240 -34932 10640
rect -34874 9240 -33274 10640
rect -33216 9240 -31616 10640
rect -31558 9240 -29958 10640
rect -29900 9240 -28300 10640
rect -94562 7604 -92962 9004
rect -92904 7604 -91304 9004
rect -91246 7604 -89646 9004
rect -89588 7604 -87988 9004
rect -87930 7604 -86330 9004
rect -86272 7604 -84672 9004
rect -84614 7604 -83014 9004
rect -82956 7604 -81356 9004
rect -81298 7604 -79698 9004
rect -79640 7604 -78040 9004
rect -77982 7604 -76382 9004
rect -76324 7604 -74724 9004
rect -74666 7604 -73066 9004
rect -73008 7604 -71408 9004
rect -71350 7604 -69750 9004
rect -69692 7604 -68092 9004
rect -68034 7604 -66434 9004
rect -66376 7604 -64776 9004
rect -64718 7604 -63118 9004
rect -63060 7604 -61460 9004
rect -61402 7604 -59802 9004
rect -59744 7604 -58144 9004
rect -58086 7604 -56486 9004
rect -56428 7604 -54828 9004
rect -54770 7604 -53170 9004
rect -53112 7604 -51512 9004
rect -51454 7604 -49854 9004
rect -49796 7604 -48196 9004
rect -48138 7604 -46538 9004
rect -46480 7604 -44880 9004
rect -44822 7604 -43222 9004
rect -43164 7604 -41564 9004
rect -41506 7604 -39906 9004
rect -39848 7604 -38248 9004
rect -38190 7604 -36590 9004
rect -36532 7604 -34932 9004
rect -34874 7604 -33274 9004
rect -33216 7604 -31616 9004
rect -31558 7604 -29958 9004
rect -29900 7604 -28300 9004
rect -94562 5968 -92962 7368
rect -92904 5968 -91304 7368
rect -91246 5968 -89646 7368
rect -89588 5968 -87988 7368
rect -87930 5968 -86330 7368
rect -86272 5968 -84672 7368
rect -84614 5968 -83014 7368
rect -82956 5968 -81356 7368
rect -81298 5968 -79698 7368
rect -79640 5968 -78040 7368
rect -77982 5968 -76382 7368
rect -76324 5968 -74724 7368
rect -74666 5968 -73066 7368
rect -73008 5968 -71408 7368
rect -71350 5968 -69750 7368
rect -69692 5968 -68092 7368
rect -68034 5968 -66434 7368
rect -66376 5968 -64776 7368
rect -64718 5968 -63118 7368
rect -63060 5968 -61460 7368
rect -61402 5968 -59802 7368
rect -59744 5968 -58144 7368
rect -58086 5968 -56486 7368
rect -56428 5968 -54828 7368
rect -54770 5968 -53170 7368
rect -53112 5968 -51512 7368
rect -51454 5968 -49854 7368
rect -49796 5968 -48196 7368
rect -48138 5968 -46538 7368
rect -46480 5968 -44880 7368
rect -44822 5968 -43222 7368
rect -43164 5968 -41564 7368
rect -41506 5968 -39906 7368
rect -39848 5968 -38248 7368
rect -38190 5968 -36590 7368
rect -36532 5968 -34932 7368
rect -34874 5968 -33274 7368
rect -33216 5968 -31616 7368
rect -31558 5968 -29958 7368
rect -29900 5968 -28300 7368
rect -94562 4332 -92962 5732
rect -92904 4332 -91304 5732
rect -91246 4332 -89646 5732
rect -89588 4332 -87988 5732
rect -87930 4332 -86330 5732
rect -86272 4332 -84672 5732
rect -84614 4332 -83014 5732
rect -82956 4332 -81356 5732
rect -81298 4332 -79698 5732
rect -79640 4332 -78040 5732
rect -77982 4332 -76382 5732
rect -76324 4332 -74724 5732
rect -74666 4332 -73066 5732
rect -73008 4332 -71408 5732
rect -71350 4332 -69750 5732
rect -69692 4332 -68092 5732
rect -68034 4332 -66434 5732
rect -66376 4332 -64776 5732
rect -64718 4332 -63118 5732
rect -63060 4332 -61460 5732
rect -61402 4332 -59802 5732
rect -59744 4332 -58144 5732
rect -58086 4332 -56486 5732
rect -56428 4332 -54828 5732
rect -54770 4332 -53170 5732
rect -53112 4332 -51512 5732
rect -51454 4332 -49854 5732
rect -49796 4332 -48196 5732
rect -48138 4332 -46538 5732
rect -46480 4332 -44880 5732
rect -44822 4332 -43222 5732
rect -43164 4332 -41564 5732
rect -41506 4332 -39906 5732
rect -39848 4332 -38248 5732
rect -38190 4332 -36590 5732
rect -36532 4332 -34932 5732
rect -34874 4332 -33274 5732
rect -33216 4332 -31616 5732
rect -31558 4332 -29958 5732
rect -29900 4332 -28300 5732
rect 2666 4916 2866 5916
rect 3322 4924 3522 5924
rect 3580 4924 3780 5924
rect 4322 4924 4522 5924
rect 4580 4924 4780 5924
rect 5228 4928 5428 5928
rect 8602 4656 8802 5656
rect 9081 4648 9281 5648
rect 9339 4648 9539 5648
rect 9739 4650 9939 5650
rect 9997 4650 10197 5650
rect 10396 4630 10596 5630
rect 13876 4528 14076 5528
rect 14270 4510 14670 5510
rect 14842 4510 15242 5510
rect 15464 4540 15664 5540
rect 9433 -7875 9633 -7675
rect 10093 -7875 10293 -7675
rect 10563 -7875 10763 -7675
rect 11166 -7876 11366 -7676
rect 11424 -7876 11624 -7676
rect 11682 -7876 11882 -7676
rect 11940 -7876 12140 -7676
rect 12198 -7876 12398 -7676
rect 12981 -7876 13181 -7676
rect 13239 -7876 13439 -7676
rect 13497 -7876 13697 -7676
rect 13755 -7876 13955 -7676
rect 14013 -7876 14213 -7676
rect 14787 -7876 14987 -7676
rect 15045 -7876 15245 -7676
rect 15303 -7876 15503 -7676
rect 15561 -7876 15761 -7676
rect 15819 -7876 16019 -7676
rect 9737 -8759 10537 -8649
rect 12407 -8759 13207 -8649
rect 15070 -8758 15870 -8648
rect 9729 -14441 10529 -14331
rect 12406 -14441 13206 -14331
rect 15070 -14440 15870 -14330
rect 9737 -20366 10537 -20256
rect 12407 -20366 13207 -20256
rect 15070 -20365 15870 -20255
<< nmoslvt >>
rect 8832 3284 9032 3684
rect 9090 3284 9290 3684
rect 9348 3284 9548 3684
rect 9846 3284 10046 3684
rect 10104 3284 10304 3684
rect 10362 3284 10562 3684
rect 8832 2728 9032 3128
rect 9090 2728 9290 3128
rect 9348 2728 9548 3128
rect 9846 2728 10046 3128
rect 10104 2728 10304 3128
rect 10362 2728 10562 3128
rect 2672 2332 2872 2532
rect 3148 2334 3948 2534
rect 4120 2334 4920 2534
rect 5206 2332 5406 2532
rect 9153 1684 9553 1884
rect 9748 1684 10148 1884
rect 13364 314 13564 3114
rect 13914 2180 14114 2980
rect 14172 2180 14372 2980
rect 14430 2180 14630 2980
rect 14914 2180 15114 2980
rect 15172 2180 15372 2980
rect 15430 2180 15630 2980
rect 13914 1224 14114 2024
rect 14172 1224 14372 2024
rect 14430 1224 14630 2024
rect 14914 1224 15114 2024
rect 15172 1224 15372 2024
rect 15430 1224 15630 2024
rect 13914 268 14114 1068
rect 14172 268 14372 1068
rect 14430 268 14630 1068
rect 14914 268 15114 1068
rect 15172 268 15372 1068
rect 15430 268 15630 1068
rect 15962 264 16162 3064
rect 9159 -9836 9359 -9636
rect 9417 -9836 9617 -9636
rect 9675 -9836 9875 -9636
rect 9933 -9836 10133 -9636
rect 10191 -9836 10391 -9636
rect 10449 -9836 10649 -9636
rect 10707 -9836 10907 -9636
rect 10965 -9836 11165 -9636
rect 11829 -9836 12029 -9636
rect 12087 -9836 12287 -9636
rect 12345 -9836 12545 -9636
rect 12603 -9836 12803 -9636
rect 12861 -9836 13061 -9636
rect 13119 -9836 13319 -9636
rect 13377 -9836 13577 -9636
rect 13635 -9836 13835 -9636
rect 14492 -9835 14692 -9635
rect 14750 -9835 14950 -9635
rect 15008 -9835 15208 -9635
rect 15266 -9835 15466 -9635
rect 15524 -9835 15724 -9635
rect 15782 -9835 15982 -9635
rect 16040 -9835 16240 -9635
rect 16298 -9835 16498 -9635
rect 9159 -10254 9359 -10054
rect 9417 -10254 9617 -10054
rect 9675 -10254 9875 -10054
rect 9933 -10254 10133 -10054
rect 10191 -10254 10391 -10054
rect 10449 -10254 10649 -10054
rect 10707 -10254 10907 -10054
rect 10965 -10254 11165 -10054
rect 11829 -10254 12029 -10054
rect 12087 -10254 12287 -10054
rect 12345 -10254 12545 -10054
rect 12603 -10254 12803 -10054
rect 12861 -10254 13061 -10054
rect 13119 -10254 13319 -10054
rect 13377 -10254 13577 -10054
rect 13635 -10254 13835 -10054
rect 14492 -10253 14692 -10053
rect 14750 -10253 14950 -10053
rect 15008 -10253 15208 -10053
rect 15266 -10253 15466 -10053
rect 15524 -10253 15724 -10053
rect 15782 -10253 15982 -10053
rect 16040 -10253 16240 -10053
rect 16298 -10253 16498 -10053
rect 9159 -10672 9359 -10472
rect 9417 -10672 9617 -10472
rect 9675 -10672 9875 -10472
rect 9933 -10672 10133 -10472
rect 10191 -10672 10391 -10472
rect 10449 -10672 10649 -10472
rect 10707 -10672 10907 -10472
rect 10965 -10672 11165 -10472
rect 11829 -10672 12029 -10472
rect 12087 -10672 12287 -10472
rect 12345 -10672 12545 -10472
rect 12603 -10672 12803 -10472
rect 12861 -10672 13061 -10472
rect 13119 -10672 13319 -10472
rect 13377 -10672 13577 -10472
rect 13635 -10672 13835 -10472
rect 14492 -10671 14692 -10471
rect 14750 -10671 14950 -10471
rect 15008 -10671 15208 -10471
rect 15266 -10671 15466 -10471
rect 15524 -10671 15724 -10471
rect 15782 -10671 15982 -10471
rect 16040 -10671 16240 -10471
rect 16298 -10671 16498 -10471
rect 9159 -11090 9359 -10890
rect 9417 -11090 9617 -10890
rect 9675 -11090 9875 -10890
rect 9933 -11090 10133 -10890
rect 10191 -11090 10391 -10890
rect 10449 -11090 10649 -10890
rect 10707 -11090 10907 -10890
rect 10965 -11090 11165 -10890
rect 11829 -11090 12029 -10890
rect 12087 -11090 12287 -10890
rect 12345 -11090 12545 -10890
rect 12603 -11090 12803 -10890
rect 12861 -11090 13061 -10890
rect 13119 -11090 13319 -10890
rect 13377 -11090 13577 -10890
rect 13635 -11090 13835 -10890
rect 14492 -11089 14692 -10889
rect 14750 -11089 14950 -10889
rect 15008 -11089 15208 -10889
rect 15266 -11089 15466 -10889
rect 15524 -11089 15724 -10889
rect 15782 -11089 15982 -10889
rect 16040 -11089 16240 -10889
rect 16298 -11089 16498 -10889
rect 9159 -11508 9359 -11308
rect 9417 -11508 9617 -11308
rect 9675 -11508 9875 -11308
rect 9933 -11508 10133 -11308
rect 10191 -11508 10391 -11308
rect 10449 -11508 10649 -11308
rect 10707 -11508 10907 -11308
rect 10965 -11508 11165 -11308
rect 11829 -11508 12029 -11308
rect 12087 -11508 12287 -11308
rect 12345 -11508 12545 -11308
rect 12603 -11508 12803 -11308
rect 12861 -11508 13061 -11308
rect 13119 -11508 13319 -11308
rect 13377 -11508 13577 -11308
rect 13635 -11508 13835 -11308
rect 14492 -11507 14692 -11307
rect 14750 -11507 14950 -11307
rect 15008 -11507 15208 -11307
rect 15266 -11507 15466 -11307
rect 15524 -11507 15724 -11307
rect 15782 -11507 15982 -11307
rect 16040 -11507 16240 -11307
rect 16298 -11507 16498 -11307
rect 9159 -11926 9359 -11726
rect 9417 -11926 9617 -11726
rect 9675 -11926 9875 -11726
rect 9933 -11926 10133 -11726
rect 10191 -11926 10391 -11726
rect 10449 -11926 10649 -11726
rect 10707 -11926 10907 -11726
rect 10965 -11926 11165 -11726
rect 11829 -11926 12029 -11726
rect 12087 -11926 12287 -11726
rect 12345 -11926 12545 -11726
rect 12603 -11926 12803 -11726
rect 12861 -11926 13061 -11726
rect 13119 -11926 13319 -11726
rect 13377 -11926 13577 -11726
rect 13635 -11926 13835 -11726
rect 14492 -11925 14692 -11725
rect 14750 -11925 14950 -11725
rect 15008 -11925 15208 -11725
rect 15266 -11925 15466 -11725
rect 15524 -11925 15724 -11725
rect 15782 -11925 15982 -11725
rect 16040 -11925 16240 -11725
rect 16298 -11925 16498 -11725
rect 9159 -12344 9359 -12144
rect 9417 -12344 9617 -12144
rect 9675 -12344 9875 -12144
rect 9933 -12344 10133 -12144
rect 10191 -12344 10391 -12144
rect 10449 -12344 10649 -12144
rect 10707 -12344 10907 -12144
rect 10965 -12344 11165 -12144
rect 11829 -12344 12029 -12144
rect 12087 -12344 12287 -12144
rect 12345 -12344 12545 -12144
rect 12603 -12344 12803 -12144
rect 12861 -12344 13061 -12144
rect 13119 -12344 13319 -12144
rect 13377 -12344 13577 -12144
rect 13635 -12344 13835 -12144
rect 14492 -12343 14692 -12143
rect 14750 -12343 14950 -12143
rect 15008 -12343 15208 -12143
rect 15266 -12343 15466 -12143
rect 15524 -12343 15724 -12143
rect 15782 -12343 15982 -12143
rect 16040 -12343 16240 -12143
rect 16298 -12343 16498 -12143
rect 9039 -12996 9239 -12796
rect 9579 -12996 9779 -12796
rect 10059 -12996 10259 -12796
rect 10562 -12994 10762 -12794
rect 11072 -12984 11272 -12784
rect 11709 -12996 11909 -12796
rect 12249 -12996 12449 -12796
rect 12729 -12996 12929 -12796
rect 13232 -12994 13432 -12794
rect 13742 -12984 13942 -12784
rect 14372 -12995 14572 -12795
rect 14912 -12995 15112 -12795
rect 15392 -12995 15592 -12795
rect 15895 -12993 16095 -12793
rect 16405 -12983 16605 -12783
rect 9159 -15553 9359 -15353
rect 9417 -15553 9617 -15353
rect 9675 -15553 9875 -15353
rect 9933 -15553 10133 -15353
rect 10191 -15553 10391 -15353
rect 10449 -15553 10649 -15353
rect 10707 -15553 10907 -15353
rect 10965 -15553 11165 -15353
rect 11829 -15553 12029 -15353
rect 12087 -15553 12287 -15353
rect 12345 -15553 12545 -15353
rect 12603 -15553 12803 -15353
rect 12861 -15553 13061 -15353
rect 13119 -15553 13319 -15353
rect 13377 -15553 13577 -15353
rect 13635 -15553 13835 -15353
rect 14492 -15552 14692 -15352
rect 14750 -15552 14950 -15352
rect 15008 -15552 15208 -15352
rect 15266 -15552 15466 -15352
rect 15524 -15552 15724 -15352
rect 15782 -15552 15982 -15352
rect 16040 -15552 16240 -15352
rect 16298 -15552 16498 -15352
rect 9159 -15971 9359 -15771
rect 9417 -15971 9617 -15771
rect 9675 -15971 9875 -15771
rect 9933 -15971 10133 -15771
rect 10191 -15971 10391 -15771
rect 10449 -15971 10649 -15771
rect 10707 -15971 10907 -15771
rect 10965 -15971 11165 -15771
rect 11829 -15971 12029 -15771
rect 12087 -15971 12287 -15771
rect 12345 -15971 12545 -15771
rect 12603 -15971 12803 -15771
rect 12861 -15971 13061 -15771
rect 13119 -15971 13319 -15771
rect 13377 -15971 13577 -15771
rect 13635 -15971 13835 -15771
rect 14492 -15970 14692 -15770
rect 14750 -15970 14950 -15770
rect 15008 -15970 15208 -15770
rect 15266 -15970 15466 -15770
rect 15524 -15970 15724 -15770
rect 15782 -15970 15982 -15770
rect 16040 -15970 16240 -15770
rect 16298 -15970 16498 -15770
rect 9159 -16389 9359 -16189
rect 9417 -16389 9617 -16189
rect 9675 -16389 9875 -16189
rect 9933 -16389 10133 -16189
rect 10191 -16389 10391 -16189
rect 10449 -16389 10649 -16189
rect 10707 -16389 10907 -16189
rect 10965 -16389 11165 -16189
rect 11829 -16389 12029 -16189
rect 12087 -16389 12287 -16189
rect 12345 -16389 12545 -16189
rect 12603 -16389 12803 -16189
rect 12861 -16389 13061 -16189
rect 13119 -16389 13319 -16189
rect 13377 -16389 13577 -16189
rect 13635 -16389 13835 -16189
rect 14492 -16388 14692 -16188
rect 14750 -16388 14950 -16188
rect 15008 -16388 15208 -16188
rect 15266 -16388 15466 -16188
rect 15524 -16388 15724 -16188
rect 15782 -16388 15982 -16188
rect 16040 -16388 16240 -16188
rect 16298 -16388 16498 -16188
rect 9159 -16807 9359 -16607
rect 9417 -16807 9617 -16607
rect 9675 -16807 9875 -16607
rect 9933 -16807 10133 -16607
rect 10191 -16807 10391 -16607
rect 10449 -16807 10649 -16607
rect 10707 -16807 10907 -16607
rect 10965 -16807 11165 -16607
rect 11829 -16807 12029 -16607
rect 12087 -16807 12287 -16607
rect 12345 -16807 12545 -16607
rect 12603 -16807 12803 -16607
rect 12861 -16807 13061 -16607
rect 13119 -16807 13319 -16607
rect 13377 -16807 13577 -16607
rect 13635 -16807 13835 -16607
rect 14492 -16806 14692 -16606
rect 14750 -16806 14950 -16606
rect 15008 -16806 15208 -16606
rect 15266 -16806 15466 -16606
rect 15524 -16806 15724 -16606
rect 15782 -16806 15982 -16606
rect 16040 -16806 16240 -16606
rect 16298 -16806 16498 -16606
rect 9159 -17225 9359 -17025
rect 9417 -17225 9617 -17025
rect 9675 -17225 9875 -17025
rect 9933 -17225 10133 -17025
rect 10191 -17225 10391 -17025
rect 10449 -17225 10649 -17025
rect 10707 -17225 10907 -17025
rect 10965 -17225 11165 -17025
rect 11829 -17225 12029 -17025
rect 12087 -17225 12287 -17025
rect 12345 -17225 12545 -17025
rect 12603 -17225 12803 -17025
rect 12861 -17225 13061 -17025
rect 13119 -17225 13319 -17025
rect 13377 -17225 13577 -17025
rect 13635 -17225 13835 -17025
rect 14492 -17224 14692 -17024
rect 14750 -17224 14950 -17024
rect 15008 -17224 15208 -17024
rect 15266 -17224 15466 -17024
rect 15524 -17224 15724 -17024
rect 15782 -17224 15982 -17024
rect 16040 -17224 16240 -17024
rect 16298 -17224 16498 -17024
rect 9159 -17643 9359 -17443
rect 9417 -17643 9617 -17443
rect 9675 -17643 9875 -17443
rect 9933 -17643 10133 -17443
rect 10191 -17643 10391 -17443
rect 10449 -17643 10649 -17443
rect 10707 -17643 10907 -17443
rect 10965 -17643 11165 -17443
rect 11829 -17643 12029 -17443
rect 12087 -17643 12287 -17443
rect 12345 -17643 12545 -17443
rect 12603 -17643 12803 -17443
rect 12861 -17643 13061 -17443
rect 13119 -17643 13319 -17443
rect 13377 -17643 13577 -17443
rect 13635 -17643 13835 -17443
rect 14492 -17642 14692 -17442
rect 14750 -17642 14950 -17442
rect 15008 -17642 15208 -17442
rect 15266 -17642 15466 -17442
rect 15524 -17642 15724 -17442
rect 15782 -17642 15982 -17442
rect 16040 -17642 16240 -17442
rect 16298 -17642 16498 -17442
rect 9159 -18061 9359 -17861
rect 9417 -18061 9617 -17861
rect 9675 -18061 9875 -17861
rect 9933 -18061 10133 -17861
rect 10191 -18061 10391 -17861
rect 10449 -18061 10649 -17861
rect 10707 -18061 10907 -17861
rect 10965 -18061 11165 -17861
rect 11829 -18061 12029 -17861
rect 12087 -18061 12287 -17861
rect 12345 -18061 12545 -17861
rect 12603 -18061 12803 -17861
rect 12861 -18061 13061 -17861
rect 13119 -18061 13319 -17861
rect 13377 -18061 13577 -17861
rect 13635 -18061 13835 -17861
rect 14492 -18060 14692 -17860
rect 14750 -18060 14950 -17860
rect 15008 -18060 15208 -17860
rect 15266 -18060 15466 -17860
rect 15524 -18060 15724 -17860
rect 15782 -18060 15982 -17860
rect 16040 -18060 16240 -17860
rect 16298 -18060 16498 -17860
rect 9039 -18713 9239 -18513
rect 9579 -18713 9779 -18513
rect 10059 -18713 10259 -18513
rect 10562 -18711 10762 -18511
rect 11072 -18701 11272 -18501
rect 11709 -18713 11909 -18513
rect 12249 -18713 12449 -18513
rect 12729 -18713 12929 -18513
rect 13232 -18711 13432 -18511
rect 13742 -18701 13942 -18501
rect 14372 -18712 14572 -18512
rect 14912 -18712 15112 -18512
rect 15392 -18712 15592 -18512
rect 15895 -18710 16095 -18510
rect 16405 -18700 16605 -18500
rect 9159 -21457 9359 -21257
rect 9417 -21457 9617 -21257
rect 9675 -21457 9875 -21257
rect 9933 -21457 10133 -21257
rect 10191 -21457 10391 -21257
rect 10449 -21457 10649 -21257
rect 10707 -21457 10907 -21257
rect 10965 -21457 11165 -21257
rect 11829 -21457 12029 -21257
rect 12087 -21457 12287 -21257
rect 12345 -21457 12545 -21257
rect 12603 -21457 12803 -21257
rect 12861 -21457 13061 -21257
rect 13119 -21457 13319 -21257
rect 13377 -21457 13577 -21257
rect 13635 -21457 13835 -21257
rect 14492 -21456 14692 -21256
rect 14750 -21456 14950 -21256
rect 15008 -21456 15208 -21256
rect 15266 -21456 15466 -21256
rect 15524 -21456 15724 -21256
rect 15782 -21456 15982 -21256
rect 16040 -21456 16240 -21256
rect 16298 -21456 16498 -21256
rect 9159 -21875 9359 -21675
rect 9417 -21875 9617 -21675
rect 9675 -21875 9875 -21675
rect 9933 -21875 10133 -21675
rect 10191 -21875 10391 -21675
rect 10449 -21875 10649 -21675
rect 10707 -21875 10907 -21675
rect 10965 -21875 11165 -21675
rect 11829 -21875 12029 -21675
rect 12087 -21875 12287 -21675
rect 12345 -21875 12545 -21675
rect 12603 -21875 12803 -21675
rect 12861 -21875 13061 -21675
rect 13119 -21875 13319 -21675
rect 13377 -21875 13577 -21675
rect 13635 -21875 13835 -21675
rect 14492 -21874 14692 -21674
rect 14750 -21874 14950 -21674
rect 15008 -21874 15208 -21674
rect 15266 -21874 15466 -21674
rect 15524 -21874 15724 -21674
rect 15782 -21874 15982 -21674
rect 16040 -21874 16240 -21674
rect 16298 -21874 16498 -21674
rect 9159 -22293 9359 -22093
rect 9417 -22293 9617 -22093
rect 9675 -22293 9875 -22093
rect 9933 -22293 10133 -22093
rect 10191 -22293 10391 -22093
rect 10449 -22293 10649 -22093
rect 10707 -22293 10907 -22093
rect 10965 -22293 11165 -22093
rect 11829 -22293 12029 -22093
rect 12087 -22293 12287 -22093
rect 12345 -22293 12545 -22093
rect 12603 -22293 12803 -22093
rect 12861 -22293 13061 -22093
rect 13119 -22293 13319 -22093
rect 13377 -22293 13577 -22093
rect 13635 -22293 13835 -22093
rect 14492 -22292 14692 -22092
rect 14750 -22292 14950 -22092
rect 15008 -22292 15208 -22092
rect 15266 -22292 15466 -22092
rect 15524 -22292 15724 -22092
rect 15782 -22292 15982 -22092
rect 16040 -22292 16240 -22092
rect 16298 -22292 16498 -22092
rect 9159 -22711 9359 -22511
rect 9417 -22711 9617 -22511
rect 9675 -22711 9875 -22511
rect 9933 -22711 10133 -22511
rect 10191 -22711 10391 -22511
rect 10449 -22711 10649 -22511
rect 10707 -22711 10907 -22511
rect 10965 -22711 11165 -22511
rect 11829 -22711 12029 -22511
rect 12087 -22711 12287 -22511
rect 12345 -22711 12545 -22511
rect 12603 -22711 12803 -22511
rect 12861 -22711 13061 -22511
rect 13119 -22711 13319 -22511
rect 13377 -22711 13577 -22511
rect 13635 -22711 13835 -22511
rect 14492 -22710 14692 -22510
rect 14750 -22710 14950 -22510
rect 15008 -22710 15208 -22510
rect 15266 -22710 15466 -22510
rect 15524 -22710 15724 -22510
rect 15782 -22710 15982 -22510
rect 16040 -22710 16240 -22510
rect 16298 -22710 16498 -22510
rect 9159 -23129 9359 -22929
rect 9417 -23129 9617 -22929
rect 9675 -23129 9875 -22929
rect 9933 -23129 10133 -22929
rect 10191 -23129 10391 -22929
rect 10449 -23129 10649 -22929
rect 10707 -23129 10907 -22929
rect 10965 -23129 11165 -22929
rect 11829 -23129 12029 -22929
rect 12087 -23129 12287 -22929
rect 12345 -23129 12545 -22929
rect 12603 -23129 12803 -22929
rect 12861 -23129 13061 -22929
rect 13119 -23129 13319 -22929
rect 13377 -23129 13577 -22929
rect 13635 -23129 13835 -22929
rect 14492 -23128 14692 -22928
rect 14750 -23128 14950 -22928
rect 15008 -23128 15208 -22928
rect 15266 -23128 15466 -22928
rect 15524 -23128 15724 -22928
rect 15782 -23128 15982 -22928
rect 16040 -23128 16240 -22928
rect 16298 -23128 16498 -22928
rect 9159 -23547 9359 -23347
rect 9417 -23547 9617 -23347
rect 9675 -23547 9875 -23347
rect 9933 -23547 10133 -23347
rect 10191 -23547 10391 -23347
rect 10449 -23547 10649 -23347
rect 10707 -23547 10907 -23347
rect 10965 -23547 11165 -23347
rect 11829 -23547 12029 -23347
rect 12087 -23547 12287 -23347
rect 12345 -23547 12545 -23347
rect 12603 -23547 12803 -23347
rect 12861 -23547 13061 -23347
rect 13119 -23547 13319 -23347
rect 13377 -23547 13577 -23347
rect 13635 -23547 13835 -23347
rect 14492 -23546 14692 -23346
rect 14750 -23546 14950 -23346
rect 15008 -23546 15208 -23346
rect 15266 -23546 15466 -23346
rect 15524 -23546 15724 -23346
rect 15782 -23546 15982 -23346
rect 16040 -23546 16240 -23346
rect 16298 -23546 16498 -23346
rect 9159 -23965 9359 -23765
rect 9417 -23965 9617 -23765
rect 9675 -23965 9875 -23765
rect 9933 -23965 10133 -23765
rect 10191 -23965 10391 -23765
rect 10449 -23965 10649 -23765
rect 10707 -23965 10907 -23765
rect 10965 -23965 11165 -23765
rect 11829 -23965 12029 -23765
rect 12087 -23965 12287 -23765
rect 12345 -23965 12545 -23765
rect 12603 -23965 12803 -23765
rect 12861 -23965 13061 -23765
rect 13119 -23965 13319 -23765
rect 13377 -23965 13577 -23765
rect 13635 -23965 13835 -23765
rect 14492 -23964 14692 -23764
rect 14750 -23964 14950 -23764
rect 15008 -23964 15208 -23764
rect 15266 -23964 15466 -23764
rect 15524 -23964 15724 -23764
rect 15782 -23964 15982 -23764
rect 16040 -23964 16240 -23764
rect 16298 -23964 16498 -23764
rect 9039 -24617 9239 -24417
rect 9579 -24617 9779 -24417
rect 10059 -24617 10259 -24417
rect 10562 -24615 10762 -24415
rect 11072 -24605 11272 -24405
rect 11709 -24617 11909 -24417
rect 12249 -24617 12449 -24417
rect 12729 -24617 12929 -24417
rect 13232 -24615 13432 -24415
rect 13742 -24605 13942 -24405
rect 14372 -24616 14572 -24416
rect 14912 -24616 15112 -24416
rect 15392 -24616 15592 -24416
rect 15895 -24614 16095 -24414
rect 16405 -24604 16605 -24404
<< ndiff >>
rect 1086 4344 1144 4400
rect 1086 4256 1098 4344
rect 1132 4256 1144 4344
rect 1086 4200 1144 4256
rect 1174 4344 1232 4400
rect 1174 4256 1186 4344
rect 1220 4256 1232 4344
rect 1174 4200 1232 4256
rect 1302 4346 1360 4402
rect 1302 4258 1314 4346
rect 1348 4258 1360 4346
rect 1302 4202 1360 4258
rect 1390 4346 1448 4402
rect 1390 4258 1402 4346
rect 1436 4258 1448 4346
rect 1390 4202 1448 4258
rect 1520 4346 1578 4402
rect 1520 4258 1532 4346
rect 1566 4258 1578 4346
rect 1520 4202 1578 4258
rect 1608 4346 1666 4402
rect 1608 4258 1620 4346
rect 1654 4258 1666 4346
rect 1608 4202 1666 4258
rect 1742 4344 1800 4400
rect 1742 4256 1754 4344
rect 1788 4256 1800 4344
rect 1742 4200 1800 4256
rect 1830 4344 1888 4400
rect 1830 4256 1842 4344
rect 1876 4256 1888 4344
rect 1830 4200 1888 4256
rect 6272 4362 6330 4418
rect 6272 4274 6284 4362
rect 6318 4274 6330 4362
rect 6272 4218 6330 4274
rect 6360 4362 6418 4418
rect 6360 4274 6372 4362
rect 6406 4274 6418 4362
rect 6360 4218 6418 4274
rect 6488 4364 6546 4420
rect 6488 4276 6500 4364
rect 6534 4276 6546 4364
rect 6488 4220 6546 4276
rect 6576 4364 6634 4420
rect 6576 4276 6588 4364
rect 6622 4276 6634 4364
rect 6576 4220 6634 4276
rect 6706 4364 6764 4420
rect 6706 4276 6718 4364
rect 6752 4276 6764 4364
rect 6706 4220 6764 4276
rect 6794 4364 6852 4420
rect 6794 4276 6806 4364
rect 6840 4276 6852 4364
rect 6794 4220 6852 4276
rect 6928 4362 6986 4418
rect 6928 4274 6940 4362
rect 6974 4274 6986 4362
rect 6928 4218 6986 4274
rect 7016 4362 7074 4418
rect 7016 4274 7028 4362
rect 7062 4274 7074 4362
rect 7016 4218 7074 4274
rect 11448 4374 11506 4430
rect 11448 4286 11460 4374
rect 11494 4286 11506 4374
rect 11448 4230 11506 4286
rect 11536 4374 11594 4430
rect 11536 4286 11548 4374
rect 11582 4286 11594 4374
rect 11536 4230 11594 4286
rect 11664 4376 11722 4432
rect 11664 4288 11676 4376
rect 11710 4288 11722 4376
rect 11664 4232 11722 4288
rect 11752 4376 11810 4432
rect 11752 4288 11764 4376
rect 11798 4288 11810 4376
rect 11752 4232 11810 4288
rect 11882 4376 11940 4432
rect 11882 4288 11894 4376
rect 11928 4288 11940 4376
rect 11882 4232 11940 4288
rect 11970 4376 12028 4432
rect 11970 4288 11982 4376
rect 12016 4288 12028 4376
rect 11970 4232 12028 4288
rect 12104 4374 12162 4430
rect 12104 4286 12116 4374
rect 12150 4286 12162 4374
rect 12104 4230 12162 4286
rect 12192 4374 12250 4430
rect 12192 4286 12204 4374
rect 12238 4286 12250 4374
rect 12192 4230 12250 4286
rect 17104 4166 17162 4222
rect 17104 4078 17116 4166
rect 17150 4078 17162 4166
rect 17104 4022 17162 4078
rect 17192 4166 17250 4222
rect 17192 4078 17204 4166
rect 17238 4078 17250 4166
rect 17192 4022 17250 4078
rect 17320 4168 17378 4224
rect 17320 4080 17332 4168
rect 17366 4080 17378 4168
rect 17320 4024 17378 4080
rect 17408 4168 17466 4224
rect 17408 4080 17420 4168
rect 17454 4080 17466 4168
rect 17408 4024 17466 4080
rect 17538 4168 17596 4224
rect 17538 4080 17550 4168
rect 17584 4080 17596 4168
rect 17538 4024 17596 4080
rect 17626 4168 17684 4224
rect 17626 4080 17638 4168
rect 17672 4080 17684 4168
rect 17626 4024 17684 4080
rect 17760 4166 17818 4222
rect 17760 4078 17772 4166
rect 17806 4078 17818 4166
rect 17760 4022 17818 4078
rect 17848 4166 17906 4222
rect 17848 4078 17860 4166
rect 17894 4078 17906 4166
rect 17848 4022 17906 4078
rect 8774 3559 8832 3684
rect 8774 3409 8786 3559
rect 8820 3409 8832 3559
rect 8774 3284 8832 3409
rect 9032 3559 9090 3684
rect 9032 3409 9044 3559
rect 9078 3409 9090 3559
rect 9032 3284 9090 3409
rect 9290 3559 9348 3684
rect 9290 3409 9302 3559
rect 9336 3409 9348 3559
rect 9290 3284 9348 3409
rect 9548 3559 9606 3684
rect 9548 3409 9560 3559
rect 9594 3409 9606 3559
rect 9548 3284 9606 3409
rect 9788 3559 9846 3684
rect 9788 3409 9800 3559
rect 9834 3409 9846 3559
rect 9788 3284 9846 3409
rect 10046 3559 10104 3684
rect 10046 3409 10058 3559
rect 10092 3409 10104 3559
rect 10046 3284 10104 3409
rect 10304 3559 10362 3684
rect 10304 3409 10316 3559
rect 10350 3409 10362 3559
rect 10304 3284 10362 3409
rect 10562 3559 10620 3684
rect 10562 3409 10574 3559
rect 10608 3409 10620 3559
rect 10562 3284 10620 3409
rect -61826 3202 -61768 3246
rect -61830 3190 -61768 3202
rect -61830 3102 -61818 3190
rect -61784 3102 -61768 3190
rect -61830 3090 -61768 3102
rect -61826 3046 -61768 3090
rect -61738 3190 -61672 3246
rect -61738 3102 -61722 3190
rect -61688 3102 -61672 3190
rect -61738 3046 -61672 3102
rect -61642 3190 -61576 3246
rect -61642 3102 -61626 3190
rect -61592 3102 -61576 3190
rect -61642 3046 -61576 3102
rect -61546 3190 -61480 3246
rect -61546 3102 -61530 3190
rect -61496 3102 -61480 3190
rect -61546 3046 -61480 3102
rect -61450 3202 -61392 3246
rect -61450 3190 -61388 3202
rect -61450 3102 -61434 3190
rect -61400 3102 -61388 3190
rect -61450 3090 -61388 3102
rect -61450 3046 -61392 3090
rect 8774 3003 8832 3128
rect 8774 2853 8786 3003
rect 8820 2853 8832 3003
rect 8774 2728 8832 2853
rect 9032 3003 9090 3128
rect 9032 2853 9044 3003
rect 9078 2853 9090 3003
rect 9032 2728 9090 2853
rect 9290 3003 9348 3128
rect 9290 2853 9302 3003
rect 9336 2853 9348 3003
rect 9290 2728 9348 2853
rect 9548 3003 9606 3128
rect 9548 2853 9560 3003
rect 9594 2853 9606 3003
rect 9548 2728 9606 2853
rect 9788 3003 9846 3128
rect 9788 2853 9800 3003
rect 9834 2853 9846 3003
rect 9788 2728 9846 2853
rect 10046 3003 10104 3128
rect 10046 2853 10058 3003
rect 10092 2853 10104 3003
rect 10046 2728 10104 2853
rect 10304 3003 10362 3128
rect 10304 2853 10316 3003
rect 10350 2853 10362 3003
rect 10304 2728 10362 2853
rect 10562 3003 10620 3128
rect 10562 2853 10574 3003
rect 10608 2853 10620 3003
rect 10562 2728 10620 2853
rect 2614 2476 2672 2532
rect 2614 2388 2626 2476
rect 2660 2388 2672 2476
rect 2614 2332 2672 2388
rect 2872 2476 2930 2532
rect 2872 2388 2884 2476
rect 2918 2388 2930 2476
rect 2872 2332 2930 2388
rect 3090 2478 3148 2534
rect 3090 2390 3102 2478
rect 3136 2390 3148 2478
rect 3090 2334 3148 2390
rect 3948 2478 4006 2534
rect 3948 2390 3960 2478
rect 3994 2390 4006 2478
rect 3948 2334 4006 2390
rect 4062 2478 4120 2534
rect 4062 2390 4074 2478
rect 4108 2390 4120 2478
rect 4062 2334 4120 2390
rect 4920 2478 4978 2534
rect 4920 2390 4932 2478
rect 4966 2390 4978 2478
rect 4920 2334 4978 2390
rect 5148 2476 5206 2532
rect 5148 2388 5160 2476
rect 5194 2388 5206 2476
rect 5148 2332 5206 2388
rect 5406 2476 5464 2532
rect 5406 2388 5418 2476
rect 5452 2388 5464 2476
rect 5406 2332 5464 2388
rect 13306 2408 13364 3114
rect 9095 1828 9153 1884
rect 9095 1740 9107 1828
rect 9141 1740 9153 1828
rect 9095 1684 9153 1740
rect 9553 1828 9611 1884
rect 9553 1740 9565 1828
rect 9599 1740 9611 1828
rect 9553 1684 9611 1740
rect 9690 1828 9748 1884
rect 9690 1740 9702 1828
rect 9736 1740 9748 1828
rect 9690 1684 9748 1740
rect 10148 1828 10206 1884
rect 10148 1740 10160 1828
rect 10194 1740 10206 1828
rect 10148 1684 10206 1740
rect 13306 1020 13318 2408
rect 13352 1020 13364 2408
rect 13306 314 13364 1020
rect 13564 2408 13622 3114
rect 13564 1020 13576 2408
rect 13610 1020 13622 2408
rect 13856 2774 13914 2980
rect 13856 2386 13868 2774
rect 13902 2386 13914 2774
rect 13856 2180 13914 2386
rect 14114 2774 14172 2980
rect 14114 2386 14126 2774
rect 14160 2386 14172 2774
rect 14114 2180 14172 2386
rect 14372 2774 14430 2980
rect 14372 2386 14384 2774
rect 14418 2386 14430 2774
rect 14372 2180 14430 2386
rect 14630 2774 14688 2980
rect 14630 2386 14642 2774
rect 14676 2386 14688 2774
rect 14630 2180 14688 2386
rect 14856 2774 14914 2980
rect 14856 2386 14868 2774
rect 14902 2386 14914 2774
rect 14856 2180 14914 2386
rect 15114 2774 15172 2980
rect 15114 2386 15126 2774
rect 15160 2386 15172 2774
rect 15114 2180 15172 2386
rect 15372 2774 15430 2980
rect 15372 2386 15384 2774
rect 15418 2386 15430 2774
rect 15372 2180 15430 2386
rect 15630 2774 15688 2980
rect 15630 2386 15642 2774
rect 15676 2386 15688 2774
rect 15630 2180 15688 2386
rect 15904 2358 15962 3064
rect 13856 1818 13914 2024
rect 13856 1430 13868 1818
rect 13902 1430 13914 1818
rect 13856 1224 13914 1430
rect 14114 1818 14172 2024
rect 14114 1430 14126 1818
rect 14160 1430 14172 1818
rect 14114 1224 14172 1430
rect 14372 1818 14430 2024
rect 14372 1430 14384 1818
rect 14418 1430 14430 1818
rect 14372 1224 14430 1430
rect 14630 1818 14688 2024
rect 14630 1430 14642 1818
rect 14676 1430 14688 1818
rect 14630 1224 14688 1430
rect 14856 1818 14914 2024
rect 14856 1430 14868 1818
rect 14902 1430 14914 1818
rect 14856 1224 14914 1430
rect 15114 1818 15172 2024
rect 15114 1430 15126 1818
rect 15160 1430 15172 1818
rect 15114 1224 15172 1430
rect 15372 1818 15430 2024
rect 15372 1430 15384 1818
rect 15418 1430 15430 1818
rect 15372 1224 15430 1430
rect 15630 1818 15688 2024
rect 15630 1430 15642 1818
rect 15676 1430 15688 1818
rect 15630 1224 15688 1430
rect 13564 314 13622 1020
rect 13856 862 13914 1068
rect 13856 474 13868 862
rect 13902 474 13914 862
rect 13856 268 13914 474
rect 14114 862 14172 1068
rect 14114 474 14126 862
rect 14160 474 14172 862
rect 14114 268 14172 474
rect 14372 862 14430 1068
rect 14372 474 14384 862
rect 14418 474 14430 862
rect 14372 268 14430 474
rect 14630 862 14688 1068
rect 14630 474 14642 862
rect 14676 474 14688 862
rect 14630 268 14688 474
rect 14856 862 14914 1068
rect 14856 474 14868 862
rect 14902 474 14914 862
rect 14856 268 14914 474
rect 15114 862 15172 1068
rect 15114 474 15126 862
rect 15160 474 15172 862
rect 15114 268 15172 474
rect 15372 862 15430 1068
rect 15372 474 15384 862
rect 15418 474 15430 862
rect 15372 268 15430 474
rect 15630 862 15688 1068
rect 15630 474 15642 862
rect 15676 474 15688 862
rect 15630 268 15688 474
rect 15904 970 15916 2358
rect 15950 970 15962 2358
rect 15904 264 15962 970
rect 16162 2358 16220 3064
rect 16162 970 16174 2358
rect 16208 970 16220 2358
rect 26874 2196 26936 2208
rect 26874 2072 26886 2196
rect 26920 2072 26936 2196
rect 26874 2060 26936 2072
rect 26966 2196 27032 2208
rect 26966 2072 26982 2196
rect 27016 2072 27032 2196
rect 26966 2060 27032 2072
rect 27062 2196 27124 2208
rect 27062 2072 27078 2196
rect 27112 2072 27124 2196
rect 27062 2060 27124 2072
rect 27486 2204 27548 2216
rect 27486 2080 27498 2204
rect 27532 2080 27548 2204
rect 27486 2068 27548 2080
rect 27578 2204 27644 2216
rect 27578 2080 27594 2204
rect 27628 2080 27644 2204
rect 27578 2068 27644 2080
rect 27674 2204 27736 2216
rect 27674 2080 27690 2204
rect 27724 2080 27736 2204
rect 27674 2068 27736 2080
rect 28064 2200 28126 2212
rect 28064 2076 28076 2200
rect 28110 2076 28126 2200
rect 28064 2064 28126 2076
rect 28156 2200 28222 2212
rect 28156 2076 28172 2200
rect 28206 2076 28222 2200
rect 28156 2064 28222 2076
rect 28252 2200 28314 2212
rect 28252 2076 28268 2200
rect 28302 2076 28314 2200
rect 28252 2064 28314 2076
rect 28638 2208 28700 2220
rect 28638 2084 28650 2208
rect 28684 2084 28700 2208
rect 28638 2072 28700 2084
rect 28730 2208 28796 2220
rect 28730 2084 28746 2208
rect 28780 2084 28796 2208
rect 28730 2072 28796 2084
rect 28826 2208 28888 2220
rect 28826 2084 28842 2208
rect 28876 2084 28888 2208
rect 28826 2072 28888 2084
rect 29216 2208 29278 2220
rect 29216 2084 29228 2208
rect 29262 2084 29278 2208
rect 29216 2072 29278 2084
rect 29308 2208 29374 2220
rect 29308 2084 29324 2208
rect 29358 2084 29374 2208
rect 29308 2072 29374 2084
rect 29404 2208 29466 2220
rect 29404 2084 29420 2208
rect 29454 2084 29466 2208
rect 29404 2072 29466 2084
rect 29794 2208 29856 2220
rect 29794 2084 29806 2208
rect 29840 2084 29856 2208
rect 29794 2072 29856 2084
rect 29886 2208 29952 2220
rect 29886 2084 29902 2208
rect 29936 2084 29952 2208
rect 29886 2072 29952 2084
rect 29982 2208 30044 2220
rect 29982 2084 29998 2208
rect 30032 2084 30044 2208
rect 29982 2072 30044 2084
rect 30376 2212 30438 2224
rect 30376 2088 30388 2212
rect 30422 2088 30438 2212
rect 30376 2076 30438 2088
rect 30468 2212 30534 2224
rect 30468 2088 30484 2212
rect 30518 2088 30534 2212
rect 30468 2076 30534 2088
rect 30564 2212 30626 2224
rect 30564 2088 30580 2212
rect 30614 2088 30626 2212
rect 30564 2076 30626 2088
rect 30952 2208 31014 2220
rect 30952 2084 30964 2208
rect 30998 2084 31014 2208
rect 30952 2072 31014 2084
rect 31044 2208 31110 2220
rect 31044 2084 31060 2208
rect 31094 2084 31110 2208
rect 31044 2072 31110 2084
rect 31140 2208 31202 2220
rect 31140 2084 31156 2208
rect 31190 2084 31202 2208
rect 31140 2072 31202 2084
rect 31522 2204 31584 2216
rect 31522 2080 31534 2204
rect 31568 2080 31584 2204
rect 31522 2068 31584 2080
rect 31614 2204 31680 2216
rect 31614 2080 31630 2204
rect 31664 2080 31680 2204
rect 31614 2068 31680 2080
rect 31710 2204 31772 2216
rect 31710 2080 31726 2204
rect 31760 2080 31772 2204
rect 31710 2068 31772 2080
rect 16162 264 16220 970
rect 28932 358 28994 370
rect 28932 -266 28944 358
rect 28978 -266 28994 358
rect 28932 -278 28994 -266
rect 29024 358 29090 370
rect 29024 -266 29040 358
rect 29074 -266 29090 358
rect 29024 -278 29090 -266
rect 29120 358 29186 370
rect 29120 -266 29136 358
rect 29170 -266 29186 358
rect 29120 -278 29186 -266
rect 29216 358 29282 370
rect 29216 -266 29232 358
rect 29266 -266 29282 358
rect 29216 -278 29282 -266
rect 29312 358 29378 370
rect 29312 -266 29328 358
rect 29362 -266 29378 358
rect 29312 -278 29378 -266
rect 29408 358 29474 370
rect 29408 -266 29424 358
rect 29458 -266 29474 358
rect 29408 -278 29474 -266
rect 29504 358 29570 370
rect 29504 -266 29520 358
rect 29554 -266 29570 358
rect 29504 -278 29570 -266
rect 29600 358 29666 370
rect 29600 -266 29616 358
rect 29650 -266 29666 358
rect 29600 -278 29666 -266
rect 29696 358 29762 370
rect 29696 -266 29712 358
rect 29746 -266 29762 358
rect 29696 -278 29762 -266
rect 29792 358 29854 370
rect 29792 -266 29808 358
rect 29842 -266 29854 358
rect 29792 -278 29854 -266
rect 8761 -1400 8813 -1388
rect 8761 -1434 8769 -1400
rect 8803 -1434 8813 -1400
rect 8761 -1472 8813 -1434
rect 8843 -1426 8897 -1388
rect 8843 -1460 8853 -1426
rect 8887 -1460 8897 -1426
rect 8843 -1472 8897 -1460
rect 8927 -1400 8979 -1388
rect 8927 -1434 8937 -1400
rect 8971 -1434 8979 -1400
rect 8927 -1472 8979 -1434
rect 9047 -1430 9152 -1388
rect 9047 -1464 9059 -1430
rect 9093 -1464 9152 -1430
rect 9047 -1472 9152 -1464
rect 9182 -1400 9232 -1388
rect 9663 -1388 9713 -1344
rect 9391 -1400 9509 -1388
rect 9182 -1424 9247 -1400
rect 9182 -1458 9192 -1424
rect 9226 -1458 9247 -1424
rect 9182 -1472 9247 -1458
rect 9277 -1424 9343 -1400
rect 9277 -1458 9299 -1424
rect 9333 -1458 9343 -1424
rect 9277 -1472 9343 -1458
rect 9373 -1472 9509 -1400
rect 9539 -1472 9581 -1388
rect 9611 -1426 9713 -1388
rect 9611 -1460 9645 -1426
rect 9679 -1460 9713 -1426
rect 9611 -1472 9713 -1460
rect 9743 -1400 9797 -1344
rect 10393 -1387 10445 -1342
rect 9967 -1400 10017 -1388
rect 9743 -1430 9812 -1400
rect 9743 -1464 9757 -1430
rect 9791 -1464 9812 -1430
rect 9743 -1472 9812 -1464
rect 9842 -1426 9921 -1400
rect 9842 -1460 9867 -1426
rect 9901 -1460 9921 -1426
rect 9842 -1472 9921 -1460
rect 9951 -1472 10017 -1400
rect 10047 -1430 10166 -1388
rect 10047 -1464 10079 -1430
rect 10113 -1464 10166 -1430
rect 10047 -1472 10166 -1464
rect 10196 -1472 10257 -1388
rect 10287 -1410 10339 -1388
rect 10287 -1444 10297 -1410
rect 10331 -1444 10339 -1410
rect 10287 -1472 10339 -1444
rect 10393 -1421 10401 -1387
rect 10435 -1421 10445 -1387
rect 10393 -1472 10445 -1421
rect 10475 -1354 10527 -1342
rect 10475 -1388 10485 -1354
rect 10519 -1388 10527 -1354
rect 10678 -1388 10730 -1342
rect 10475 -1422 10527 -1388
rect 10475 -1456 10485 -1422
rect 10519 -1456 10527 -1422
rect 10475 -1472 10527 -1456
rect 10581 -1400 10633 -1388
rect 10581 -1434 10589 -1400
rect 10623 -1434 10633 -1400
rect 10581 -1472 10633 -1434
rect 10663 -1406 10730 -1388
rect 10663 -1440 10686 -1406
rect 10720 -1440 10730 -1406
rect 10663 -1472 10730 -1440
rect 10760 -1376 10812 -1342
rect 10760 -1410 10770 -1376
rect 10804 -1410 10812 -1376
rect 10760 -1472 10812 -1410
rect 11227 -1400 11279 -1388
rect 11227 -1434 11235 -1400
rect 11269 -1434 11279 -1400
rect 11227 -1472 11279 -1434
rect 11309 -1426 11363 -1388
rect 11309 -1460 11319 -1426
rect 11353 -1460 11363 -1426
rect 11309 -1472 11363 -1460
rect 11393 -1400 11445 -1388
rect 11393 -1434 11403 -1400
rect 11437 -1434 11445 -1400
rect 11393 -1472 11445 -1434
rect 11513 -1430 11618 -1388
rect 11513 -1464 11525 -1430
rect 11559 -1464 11618 -1430
rect 11513 -1472 11618 -1464
rect 11648 -1400 11698 -1388
rect 12129 -1388 12179 -1344
rect 11857 -1400 11975 -1388
rect 11648 -1424 11713 -1400
rect 11648 -1458 11658 -1424
rect 11692 -1458 11713 -1424
rect 11648 -1472 11713 -1458
rect 11743 -1424 11809 -1400
rect 11743 -1458 11765 -1424
rect 11799 -1458 11809 -1424
rect 11743 -1472 11809 -1458
rect 11839 -1472 11975 -1400
rect 12005 -1472 12047 -1388
rect 12077 -1426 12179 -1388
rect 12077 -1460 12111 -1426
rect 12145 -1460 12179 -1426
rect 12077 -1472 12179 -1460
rect 12209 -1400 12263 -1344
rect 12859 -1387 12911 -1342
rect 12433 -1400 12483 -1388
rect 12209 -1430 12278 -1400
rect 12209 -1464 12223 -1430
rect 12257 -1464 12278 -1430
rect 12209 -1472 12278 -1464
rect 12308 -1426 12387 -1400
rect 12308 -1460 12333 -1426
rect 12367 -1460 12387 -1426
rect 12308 -1472 12387 -1460
rect 12417 -1472 12483 -1400
rect 12513 -1430 12632 -1388
rect 12513 -1464 12545 -1430
rect 12579 -1464 12632 -1430
rect 12513 -1472 12632 -1464
rect 12662 -1472 12723 -1388
rect 12753 -1410 12805 -1388
rect 12753 -1444 12763 -1410
rect 12797 -1444 12805 -1410
rect 12753 -1472 12805 -1444
rect 12859 -1421 12867 -1387
rect 12901 -1421 12911 -1387
rect 12859 -1472 12911 -1421
rect 12941 -1354 12993 -1342
rect 12941 -1388 12951 -1354
rect 12985 -1388 12993 -1354
rect 13144 -1388 13196 -1342
rect 12941 -1422 12993 -1388
rect 12941 -1456 12951 -1422
rect 12985 -1456 12993 -1422
rect 12941 -1472 12993 -1456
rect 13047 -1400 13099 -1388
rect 13047 -1434 13055 -1400
rect 13089 -1434 13099 -1400
rect 13047 -1472 13099 -1434
rect 13129 -1406 13196 -1388
rect 13129 -1440 13152 -1406
rect 13186 -1440 13196 -1406
rect 13129 -1472 13196 -1440
rect 13226 -1376 13278 -1342
rect 13226 -1410 13236 -1376
rect 13270 -1410 13278 -1376
rect 13226 -1472 13278 -1410
rect 10181 -2156 10233 -2144
rect 10181 -2190 10189 -2156
rect 10223 -2190 10233 -2156
rect 10181 -2228 10233 -2190
rect 10181 -2262 10189 -2228
rect 10223 -2262 10233 -2228
rect 10181 -2274 10233 -2262
rect 10263 -2156 10317 -2144
rect 10263 -2190 10273 -2156
rect 10307 -2190 10317 -2156
rect 10263 -2228 10317 -2190
rect 10263 -2262 10273 -2228
rect 10307 -2262 10317 -2228
rect 10263 -2274 10317 -2262
rect 10347 -2156 10399 -2144
rect 10347 -2190 10357 -2156
rect 10391 -2190 10399 -2156
rect 10347 -2228 10399 -2190
rect 10347 -2262 10357 -2228
rect 10391 -2262 10399 -2228
rect 10347 -2274 10399 -2262
rect 11227 -2202 11279 -2190
rect 11227 -2236 11235 -2202
rect 11269 -2236 11279 -2202
rect 11227 -2274 11279 -2236
rect 11309 -2228 11363 -2190
rect 11309 -2262 11319 -2228
rect 11353 -2262 11363 -2228
rect 11309 -2274 11363 -2262
rect 11393 -2202 11445 -2190
rect 11393 -2236 11403 -2202
rect 11437 -2236 11445 -2202
rect 11393 -2274 11445 -2236
rect 11513 -2232 11618 -2190
rect 11513 -2266 11525 -2232
rect 11559 -2266 11618 -2232
rect 11513 -2274 11618 -2266
rect 11648 -2202 11698 -2190
rect 12129 -2190 12179 -2146
rect 11857 -2202 11975 -2190
rect 11648 -2226 11713 -2202
rect 11648 -2260 11658 -2226
rect 11692 -2260 11713 -2226
rect 11648 -2274 11713 -2260
rect 11743 -2226 11809 -2202
rect 11743 -2260 11765 -2226
rect 11799 -2260 11809 -2226
rect 11743 -2274 11809 -2260
rect 11839 -2274 11975 -2202
rect 12005 -2274 12047 -2190
rect 12077 -2228 12179 -2190
rect 12077 -2262 12111 -2228
rect 12145 -2262 12179 -2228
rect 12077 -2274 12179 -2262
rect 12209 -2202 12263 -2146
rect 12859 -2189 12911 -2144
rect 12433 -2202 12483 -2190
rect 12209 -2232 12278 -2202
rect 12209 -2266 12223 -2232
rect 12257 -2266 12278 -2232
rect 12209 -2274 12278 -2266
rect 12308 -2228 12387 -2202
rect 12308 -2262 12333 -2228
rect 12367 -2262 12387 -2228
rect 12308 -2274 12387 -2262
rect 12417 -2274 12483 -2202
rect 12513 -2232 12632 -2190
rect 12513 -2266 12545 -2232
rect 12579 -2266 12632 -2232
rect 12513 -2274 12632 -2266
rect 12662 -2274 12723 -2190
rect 12753 -2212 12805 -2190
rect 12753 -2246 12763 -2212
rect 12797 -2246 12805 -2212
rect 12753 -2274 12805 -2246
rect 12859 -2223 12867 -2189
rect 12901 -2223 12911 -2189
rect 12859 -2274 12911 -2223
rect 12941 -2156 12993 -2144
rect 12941 -2190 12951 -2156
rect 12985 -2190 12993 -2156
rect 13144 -2190 13196 -2144
rect 12941 -2224 12993 -2190
rect 12941 -2258 12951 -2224
rect 12985 -2258 12993 -2224
rect 12941 -2274 12993 -2258
rect 13047 -2202 13099 -2190
rect 13047 -2236 13055 -2202
rect 13089 -2236 13099 -2202
rect 13047 -2274 13099 -2236
rect 13129 -2208 13196 -2190
rect 13129 -2242 13152 -2208
rect 13186 -2242 13196 -2208
rect 13129 -2274 13196 -2242
rect 13226 -2178 13278 -2144
rect 13226 -2212 13236 -2178
rect 13270 -2212 13278 -2178
rect 13226 -2274 13278 -2212
rect -9131 -4670 -9079 -4658
rect -9131 -4704 -9123 -4670
rect -9089 -4704 -9079 -4670
rect -9131 -4742 -9079 -4704
rect -9049 -4696 -8995 -4658
rect -9049 -4730 -9039 -4696
rect -9005 -4730 -8995 -4696
rect -9049 -4742 -8995 -4730
rect -8965 -4670 -8913 -4658
rect -8965 -4704 -8955 -4670
rect -8921 -4704 -8913 -4670
rect -8965 -4742 -8913 -4704
rect -8845 -4700 -8740 -4658
rect -8845 -4734 -8833 -4700
rect -8799 -4734 -8740 -4700
rect -8845 -4742 -8740 -4734
rect -8710 -4670 -8660 -4658
rect -8229 -4658 -8179 -4614
rect -8501 -4670 -8383 -4658
rect -8710 -4694 -8645 -4670
rect -8710 -4728 -8700 -4694
rect -8666 -4728 -8645 -4694
rect -8710 -4742 -8645 -4728
rect -8615 -4694 -8549 -4670
rect -8615 -4728 -8593 -4694
rect -8559 -4728 -8549 -4694
rect -8615 -4742 -8549 -4728
rect -8519 -4742 -8383 -4670
rect -8353 -4742 -8311 -4658
rect -8281 -4696 -8179 -4658
rect -8281 -4730 -8247 -4696
rect -8213 -4730 -8179 -4696
rect -8281 -4742 -8179 -4730
rect -8149 -4670 -8095 -4614
rect -7499 -4657 -7447 -4612
rect -7925 -4670 -7875 -4658
rect -8149 -4700 -8080 -4670
rect -8149 -4734 -8135 -4700
rect -8101 -4734 -8080 -4700
rect -8149 -4742 -8080 -4734
rect -8050 -4696 -7971 -4670
rect -8050 -4730 -8025 -4696
rect -7991 -4730 -7971 -4696
rect -8050 -4742 -7971 -4730
rect -7941 -4742 -7875 -4670
rect -7845 -4700 -7726 -4658
rect -7845 -4734 -7813 -4700
rect -7779 -4734 -7726 -4700
rect -7845 -4742 -7726 -4734
rect -7696 -4742 -7635 -4658
rect -7605 -4680 -7553 -4658
rect -7605 -4714 -7595 -4680
rect -7561 -4714 -7553 -4680
rect -7605 -4742 -7553 -4714
rect -7499 -4691 -7491 -4657
rect -7457 -4691 -7447 -4657
rect -7499 -4742 -7447 -4691
rect -7417 -4624 -7365 -4612
rect -7417 -4658 -7407 -4624
rect -7373 -4658 -7365 -4624
rect -7214 -4658 -7162 -4612
rect -7417 -4692 -7365 -4658
rect -7417 -4726 -7407 -4692
rect -7373 -4726 -7365 -4692
rect -7417 -4742 -7365 -4726
rect -7311 -4670 -7259 -4658
rect -7311 -4704 -7303 -4670
rect -7269 -4704 -7259 -4670
rect -7311 -4742 -7259 -4704
rect -7229 -4676 -7162 -4658
rect -7229 -4710 -7206 -4676
rect -7172 -4710 -7162 -4676
rect -7229 -4742 -7162 -4710
rect -7132 -4646 -7080 -4612
rect -7132 -4680 -7122 -4646
rect -7088 -4680 -7080 -4646
rect -7132 -4742 -7080 -4680
rect -7015 -4670 -6963 -4658
rect -7015 -4704 -7007 -4670
rect -6973 -4704 -6963 -4670
rect -7015 -4742 -6963 -4704
rect -6933 -4696 -6879 -4658
rect -6933 -4730 -6923 -4696
rect -6889 -4730 -6879 -4696
rect -6933 -4742 -6879 -4730
rect -6849 -4670 -6797 -4658
rect -6849 -4704 -6839 -4670
rect -6805 -4704 -6797 -4670
rect -6849 -4742 -6797 -4704
rect -6729 -4700 -6624 -4658
rect -6729 -4734 -6717 -4700
rect -6683 -4734 -6624 -4700
rect -6729 -4742 -6624 -4734
rect -6594 -4670 -6544 -4658
rect -6113 -4658 -6063 -4614
rect -6385 -4670 -6267 -4658
rect -6594 -4694 -6529 -4670
rect -6594 -4728 -6584 -4694
rect -6550 -4728 -6529 -4694
rect -6594 -4742 -6529 -4728
rect -6499 -4694 -6433 -4670
rect -6499 -4728 -6477 -4694
rect -6443 -4728 -6433 -4694
rect -6499 -4742 -6433 -4728
rect -6403 -4742 -6267 -4670
rect -6237 -4742 -6195 -4658
rect -6165 -4696 -6063 -4658
rect -6165 -4730 -6131 -4696
rect -6097 -4730 -6063 -4696
rect -6165 -4742 -6063 -4730
rect -6033 -4670 -5979 -4614
rect -5383 -4657 -5331 -4612
rect -5809 -4670 -5759 -4658
rect -6033 -4700 -5964 -4670
rect -6033 -4734 -6019 -4700
rect -5985 -4734 -5964 -4700
rect -6033 -4742 -5964 -4734
rect -5934 -4696 -5855 -4670
rect -5934 -4730 -5909 -4696
rect -5875 -4730 -5855 -4696
rect -5934 -4742 -5855 -4730
rect -5825 -4742 -5759 -4670
rect -5729 -4700 -5610 -4658
rect -5729 -4734 -5697 -4700
rect -5663 -4734 -5610 -4700
rect -5729 -4742 -5610 -4734
rect -5580 -4742 -5519 -4658
rect -5489 -4680 -5437 -4658
rect -5489 -4714 -5479 -4680
rect -5445 -4714 -5437 -4680
rect -5489 -4742 -5437 -4714
rect -5383 -4691 -5375 -4657
rect -5341 -4691 -5331 -4657
rect -5383 -4742 -5331 -4691
rect -5301 -4624 -5249 -4612
rect -5301 -4658 -5291 -4624
rect -5257 -4658 -5249 -4624
rect -5098 -4658 -5046 -4612
rect -5301 -4692 -5249 -4658
rect -5301 -4726 -5291 -4692
rect -5257 -4726 -5249 -4692
rect -5301 -4742 -5249 -4726
rect -5195 -4670 -5143 -4658
rect -5195 -4704 -5187 -4670
rect -5153 -4704 -5143 -4670
rect -5195 -4742 -5143 -4704
rect -5113 -4676 -5046 -4658
rect -5113 -4710 -5090 -4676
rect -5056 -4710 -5046 -4676
rect -5113 -4742 -5046 -4710
rect -5016 -4646 -4964 -4612
rect -5016 -4680 -5006 -4646
rect -4972 -4680 -4964 -4646
rect -5016 -4742 -4964 -4680
rect -4899 -4670 -4847 -4658
rect -4899 -4704 -4891 -4670
rect -4857 -4704 -4847 -4670
rect -4899 -4742 -4847 -4704
rect -4817 -4696 -4763 -4658
rect -4817 -4730 -4807 -4696
rect -4773 -4730 -4763 -4696
rect -4817 -4742 -4763 -4730
rect -4733 -4670 -4681 -4658
rect -4733 -4704 -4723 -4670
rect -4689 -4704 -4681 -4670
rect -4733 -4742 -4681 -4704
rect -4613 -4700 -4508 -4658
rect -4613 -4734 -4601 -4700
rect -4567 -4734 -4508 -4700
rect -4613 -4742 -4508 -4734
rect -4478 -4670 -4428 -4658
rect -3997 -4658 -3947 -4614
rect -4269 -4670 -4151 -4658
rect -4478 -4694 -4413 -4670
rect -4478 -4728 -4468 -4694
rect -4434 -4728 -4413 -4694
rect -4478 -4742 -4413 -4728
rect -4383 -4694 -4317 -4670
rect -4383 -4728 -4361 -4694
rect -4327 -4728 -4317 -4694
rect -4383 -4742 -4317 -4728
rect -4287 -4742 -4151 -4670
rect -4121 -4742 -4079 -4658
rect -4049 -4696 -3947 -4658
rect -4049 -4730 -4015 -4696
rect -3981 -4730 -3947 -4696
rect -4049 -4742 -3947 -4730
rect -3917 -4670 -3863 -4614
rect -3267 -4657 -3215 -4612
rect -3693 -4670 -3643 -4658
rect -3917 -4700 -3848 -4670
rect -3917 -4734 -3903 -4700
rect -3869 -4734 -3848 -4700
rect -3917 -4742 -3848 -4734
rect -3818 -4696 -3739 -4670
rect -3818 -4730 -3793 -4696
rect -3759 -4730 -3739 -4696
rect -3818 -4742 -3739 -4730
rect -3709 -4742 -3643 -4670
rect -3613 -4700 -3494 -4658
rect -3613 -4734 -3581 -4700
rect -3547 -4734 -3494 -4700
rect -3613 -4742 -3494 -4734
rect -3464 -4742 -3403 -4658
rect -3373 -4680 -3321 -4658
rect -3373 -4714 -3363 -4680
rect -3329 -4714 -3321 -4680
rect -3373 -4742 -3321 -4714
rect -3267 -4691 -3259 -4657
rect -3225 -4691 -3215 -4657
rect -3267 -4742 -3215 -4691
rect -3185 -4624 -3133 -4612
rect -3185 -4658 -3175 -4624
rect -3141 -4658 -3133 -4624
rect -2982 -4658 -2930 -4612
rect -3185 -4692 -3133 -4658
rect -3185 -4726 -3175 -4692
rect -3141 -4726 -3133 -4692
rect -3185 -4742 -3133 -4726
rect -3079 -4670 -3027 -4658
rect -3079 -4704 -3071 -4670
rect -3037 -4704 -3027 -4670
rect -3079 -4742 -3027 -4704
rect -2997 -4676 -2930 -4658
rect -2997 -4710 -2974 -4676
rect -2940 -4710 -2930 -4676
rect -2997 -4742 -2930 -4710
rect -2900 -4646 -2848 -4612
rect -2900 -4680 -2890 -4646
rect -2856 -4680 -2848 -4646
rect -2900 -4742 -2848 -4680
rect -2783 -4670 -2731 -4658
rect -2783 -4704 -2775 -4670
rect -2741 -4704 -2731 -4670
rect -2783 -4742 -2731 -4704
rect -2701 -4696 -2647 -4658
rect -2701 -4730 -2691 -4696
rect -2657 -4730 -2647 -4696
rect -2701 -4742 -2647 -4730
rect -2617 -4670 -2565 -4658
rect -2617 -4704 -2607 -4670
rect -2573 -4704 -2565 -4670
rect -2617 -4742 -2565 -4704
rect -2497 -4700 -2392 -4658
rect -2497 -4734 -2485 -4700
rect -2451 -4734 -2392 -4700
rect -2497 -4742 -2392 -4734
rect -2362 -4670 -2312 -4658
rect -1881 -4658 -1831 -4614
rect -2153 -4670 -2035 -4658
rect -2362 -4694 -2297 -4670
rect -2362 -4728 -2352 -4694
rect -2318 -4728 -2297 -4694
rect -2362 -4742 -2297 -4728
rect -2267 -4694 -2201 -4670
rect -2267 -4728 -2245 -4694
rect -2211 -4728 -2201 -4694
rect -2267 -4742 -2201 -4728
rect -2171 -4742 -2035 -4670
rect -2005 -4742 -1963 -4658
rect -1933 -4696 -1831 -4658
rect -1933 -4730 -1899 -4696
rect -1865 -4730 -1831 -4696
rect -1933 -4742 -1831 -4730
rect -1801 -4670 -1747 -4614
rect -1151 -4657 -1099 -4612
rect -1577 -4670 -1527 -4658
rect -1801 -4700 -1732 -4670
rect -1801 -4734 -1787 -4700
rect -1753 -4734 -1732 -4700
rect -1801 -4742 -1732 -4734
rect -1702 -4696 -1623 -4670
rect -1702 -4730 -1677 -4696
rect -1643 -4730 -1623 -4696
rect -1702 -4742 -1623 -4730
rect -1593 -4742 -1527 -4670
rect -1497 -4700 -1378 -4658
rect -1497 -4734 -1465 -4700
rect -1431 -4734 -1378 -4700
rect -1497 -4742 -1378 -4734
rect -1348 -4742 -1287 -4658
rect -1257 -4680 -1205 -4658
rect -1257 -4714 -1247 -4680
rect -1213 -4714 -1205 -4680
rect -1257 -4742 -1205 -4714
rect -1151 -4691 -1143 -4657
rect -1109 -4691 -1099 -4657
rect -1151 -4742 -1099 -4691
rect -1069 -4624 -1017 -4612
rect -1069 -4658 -1059 -4624
rect -1025 -4658 -1017 -4624
rect -866 -4658 -814 -4612
rect -1069 -4692 -1017 -4658
rect -1069 -4726 -1059 -4692
rect -1025 -4726 -1017 -4692
rect -1069 -4742 -1017 -4726
rect -963 -4670 -911 -4658
rect -963 -4704 -955 -4670
rect -921 -4704 -911 -4670
rect -963 -4742 -911 -4704
rect -881 -4676 -814 -4658
rect -881 -4710 -858 -4676
rect -824 -4710 -814 -4676
rect -881 -4742 -814 -4710
rect -784 -4646 -732 -4612
rect -784 -4680 -774 -4646
rect -740 -4680 -732 -4646
rect -784 -4742 -732 -4680
rect -667 -4670 -615 -4658
rect -667 -4704 -659 -4670
rect -625 -4704 -615 -4670
rect -667 -4742 -615 -4704
rect -585 -4696 -531 -4658
rect -585 -4730 -575 -4696
rect -541 -4730 -531 -4696
rect -585 -4742 -531 -4730
rect -501 -4670 -449 -4658
rect -501 -4704 -491 -4670
rect -457 -4704 -449 -4670
rect -501 -4742 -449 -4704
rect -381 -4700 -276 -4658
rect -381 -4734 -369 -4700
rect -335 -4734 -276 -4700
rect -381 -4742 -276 -4734
rect -246 -4670 -196 -4658
rect 235 -4658 285 -4614
rect -37 -4670 81 -4658
rect -246 -4694 -181 -4670
rect -246 -4728 -236 -4694
rect -202 -4728 -181 -4694
rect -246 -4742 -181 -4728
rect -151 -4694 -85 -4670
rect -151 -4728 -129 -4694
rect -95 -4728 -85 -4694
rect -151 -4742 -85 -4728
rect -55 -4742 81 -4670
rect 111 -4742 153 -4658
rect 183 -4696 285 -4658
rect 183 -4730 217 -4696
rect 251 -4730 285 -4696
rect 183 -4742 285 -4730
rect 315 -4670 369 -4614
rect 965 -4657 1017 -4612
rect 539 -4670 589 -4658
rect 315 -4700 384 -4670
rect 315 -4734 329 -4700
rect 363 -4734 384 -4700
rect 315 -4742 384 -4734
rect 414 -4696 493 -4670
rect 414 -4730 439 -4696
rect 473 -4730 493 -4696
rect 414 -4742 493 -4730
rect 523 -4742 589 -4670
rect 619 -4700 738 -4658
rect 619 -4734 651 -4700
rect 685 -4734 738 -4700
rect 619 -4742 738 -4734
rect 768 -4742 829 -4658
rect 859 -4680 911 -4658
rect 859 -4714 869 -4680
rect 903 -4714 911 -4680
rect 859 -4742 911 -4714
rect 965 -4691 973 -4657
rect 1007 -4691 1017 -4657
rect 965 -4742 1017 -4691
rect 1047 -4624 1099 -4612
rect 1047 -4658 1057 -4624
rect 1091 -4658 1099 -4624
rect 1250 -4658 1302 -4612
rect 1047 -4692 1099 -4658
rect 1047 -4726 1057 -4692
rect 1091 -4726 1099 -4692
rect 1047 -4742 1099 -4726
rect 1153 -4670 1205 -4658
rect 1153 -4704 1161 -4670
rect 1195 -4704 1205 -4670
rect 1153 -4742 1205 -4704
rect 1235 -4676 1302 -4658
rect 1235 -4710 1258 -4676
rect 1292 -4710 1302 -4676
rect 1235 -4742 1302 -4710
rect 1332 -4646 1384 -4612
rect 1332 -4680 1342 -4646
rect 1376 -4680 1384 -4646
rect 1332 -4742 1384 -4680
rect 1449 -4670 1501 -4658
rect 1449 -4704 1457 -4670
rect 1491 -4704 1501 -4670
rect 1449 -4742 1501 -4704
rect 1531 -4696 1585 -4658
rect 1531 -4730 1541 -4696
rect 1575 -4730 1585 -4696
rect 1531 -4742 1585 -4730
rect 1615 -4670 1667 -4658
rect 1615 -4704 1625 -4670
rect 1659 -4704 1667 -4670
rect 1615 -4742 1667 -4704
rect 1735 -4700 1840 -4658
rect 1735 -4734 1747 -4700
rect 1781 -4734 1840 -4700
rect 1735 -4742 1840 -4734
rect 1870 -4670 1920 -4658
rect 2351 -4658 2401 -4614
rect 2079 -4670 2197 -4658
rect 1870 -4694 1935 -4670
rect 1870 -4728 1880 -4694
rect 1914 -4728 1935 -4694
rect 1870 -4742 1935 -4728
rect 1965 -4694 2031 -4670
rect 1965 -4728 1987 -4694
rect 2021 -4728 2031 -4694
rect 1965 -4742 2031 -4728
rect 2061 -4742 2197 -4670
rect 2227 -4742 2269 -4658
rect 2299 -4696 2401 -4658
rect 2299 -4730 2333 -4696
rect 2367 -4730 2401 -4696
rect 2299 -4742 2401 -4730
rect 2431 -4670 2485 -4614
rect 3081 -4657 3133 -4612
rect 2655 -4670 2705 -4658
rect 2431 -4700 2500 -4670
rect 2431 -4734 2445 -4700
rect 2479 -4734 2500 -4700
rect 2431 -4742 2500 -4734
rect 2530 -4696 2609 -4670
rect 2530 -4730 2555 -4696
rect 2589 -4730 2609 -4696
rect 2530 -4742 2609 -4730
rect 2639 -4742 2705 -4670
rect 2735 -4700 2854 -4658
rect 2735 -4734 2767 -4700
rect 2801 -4734 2854 -4700
rect 2735 -4742 2854 -4734
rect 2884 -4742 2945 -4658
rect 2975 -4680 3027 -4658
rect 2975 -4714 2985 -4680
rect 3019 -4714 3027 -4680
rect 2975 -4742 3027 -4714
rect 3081 -4691 3089 -4657
rect 3123 -4691 3133 -4657
rect 3081 -4742 3133 -4691
rect 3163 -4624 3215 -4612
rect 3163 -4658 3173 -4624
rect 3207 -4658 3215 -4624
rect 3366 -4658 3418 -4612
rect 3163 -4692 3215 -4658
rect 3163 -4726 3173 -4692
rect 3207 -4726 3215 -4692
rect 3163 -4742 3215 -4726
rect 3269 -4670 3321 -4658
rect 3269 -4704 3277 -4670
rect 3311 -4704 3321 -4670
rect 3269 -4742 3321 -4704
rect 3351 -4676 3418 -4658
rect 3351 -4710 3374 -4676
rect 3408 -4710 3418 -4676
rect 3351 -4742 3418 -4710
rect 3448 -4646 3500 -4612
rect 3448 -4680 3458 -4646
rect 3492 -4680 3500 -4646
rect 3448 -4742 3500 -4680
rect 3565 -4670 3617 -4658
rect 3565 -4704 3573 -4670
rect 3607 -4704 3617 -4670
rect 3565 -4742 3617 -4704
rect 3647 -4696 3701 -4658
rect 3647 -4730 3657 -4696
rect 3691 -4730 3701 -4696
rect 3647 -4742 3701 -4730
rect 3731 -4670 3783 -4658
rect 3731 -4704 3741 -4670
rect 3775 -4704 3783 -4670
rect 3731 -4742 3783 -4704
rect 3851 -4700 3956 -4658
rect 3851 -4734 3863 -4700
rect 3897 -4734 3956 -4700
rect 3851 -4742 3956 -4734
rect 3986 -4670 4036 -4658
rect 4467 -4658 4517 -4614
rect 4195 -4670 4313 -4658
rect 3986 -4694 4051 -4670
rect 3986 -4728 3996 -4694
rect 4030 -4728 4051 -4694
rect 3986 -4742 4051 -4728
rect 4081 -4694 4147 -4670
rect 4081 -4728 4103 -4694
rect 4137 -4728 4147 -4694
rect 4081 -4742 4147 -4728
rect 4177 -4742 4313 -4670
rect 4343 -4742 4385 -4658
rect 4415 -4696 4517 -4658
rect 4415 -4730 4449 -4696
rect 4483 -4730 4517 -4696
rect 4415 -4742 4517 -4730
rect 4547 -4670 4601 -4614
rect 5197 -4657 5249 -4612
rect 4771 -4670 4821 -4658
rect 4547 -4700 4616 -4670
rect 4547 -4734 4561 -4700
rect 4595 -4734 4616 -4700
rect 4547 -4742 4616 -4734
rect 4646 -4696 4725 -4670
rect 4646 -4730 4671 -4696
rect 4705 -4730 4725 -4696
rect 4646 -4742 4725 -4730
rect 4755 -4742 4821 -4670
rect 4851 -4700 4970 -4658
rect 4851 -4734 4883 -4700
rect 4917 -4734 4970 -4700
rect 4851 -4742 4970 -4734
rect 5000 -4742 5061 -4658
rect 5091 -4680 5143 -4658
rect 5091 -4714 5101 -4680
rect 5135 -4714 5143 -4680
rect 5091 -4742 5143 -4714
rect 5197 -4691 5205 -4657
rect 5239 -4691 5249 -4657
rect 5197 -4742 5249 -4691
rect 5279 -4624 5331 -4612
rect 5279 -4658 5289 -4624
rect 5323 -4658 5331 -4624
rect 5482 -4658 5534 -4612
rect 5279 -4692 5331 -4658
rect 5279 -4726 5289 -4692
rect 5323 -4726 5331 -4692
rect 5279 -4742 5331 -4726
rect 5385 -4670 5437 -4658
rect 5385 -4704 5393 -4670
rect 5427 -4704 5437 -4670
rect 5385 -4742 5437 -4704
rect 5467 -4676 5534 -4658
rect 5467 -4710 5490 -4676
rect 5524 -4710 5534 -4676
rect 5467 -4742 5534 -4710
rect 5564 -4646 5616 -4612
rect 5564 -4680 5574 -4646
rect 5608 -4680 5616 -4646
rect 5564 -4742 5616 -4680
rect 5681 -4670 5733 -4658
rect 5681 -4704 5689 -4670
rect 5723 -4704 5733 -4670
rect 5681 -4742 5733 -4704
rect 5763 -4696 5817 -4658
rect 5763 -4730 5773 -4696
rect 5807 -4730 5817 -4696
rect 5763 -4742 5817 -4730
rect 5847 -4670 5899 -4658
rect 5847 -4704 5857 -4670
rect 5891 -4704 5899 -4670
rect 5847 -4742 5899 -4704
rect 5967 -4700 6072 -4658
rect 5967 -4734 5979 -4700
rect 6013 -4734 6072 -4700
rect 5967 -4742 6072 -4734
rect 6102 -4670 6152 -4658
rect 6583 -4658 6633 -4614
rect 6311 -4670 6429 -4658
rect 6102 -4694 6167 -4670
rect 6102 -4728 6112 -4694
rect 6146 -4728 6167 -4694
rect 6102 -4742 6167 -4728
rect 6197 -4694 6263 -4670
rect 6197 -4728 6219 -4694
rect 6253 -4728 6263 -4694
rect 6197 -4742 6263 -4728
rect 6293 -4742 6429 -4670
rect 6459 -4742 6501 -4658
rect 6531 -4696 6633 -4658
rect 6531 -4730 6565 -4696
rect 6599 -4730 6633 -4696
rect 6531 -4742 6633 -4730
rect 6663 -4670 6717 -4614
rect 7313 -4657 7365 -4612
rect 6887 -4670 6937 -4658
rect 6663 -4700 6732 -4670
rect 6663 -4734 6677 -4700
rect 6711 -4734 6732 -4700
rect 6663 -4742 6732 -4734
rect 6762 -4696 6841 -4670
rect 6762 -4730 6787 -4696
rect 6821 -4730 6841 -4696
rect 6762 -4742 6841 -4730
rect 6871 -4742 6937 -4670
rect 6967 -4700 7086 -4658
rect 6967 -4734 6999 -4700
rect 7033 -4734 7086 -4700
rect 6967 -4742 7086 -4734
rect 7116 -4742 7177 -4658
rect 7207 -4680 7259 -4658
rect 7207 -4714 7217 -4680
rect 7251 -4714 7259 -4680
rect 7207 -4742 7259 -4714
rect 7313 -4691 7321 -4657
rect 7355 -4691 7365 -4657
rect 7313 -4742 7365 -4691
rect 7395 -4624 7447 -4612
rect 7395 -4658 7405 -4624
rect 7439 -4658 7447 -4624
rect 7598 -4658 7650 -4612
rect 7395 -4692 7447 -4658
rect 7395 -4726 7405 -4692
rect 7439 -4726 7447 -4692
rect 7395 -4742 7447 -4726
rect 7501 -4670 7553 -4658
rect 7501 -4704 7509 -4670
rect 7543 -4704 7553 -4670
rect 7501 -4742 7553 -4704
rect 7583 -4676 7650 -4658
rect 7583 -4710 7606 -4676
rect 7640 -4710 7650 -4676
rect 7583 -4742 7650 -4710
rect 7680 -4646 7732 -4612
rect 7680 -4680 7690 -4646
rect 7724 -4680 7732 -4646
rect 7680 -4742 7732 -4680
rect 7797 -4670 7849 -4658
rect 7797 -4704 7805 -4670
rect 7839 -4704 7849 -4670
rect 7797 -4742 7849 -4704
rect 7879 -4696 7933 -4658
rect 7879 -4730 7889 -4696
rect 7923 -4730 7933 -4696
rect 7879 -4742 7933 -4730
rect 7963 -4670 8015 -4658
rect 7963 -4704 7973 -4670
rect 8007 -4704 8015 -4670
rect 7963 -4742 8015 -4704
rect 8083 -4700 8188 -4658
rect 8083 -4734 8095 -4700
rect 8129 -4734 8188 -4700
rect 8083 -4742 8188 -4734
rect 8218 -4670 8268 -4658
rect 8699 -4658 8749 -4614
rect 8427 -4670 8545 -4658
rect 8218 -4694 8283 -4670
rect 8218 -4728 8228 -4694
rect 8262 -4728 8283 -4694
rect 8218 -4742 8283 -4728
rect 8313 -4694 8379 -4670
rect 8313 -4728 8335 -4694
rect 8369 -4728 8379 -4694
rect 8313 -4742 8379 -4728
rect 8409 -4742 8545 -4670
rect 8575 -4742 8617 -4658
rect 8647 -4696 8749 -4658
rect 8647 -4730 8681 -4696
rect 8715 -4730 8749 -4696
rect 8647 -4742 8749 -4730
rect 8779 -4670 8833 -4614
rect 9429 -4657 9481 -4612
rect 9003 -4670 9053 -4658
rect 8779 -4700 8848 -4670
rect 8779 -4734 8793 -4700
rect 8827 -4734 8848 -4700
rect 8779 -4742 8848 -4734
rect 8878 -4696 8957 -4670
rect 8878 -4730 8903 -4696
rect 8937 -4730 8957 -4696
rect 8878 -4742 8957 -4730
rect 8987 -4742 9053 -4670
rect 9083 -4700 9202 -4658
rect 9083 -4734 9115 -4700
rect 9149 -4734 9202 -4700
rect 9083 -4742 9202 -4734
rect 9232 -4742 9293 -4658
rect 9323 -4680 9375 -4658
rect 9323 -4714 9333 -4680
rect 9367 -4714 9375 -4680
rect 9323 -4742 9375 -4714
rect 9429 -4691 9437 -4657
rect 9471 -4691 9481 -4657
rect 9429 -4742 9481 -4691
rect 9511 -4624 9563 -4612
rect 9511 -4658 9521 -4624
rect 9555 -4658 9563 -4624
rect 9714 -4658 9766 -4612
rect 9511 -4692 9563 -4658
rect 9511 -4726 9521 -4692
rect 9555 -4726 9563 -4692
rect 9511 -4742 9563 -4726
rect 9617 -4670 9669 -4658
rect 9617 -4704 9625 -4670
rect 9659 -4704 9669 -4670
rect 9617 -4742 9669 -4704
rect 9699 -4676 9766 -4658
rect 9699 -4710 9722 -4676
rect 9756 -4710 9766 -4676
rect 9699 -4742 9766 -4710
rect 9796 -4646 9848 -4612
rect 9796 -4680 9806 -4646
rect 9840 -4680 9848 -4646
rect 9796 -4742 9848 -4680
rect 9913 -4670 9965 -4658
rect 9913 -4704 9921 -4670
rect 9955 -4704 9965 -4670
rect 9913 -4742 9965 -4704
rect 9995 -4696 10049 -4658
rect 9995 -4730 10005 -4696
rect 10039 -4730 10049 -4696
rect 9995 -4742 10049 -4730
rect 10079 -4670 10131 -4658
rect 10079 -4704 10089 -4670
rect 10123 -4704 10131 -4670
rect 10079 -4742 10131 -4704
rect 10199 -4700 10304 -4658
rect 10199 -4734 10211 -4700
rect 10245 -4734 10304 -4700
rect 10199 -4742 10304 -4734
rect 10334 -4670 10384 -4658
rect 10815 -4658 10865 -4614
rect 10543 -4670 10661 -4658
rect 10334 -4694 10399 -4670
rect 10334 -4728 10344 -4694
rect 10378 -4728 10399 -4694
rect 10334 -4742 10399 -4728
rect 10429 -4694 10495 -4670
rect 10429 -4728 10451 -4694
rect 10485 -4728 10495 -4694
rect 10429 -4742 10495 -4728
rect 10525 -4742 10661 -4670
rect 10691 -4742 10733 -4658
rect 10763 -4696 10865 -4658
rect 10763 -4730 10797 -4696
rect 10831 -4730 10865 -4696
rect 10763 -4742 10865 -4730
rect 10895 -4670 10949 -4614
rect 11545 -4657 11597 -4612
rect 11119 -4670 11169 -4658
rect 10895 -4700 10964 -4670
rect 10895 -4734 10909 -4700
rect 10943 -4734 10964 -4700
rect 10895 -4742 10964 -4734
rect 10994 -4696 11073 -4670
rect 10994 -4730 11019 -4696
rect 11053 -4730 11073 -4696
rect 10994 -4742 11073 -4730
rect 11103 -4742 11169 -4670
rect 11199 -4700 11318 -4658
rect 11199 -4734 11231 -4700
rect 11265 -4734 11318 -4700
rect 11199 -4742 11318 -4734
rect 11348 -4742 11409 -4658
rect 11439 -4680 11491 -4658
rect 11439 -4714 11449 -4680
rect 11483 -4714 11491 -4680
rect 11439 -4742 11491 -4714
rect 11545 -4691 11553 -4657
rect 11587 -4691 11597 -4657
rect 11545 -4742 11597 -4691
rect 11627 -4624 11679 -4612
rect 11627 -4658 11637 -4624
rect 11671 -4658 11679 -4624
rect 11830 -4658 11882 -4612
rect 11627 -4692 11679 -4658
rect 11627 -4726 11637 -4692
rect 11671 -4726 11679 -4692
rect 11627 -4742 11679 -4726
rect 11733 -4670 11785 -4658
rect 11733 -4704 11741 -4670
rect 11775 -4704 11785 -4670
rect 11733 -4742 11785 -4704
rect 11815 -4676 11882 -4658
rect 11815 -4710 11838 -4676
rect 11872 -4710 11882 -4676
rect 11815 -4742 11882 -4710
rect 11912 -4646 11964 -4612
rect 11912 -4680 11922 -4646
rect 11956 -4680 11964 -4646
rect 11912 -4742 11964 -4680
rect 12029 -4670 12081 -4658
rect 12029 -4704 12037 -4670
rect 12071 -4704 12081 -4670
rect 12029 -4742 12081 -4704
rect 12111 -4696 12165 -4658
rect 12111 -4730 12121 -4696
rect 12155 -4730 12165 -4696
rect 12111 -4742 12165 -4730
rect 12195 -4670 12247 -4658
rect 12195 -4704 12205 -4670
rect 12239 -4704 12247 -4670
rect 12195 -4742 12247 -4704
rect 12315 -4700 12420 -4658
rect 12315 -4734 12327 -4700
rect 12361 -4734 12420 -4700
rect 12315 -4742 12420 -4734
rect 12450 -4670 12500 -4658
rect 12931 -4658 12981 -4614
rect 12659 -4670 12777 -4658
rect 12450 -4694 12515 -4670
rect 12450 -4728 12460 -4694
rect 12494 -4728 12515 -4694
rect 12450 -4742 12515 -4728
rect 12545 -4694 12611 -4670
rect 12545 -4728 12567 -4694
rect 12601 -4728 12611 -4694
rect 12545 -4742 12611 -4728
rect 12641 -4742 12777 -4670
rect 12807 -4742 12849 -4658
rect 12879 -4696 12981 -4658
rect 12879 -4730 12913 -4696
rect 12947 -4730 12981 -4696
rect 12879 -4742 12981 -4730
rect 13011 -4670 13065 -4614
rect 13661 -4657 13713 -4612
rect 13235 -4670 13285 -4658
rect 13011 -4700 13080 -4670
rect 13011 -4734 13025 -4700
rect 13059 -4734 13080 -4700
rect 13011 -4742 13080 -4734
rect 13110 -4696 13189 -4670
rect 13110 -4730 13135 -4696
rect 13169 -4730 13189 -4696
rect 13110 -4742 13189 -4730
rect 13219 -4742 13285 -4670
rect 13315 -4700 13434 -4658
rect 13315 -4734 13347 -4700
rect 13381 -4734 13434 -4700
rect 13315 -4742 13434 -4734
rect 13464 -4742 13525 -4658
rect 13555 -4680 13607 -4658
rect 13555 -4714 13565 -4680
rect 13599 -4714 13607 -4680
rect 13555 -4742 13607 -4714
rect 13661 -4691 13669 -4657
rect 13703 -4691 13713 -4657
rect 13661 -4742 13713 -4691
rect 13743 -4624 13795 -4612
rect 13743 -4658 13753 -4624
rect 13787 -4658 13795 -4624
rect 13946 -4658 13998 -4612
rect 13743 -4692 13795 -4658
rect 13743 -4726 13753 -4692
rect 13787 -4726 13795 -4692
rect 13743 -4742 13795 -4726
rect 13849 -4670 13901 -4658
rect 13849 -4704 13857 -4670
rect 13891 -4704 13901 -4670
rect 13849 -4742 13901 -4704
rect 13931 -4676 13998 -4658
rect 13931 -4710 13954 -4676
rect 13988 -4710 13998 -4676
rect 13931 -4742 13998 -4710
rect 14028 -4646 14080 -4612
rect 14028 -4680 14038 -4646
rect 14072 -4680 14080 -4646
rect 14028 -4742 14080 -4680
rect 14145 -4670 14197 -4658
rect 14145 -4704 14153 -4670
rect 14187 -4704 14197 -4670
rect 14145 -4742 14197 -4704
rect 14227 -4696 14281 -4658
rect 14227 -4730 14237 -4696
rect 14271 -4730 14281 -4696
rect 14227 -4742 14281 -4730
rect 14311 -4670 14363 -4658
rect 14311 -4704 14321 -4670
rect 14355 -4704 14363 -4670
rect 14311 -4742 14363 -4704
rect 14431 -4700 14536 -4658
rect 14431 -4734 14443 -4700
rect 14477 -4734 14536 -4700
rect 14431 -4742 14536 -4734
rect 14566 -4670 14616 -4658
rect 15047 -4658 15097 -4614
rect 14775 -4670 14893 -4658
rect 14566 -4694 14631 -4670
rect 14566 -4728 14576 -4694
rect 14610 -4728 14631 -4694
rect 14566 -4742 14631 -4728
rect 14661 -4694 14727 -4670
rect 14661 -4728 14683 -4694
rect 14717 -4728 14727 -4694
rect 14661 -4742 14727 -4728
rect 14757 -4742 14893 -4670
rect 14923 -4742 14965 -4658
rect 14995 -4696 15097 -4658
rect 14995 -4730 15029 -4696
rect 15063 -4730 15097 -4696
rect 14995 -4742 15097 -4730
rect 15127 -4670 15181 -4614
rect 15777 -4657 15829 -4612
rect 15351 -4670 15401 -4658
rect 15127 -4700 15196 -4670
rect 15127 -4734 15141 -4700
rect 15175 -4734 15196 -4700
rect 15127 -4742 15196 -4734
rect 15226 -4696 15305 -4670
rect 15226 -4730 15251 -4696
rect 15285 -4730 15305 -4696
rect 15226 -4742 15305 -4730
rect 15335 -4742 15401 -4670
rect 15431 -4700 15550 -4658
rect 15431 -4734 15463 -4700
rect 15497 -4734 15550 -4700
rect 15431 -4742 15550 -4734
rect 15580 -4742 15641 -4658
rect 15671 -4680 15723 -4658
rect 15671 -4714 15681 -4680
rect 15715 -4714 15723 -4680
rect 15671 -4742 15723 -4714
rect 15777 -4691 15785 -4657
rect 15819 -4691 15829 -4657
rect 15777 -4742 15829 -4691
rect 15859 -4624 15911 -4612
rect 15859 -4658 15869 -4624
rect 15903 -4658 15911 -4624
rect 16062 -4658 16114 -4612
rect 15859 -4692 15911 -4658
rect 15859 -4726 15869 -4692
rect 15903 -4726 15911 -4692
rect 15859 -4742 15911 -4726
rect 15965 -4670 16017 -4658
rect 15965 -4704 15973 -4670
rect 16007 -4704 16017 -4670
rect 15965 -4742 16017 -4704
rect 16047 -4676 16114 -4658
rect 16047 -4710 16070 -4676
rect 16104 -4710 16114 -4676
rect 16047 -4742 16114 -4710
rect 16144 -4646 16196 -4612
rect 16144 -4680 16154 -4646
rect 16188 -4680 16196 -4646
rect 16144 -4742 16196 -4680
rect 16261 -4670 16313 -4658
rect 16261 -4704 16269 -4670
rect 16303 -4704 16313 -4670
rect 16261 -4742 16313 -4704
rect 16343 -4696 16397 -4658
rect 16343 -4730 16353 -4696
rect 16387 -4730 16397 -4696
rect 16343 -4742 16397 -4730
rect 16427 -4670 16479 -4658
rect 16427 -4704 16437 -4670
rect 16471 -4704 16479 -4670
rect 16427 -4742 16479 -4704
rect 16547 -4700 16652 -4658
rect 16547 -4734 16559 -4700
rect 16593 -4734 16652 -4700
rect 16547 -4742 16652 -4734
rect 16682 -4670 16732 -4658
rect 17163 -4658 17213 -4614
rect 16891 -4670 17009 -4658
rect 16682 -4694 16747 -4670
rect 16682 -4728 16692 -4694
rect 16726 -4728 16747 -4694
rect 16682 -4742 16747 -4728
rect 16777 -4694 16843 -4670
rect 16777 -4728 16799 -4694
rect 16833 -4728 16843 -4694
rect 16777 -4742 16843 -4728
rect 16873 -4742 17009 -4670
rect 17039 -4742 17081 -4658
rect 17111 -4696 17213 -4658
rect 17111 -4730 17145 -4696
rect 17179 -4730 17213 -4696
rect 17111 -4742 17213 -4730
rect 17243 -4670 17297 -4614
rect 17893 -4657 17945 -4612
rect 17467 -4670 17517 -4658
rect 17243 -4700 17312 -4670
rect 17243 -4734 17257 -4700
rect 17291 -4734 17312 -4700
rect 17243 -4742 17312 -4734
rect 17342 -4696 17421 -4670
rect 17342 -4730 17367 -4696
rect 17401 -4730 17421 -4696
rect 17342 -4742 17421 -4730
rect 17451 -4742 17517 -4670
rect 17547 -4700 17666 -4658
rect 17547 -4734 17579 -4700
rect 17613 -4734 17666 -4700
rect 17547 -4742 17666 -4734
rect 17696 -4742 17757 -4658
rect 17787 -4680 17839 -4658
rect 17787 -4714 17797 -4680
rect 17831 -4714 17839 -4680
rect 17787 -4742 17839 -4714
rect 17893 -4691 17901 -4657
rect 17935 -4691 17945 -4657
rect 17893 -4742 17945 -4691
rect 17975 -4624 18027 -4612
rect 17975 -4658 17985 -4624
rect 18019 -4658 18027 -4624
rect 18178 -4658 18230 -4612
rect 17975 -4692 18027 -4658
rect 17975 -4726 17985 -4692
rect 18019 -4726 18027 -4692
rect 17975 -4742 18027 -4726
rect 18081 -4670 18133 -4658
rect 18081 -4704 18089 -4670
rect 18123 -4704 18133 -4670
rect 18081 -4742 18133 -4704
rect 18163 -4676 18230 -4658
rect 18163 -4710 18186 -4676
rect 18220 -4710 18230 -4676
rect 18163 -4742 18230 -4710
rect 18260 -4646 18312 -4612
rect 18260 -4680 18270 -4646
rect 18304 -4680 18312 -4646
rect 18260 -4742 18312 -4680
rect 18377 -4670 18429 -4658
rect 18377 -4704 18385 -4670
rect 18419 -4704 18429 -4670
rect 18377 -4742 18429 -4704
rect 18459 -4696 18513 -4658
rect 18459 -4730 18469 -4696
rect 18503 -4730 18513 -4696
rect 18459 -4742 18513 -4730
rect 18543 -4670 18595 -4658
rect 18543 -4704 18553 -4670
rect 18587 -4704 18595 -4670
rect 18543 -4742 18595 -4704
rect 18663 -4700 18768 -4658
rect 18663 -4734 18675 -4700
rect 18709 -4734 18768 -4700
rect 18663 -4742 18768 -4734
rect 18798 -4670 18848 -4658
rect 19279 -4658 19329 -4614
rect 19007 -4670 19125 -4658
rect 18798 -4694 18863 -4670
rect 18798 -4728 18808 -4694
rect 18842 -4728 18863 -4694
rect 18798 -4742 18863 -4728
rect 18893 -4694 18959 -4670
rect 18893 -4728 18915 -4694
rect 18949 -4728 18959 -4694
rect 18893 -4742 18959 -4728
rect 18989 -4742 19125 -4670
rect 19155 -4742 19197 -4658
rect 19227 -4696 19329 -4658
rect 19227 -4730 19261 -4696
rect 19295 -4730 19329 -4696
rect 19227 -4742 19329 -4730
rect 19359 -4670 19413 -4614
rect 20009 -4657 20061 -4612
rect 19583 -4670 19633 -4658
rect 19359 -4700 19428 -4670
rect 19359 -4734 19373 -4700
rect 19407 -4734 19428 -4700
rect 19359 -4742 19428 -4734
rect 19458 -4696 19537 -4670
rect 19458 -4730 19483 -4696
rect 19517 -4730 19537 -4696
rect 19458 -4742 19537 -4730
rect 19567 -4742 19633 -4670
rect 19663 -4700 19782 -4658
rect 19663 -4734 19695 -4700
rect 19729 -4734 19782 -4700
rect 19663 -4742 19782 -4734
rect 19812 -4742 19873 -4658
rect 19903 -4680 19955 -4658
rect 19903 -4714 19913 -4680
rect 19947 -4714 19955 -4680
rect 19903 -4742 19955 -4714
rect 20009 -4691 20017 -4657
rect 20051 -4691 20061 -4657
rect 20009 -4742 20061 -4691
rect 20091 -4624 20143 -4612
rect 20091 -4658 20101 -4624
rect 20135 -4658 20143 -4624
rect 20294 -4658 20346 -4612
rect 20091 -4692 20143 -4658
rect 20091 -4726 20101 -4692
rect 20135 -4726 20143 -4692
rect 20091 -4742 20143 -4726
rect 20197 -4670 20249 -4658
rect 20197 -4704 20205 -4670
rect 20239 -4704 20249 -4670
rect 20197 -4742 20249 -4704
rect 20279 -4676 20346 -4658
rect 20279 -4710 20302 -4676
rect 20336 -4710 20346 -4676
rect 20279 -4742 20346 -4710
rect 20376 -4646 20428 -4612
rect 20376 -4680 20386 -4646
rect 20420 -4680 20428 -4646
rect 20376 -4742 20428 -4680
rect 20493 -4670 20545 -4658
rect 20493 -4704 20501 -4670
rect 20535 -4704 20545 -4670
rect 20493 -4742 20545 -4704
rect 20575 -4696 20629 -4658
rect 20575 -4730 20585 -4696
rect 20619 -4730 20629 -4696
rect 20575 -4742 20629 -4730
rect 20659 -4670 20711 -4658
rect 20659 -4704 20669 -4670
rect 20703 -4704 20711 -4670
rect 20659 -4742 20711 -4704
rect 20779 -4700 20884 -4658
rect 20779 -4734 20791 -4700
rect 20825 -4734 20884 -4700
rect 20779 -4742 20884 -4734
rect 20914 -4670 20964 -4658
rect 21395 -4658 21445 -4614
rect 21123 -4670 21241 -4658
rect 20914 -4694 20979 -4670
rect 20914 -4728 20924 -4694
rect 20958 -4728 20979 -4694
rect 20914 -4742 20979 -4728
rect 21009 -4694 21075 -4670
rect 21009 -4728 21031 -4694
rect 21065 -4728 21075 -4694
rect 21009 -4742 21075 -4728
rect 21105 -4742 21241 -4670
rect 21271 -4742 21313 -4658
rect 21343 -4696 21445 -4658
rect 21343 -4730 21377 -4696
rect 21411 -4730 21445 -4696
rect 21343 -4742 21445 -4730
rect 21475 -4670 21529 -4614
rect 22125 -4657 22177 -4612
rect 21699 -4670 21749 -4658
rect 21475 -4700 21544 -4670
rect 21475 -4734 21489 -4700
rect 21523 -4734 21544 -4700
rect 21475 -4742 21544 -4734
rect 21574 -4696 21653 -4670
rect 21574 -4730 21599 -4696
rect 21633 -4730 21653 -4696
rect 21574 -4742 21653 -4730
rect 21683 -4742 21749 -4670
rect 21779 -4700 21898 -4658
rect 21779 -4734 21811 -4700
rect 21845 -4734 21898 -4700
rect 21779 -4742 21898 -4734
rect 21928 -4742 21989 -4658
rect 22019 -4680 22071 -4658
rect 22019 -4714 22029 -4680
rect 22063 -4714 22071 -4680
rect 22019 -4742 22071 -4714
rect 22125 -4691 22133 -4657
rect 22167 -4691 22177 -4657
rect 22125 -4742 22177 -4691
rect 22207 -4624 22259 -4612
rect 22207 -4658 22217 -4624
rect 22251 -4658 22259 -4624
rect 22410 -4658 22462 -4612
rect 22207 -4692 22259 -4658
rect 22207 -4726 22217 -4692
rect 22251 -4726 22259 -4692
rect 22207 -4742 22259 -4726
rect 22313 -4670 22365 -4658
rect 22313 -4704 22321 -4670
rect 22355 -4704 22365 -4670
rect 22313 -4742 22365 -4704
rect 22395 -4676 22462 -4658
rect 22395 -4710 22418 -4676
rect 22452 -4710 22462 -4676
rect 22395 -4742 22462 -4710
rect 22492 -4646 22544 -4612
rect 22492 -4680 22502 -4646
rect 22536 -4680 22544 -4646
rect 22492 -4742 22544 -4680
rect 22609 -4670 22661 -4658
rect 22609 -4704 22617 -4670
rect 22651 -4704 22661 -4670
rect 22609 -4742 22661 -4704
rect 22691 -4696 22745 -4658
rect 22691 -4730 22701 -4696
rect 22735 -4730 22745 -4696
rect 22691 -4742 22745 -4730
rect 22775 -4670 22827 -4658
rect 22775 -4704 22785 -4670
rect 22819 -4704 22827 -4670
rect 22775 -4742 22827 -4704
rect 22895 -4700 23000 -4658
rect 22895 -4734 22907 -4700
rect 22941 -4734 23000 -4700
rect 22895 -4742 23000 -4734
rect 23030 -4670 23080 -4658
rect 23511 -4658 23561 -4614
rect 23239 -4670 23357 -4658
rect 23030 -4694 23095 -4670
rect 23030 -4728 23040 -4694
rect 23074 -4728 23095 -4694
rect 23030 -4742 23095 -4728
rect 23125 -4694 23191 -4670
rect 23125 -4728 23147 -4694
rect 23181 -4728 23191 -4694
rect 23125 -4742 23191 -4728
rect 23221 -4742 23357 -4670
rect 23387 -4742 23429 -4658
rect 23459 -4696 23561 -4658
rect 23459 -4730 23493 -4696
rect 23527 -4730 23561 -4696
rect 23459 -4742 23561 -4730
rect 23591 -4670 23645 -4614
rect 24241 -4657 24293 -4612
rect 23815 -4670 23865 -4658
rect 23591 -4700 23660 -4670
rect 23591 -4734 23605 -4700
rect 23639 -4734 23660 -4700
rect 23591 -4742 23660 -4734
rect 23690 -4696 23769 -4670
rect 23690 -4730 23715 -4696
rect 23749 -4730 23769 -4696
rect 23690 -4742 23769 -4730
rect 23799 -4742 23865 -4670
rect 23895 -4700 24014 -4658
rect 23895 -4734 23927 -4700
rect 23961 -4734 24014 -4700
rect 23895 -4742 24014 -4734
rect 24044 -4742 24105 -4658
rect 24135 -4680 24187 -4658
rect 24135 -4714 24145 -4680
rect 24179 -4714 24187 -4680
rect 24135 -4742 24187 -4714
rect 24241 -4691 24249 -4657
rect 24283 -4691 24293 -4657
rect 24241 -4742 24293 -4691
rect 24323 -4624 24375 -4612
rect 24323 -4658 24333 -4624
rect 24367 -4658 24375 -4624
rect 24526 -4658 24578 -4612
rect 24323 -4692 24375 -4658
rect 24323 -4726 24333 -4692
rect 24367 -4726 24375 -4692
rect 24323 -4742 24375 -4726
rect 24429 -4670 24481 -4658
rect 24429 -4704 24437 -4670
rect 24471 -4704 24481 -4670
rect 24429 -4742 24481 -4704
rect 24511 -4676 24578 -4658
rect 24511 -4710 24534 -4676
rect 24568 -4710 24578 -4676
rect 24511 -4742 24578 -4710
rect 24608 -4646 24660 -4612
rect 24608 -4680 24618 -4646
rect 24652 -4680 24660 -4646
rect 24608 -4742 24660 -4680
rect 24725 -4670 24777 -4658
rect 24725 -4704 24733 -4670
rect 24767 -4704 24777 -4670
rect 24725 -4742 24777 -4704
rect 24807 -4696 24861 -4658
rect 24807 -4730 24817 -4696
rect 24851 -4730 24861 -4696
rect 24807 -4742 24861 -4730
rect 24891 -4670 24943 -4658
rect 24891 -4704 24901 -4670
rect 24935 -4704 24943 -4670
rect 24891 -4742 24943 -4704
rect 25011 -4700 25116 -4658
rect 25011 -4734 25023 -4700
rect 25057 -4734 25116 -4700
rect 25011 -4742 25116 -4734
rect 25146 -4670 25196 -4658
rect 25627 -4658 25677 -4614
rect 25355 -4670 25473 -4658
rect 25146 -4694 25211 -4670
rect 25146 -4728 25156 -4694
rect 25190 -4728 25211 -4694
rect 25146 -4742 25211 -4728
rect 25241 -4694 25307 -4670
rect 25241 -4728 25263 -4694
rect 25297 -4728 25307 -4694
rect 25241 -4742 25307 -4728
rect 25337 -4742 25473 -4670
rect 25503 -4742 25545 -4658
rect 25575 -4696 25677 -4658
rect 25575 -4730 25609 -4696
rect 25643 -4730 25677 -4696
rect 25575 -4742 25677 -4730
rect 25707 -4670 25761 -4614
rect 26357 -4657 26409 -4612
rect 25931 -4670 25981 -4658
rect 25707 -4700 25776 -4670
rect 25707 -4734 25721 -4700
rect 25755 -4734 25776 -4700
rect 25707 -4742 25776 -4734
rect 25806 -4696 25885 -4670
rect 25806 -4730 25831 -4696
rect 25865 -4730 25885 -4696
rect 25806 -4742 25885 -4730
rect 25915 -4742 25981 -4670
rect 26011 -4700 26130 -4658
rect 26011 -4734 26043 -4700
rect 26077 -4734 26130 -4700
rect 26011 -4742 26130 -4734
rect 26160 -4742 26221 -4658
rect 26251 -4680 26303 -4658
rect 26251 -4714 26261 -4680
rect 26295 -4714 26303 -4680
rect 26251 -4742 26303 -4714
rect 26357 -4691 26365 -4657
rect 26399 -4691 26409 -4657
rect 26357 -4742 26409 -4691
rect 26439 -4624 26491 -4612
rect 26439 -4658 26449 -4624
rect 26483 -4658 26491 -4624
rect 26642 -4658 26694 -4612
rect 26439 -4692 26491 -4658
rect 26439 -4726 26449 -4692
rect 26483 -4726 26491 -4692
rect 26439 -4742 26491 -4726
rect 26545 -4670 26597 -4658
rect 26545 -4704 26553 -4670
rect 26587 -4704 26597 -4670
rect 26545 -4742 26597 -4704
rect 26627 -4676 26694 -4658
rect 26627 -4710 26650 -4676
rect 26684 -4710 26694 -4676
rect 26627 -4742 26694 -4710
rect 26724 -4646 26776 -4612
rect 26724 -4680 26734 -4646
rect 26768 -4680 26776 -4646
rect 26724 -4742 26776 -4680
rect 26841 -4670 26893 -4658
rect 26841 -4704 26849 -4670
rect 26883 -4704 26893 -4670
rect 26841 -4742 26893 -4704
rect 26923 -4696 26977 -4658
rect 26923 -4730 26933 -4696
rect 26967 -4730 26977 -4696
rect 26923 -4742 26977 -4730
rect 27007 -4670 27059 -4658
rect 27007 -4704 27017 -4670
rect 27051 -4704 27059 -4670
rect 27007 -4742 27059 -4704
rect 27127 -4700 27232 -4658
rect 27127 -4734 27139 -4700
rect 27173 -4734 27232 -4700
rect 27127 -4742 27232 -4734
rect 27262 -4670 27312 -4658
rect 27743 -4658 27793 -4614
rect 27471 -4670 27589 -4658
rect 27262 -4694 27327 -4670
rect 27262 -4728 27272 -4694
rect 27306 -4728 27327 -4694
rect 27262 -4742 27327 -4728
rect 27357 -4694 27423 -4670
rect 27357 -4728 27379 -4694
rect 27413 -4728 27423 -4694
rect 27357 -4742 27423 -4728
rect 27453 -4742 27589 -4670
rect 27619 -4742 27661 -4658
rect 27691 -4696 27793 -4658
rect 27691 -4730 27725 -4696
rect 27759 -4730 27793 -4696
rect 27691 -4742 27793 -4730
rect 27823 -4670 27877 -4614
rect 28473 -4657 28525 -4612
rect 28047 -4670 28097 -4658
rect 27823 -4700 27892 -4670
rect 27823 -4734 27837 -4700
rect 27871 -4734 27892 -4700
rect 27823 -4742 27892 -4734
rect 27922 -4696 28001 -4670
rect 27922 -4730 27947 -4696
rect 27981 -4730 28001 -4696
rect 27922 -4742 28001 -4730
rect 28031 -4742 28097 -4670
rect 28127 -4700 28246 -4658
rect 28127 -4734 28159 -4700
rect 28193 -4734 28246 -4700
rect 28127 -4742 28246 -4734
rect 28276 -4742 28337 -4658
rect 28367 -4680 28419 -4658
rect 28367 -4714 28377 -4680
rect 28411 -4714 28419 -4680
rect 28367 -4742 28419 -4714
rect 28473 -4691 28481 -4657
rect 28515 -4691 28525 -4657
rect 28473 -4742 28525 -4691
rect 28555 -4624 28607 -4612
rect 28555 -4658 28565 -4624
rect 28599 -4658 28607 -4624
rect 28758 -4658 28810 -4612
rect 28555 -4692 28607 -4658
rect 28555 -4726 28565 -4692
rect 28599 -4726 28607 -4692
rect 28555 -4742 28607 -4726
rect 28661 -4670 28713 -4658
rect 28661 -4704 28669 -4670
rect 28703 -4704 28713 -4670
rect 28661 -4742 28713 -4704
rect 28743 -4676 28810 -4658
rect 28743 -4710 28766 -4676
rect 28800 -4710 28810 -4676
rect 28743 -4742 28810 -4710
rect 28840 -4646 28892 -4612
rect 28840 -4680 28850 -4646
rect 28884 -4680 28892 -4646
rect 28840 -4742 28892 -4680
rect 28957 -4670 29009 -4658
rect 28957 -4704 28965 -4670
rect 28999 -4704 29009 -4670
rect 28957 -4742 29009 -4704
rect 29039 -4696 29093 -4658
rect 29039 -4730 29049 -4696
rect 29083 -4730 29093 -4696
rect 29039 -4742 29093 -4730
rect 29123 -4670 29175 -4658
rect 29123 -4704 29133 -4670
rect 29167 -4704 29175 -4670
rect 29123 -4742 29175 -4704
rect 29243 -4700 29348 -4658
rect 29243 -4734 29255 -4700
rect 29289 -4734 29348 -4700
rect 29243 -4742 29348 -4734
rect 29378 -4670 29428 -4658
rect 29859 -4658 29909 -4614
rect 29587 -4670 29705 -4658
rect 29378 -4694 29443 -4670
rect 29378 -4728 29388 -4694
rect 29422 -4728 29443 -4694
rect 29378 -4742 29443 -4728
rect 29473 -4694 29539 -4670
rect 29473 -4728 29495 -4694
rect 29529 -4728 29539 -4694
rect 29473 -4742 29539 -4728
rect 29569 -4742 29705 -4670
rect 29735 -4742 29777 -4658
rect 29807 -4696 29909 -4658
rect 29807 -4730 29841 -4696
rect 29875 -4730 29909 -4696
rect 29807 -4742 29909 -4730
rect 29939 -4670 29993 -4614
rect 30589 -4657 30641 -4612
rect 30163 -4670 30213 -4658
rect 29939 -4700 30008 -4670
rect 29939 -4734 29953 -4700
rect 29987 -4734 30008 -4700
rect 29939 -4742 30008 -4734
rect 30038 -4696 30117 -4670
rect 30038 -4730 30063 -4696
rect 30097 -4730 30117 -4696
rect 30038 -4742 30117 -4730
rect 30147 -4742 30213 -4670
rect 30243 -4700 30362 -4658
rect 30243 -4734 30275 -4700
rect 30309 -4734 30362 -4700
rect 30243 -4742 30362 -4734
rect 30392 -4742 30453 -4658
rect 30483 -4680 30535 -4658
rect 30483 -4714 30493 -4680
rect 30527 -4714 30535 -4680
rect 30483 -4742 30535 -4714
rect 30589 -4691 30597 -4657
rect 30631 -4691 30641 -4657
rect 30589 -4742 30641 -4691
rect 30671 -4624 30723 -4612
rect 30671 -4658 30681 -4624
rect 30715 -4658 30723 -4624
rect 30874 -4658 30926 -4612
rect 30671 -4692 30723 -4658
rect 30671 -4726 30681 -4692
rect 30715 -4726 30723 -4692
rect 30671 -4742 30723 -4726
rect 30777 -4670 30829 -4658
rect 30777 -4704 30785 -4670
rect 30819 -4704 30829 -4670
rect 30777 -4742 30829 -4704
rect 30859 -4676 30926 -4658
rect 30859 -4710 30882 -4676
rect 30916 -4710 30926 -4676
rect 30859 -4742 30926 -4710
rect 30956 -4646 31008 -4612
rect 30956 -4680 30966 -4646
rect 31000 -4680 31008 -4646
rect 30956 -4742 31008 -4680
rect 31073 -4670 31125 -4658
rect 31073 -4704 31081 -4670
rect 31115 -4704 31125 -4670
rect 31073 -4742 31125 -4704
rect 31155 -4696 31209 -4658
rect 31155 -4730 31165 -4696
rect 31199 -4730 31209 -4696
rect 31155 -4742 31209 -4730
rect 31239 -4670 31291 -4658
rect 31239 -4704 31249 -4670
rect 31283 -4704 31291 -4670
rect 31239 -4742 31291 -4704
rect 31359 -4700 31464 -4658
rect 31359 -4734 31371 -4700
rect 31405 -4734 31464 -4700
rect 31359 -4742 31464 -4734
rect 31494 -4670 31544 -4658
rect 31975 -4658 32025 -4614
rect 31703 -4670 31821 -4658
rect 31494 -4694 31559 -4670
rect 31494 -4728 31504 -4694
rect 31538 -4728 31559 -4694
rect 31494 -4742 31559 -4728
rect 31589 -4694 31655 -4670
rect 31589 -4728 31611 -4694
rect 31645 -4728 31655 -4694
rect 31589 -4742 31655 -4728
rect 31685 -4742 31821 -4670
rect 31851 -4742 31893 -4658
rect 31923 -4696 32025 -4658
rect 31923 -4730 31957 -4696
rect 31991 -4730 32025 -4696
rect 31923 -4742 32025 -4730
rect 32055 -4670 32109 -4614
rect 32705 -4657 32757 -4612
rect 32279 -4670 32329 -4658
rect 32055 -4700 32124 -4670
rect 32055 -4734 32069 -4700
rect 32103 -4734 32124 -4700
rect 32055 -4742 32124 -4734
rect 32154 -4696 32233 -4670
rect 32154 -4730 32179 -4696
rect 32213 -4730 32233 -4696
rect 32154 -4742 32233 -4730
rect 32263 -4742 32329 -4670
rect 32359 -4700 32478 -4658
rect 32359 -4734 32391 -4700
rect 32425 -4734 32478 -4700
rect 32359 -4742 32478 -4734
rect 32508 -4742 32569 -4658
rect 32599 -4680 32651 -4658
rect 32599 -4714 32609 -4680
rect 32643 -4714 32651 -4680
rect 32599 -4742 32651 -4714
rect 32705 -4691 32713 -4657
rect 32747 -4691 32757 -4657
rect 32705 -4742 32757 -4691
rect 32787 -4624 32839 -4612
rect 32787 -4658 32797 -4624
rect 32831 -4658 32839 -4624
rect 32990 -4658 33042 -4612
rect 32787 -4692 32839 -4658
rect 32787 -4726 32797 -4692
rect 32831 -4726 32839 -4692
rect 32787 -4742 32839 -4726
rect 32893 -4670 32945 -4658
rect 32893 -4704 32901 -4670
rect 32935 -4704 32945 -4670
rect 32893 -4742 32945 -4704
rect 32975 -4676 33042 -4658
rect 32975 -4710 32998 -4676
rect 33032 -4710 33042 -4676
rect 32975 -4742 33042 -4710
rect 33072 -4646 33124 -4612
rect 33072 -4680 33082 -4646
rect 33116 -4680 33124 -4646
rect 33072 -4742 33124 -4680
rect 4357 -7635 4415 -7623
rect 4357 -9011 4369 -7635
rect 4403 -9011 4415 -7635
rect 4357 -9023 4415 -9011
rect 6015 -7635 6073 -7623
rect 6015 -9011 6027 -7635
rect 6061 -9011 6073 -7635
rect 6015 -9023 6073 -9011
rect 7673 -7635 7731 -7623
rect 7673 -9011 7685 -7635
rect 7719 -9011 7731 -7635
rect 7673 -9023 7731 -9011
rect 4357 -9145 4415 -9133
rect 4357 -10521 4369 -9145
rect 4403 -10521 4415 -9145
rect 4357 -10533 4415 -10521
rect 6015 -9145 6073 -9133
rect 6015 -10521 6027 -9145
rect 6061 -10521 6073 -9145
rect 6015 -10533 6073 -10521
rect 7673 -9145 7731 -9133
rect 7673 -10521 7685 -9145
rect 7719 -10521 7731 -9145
rect 7673 -10533 7731 -10521
rect 4357 -10655 4415 -10643
rect 4357 -12031 4369 -10655
rect 4403 -12031 4415 -10655
rect 4357 -12043 4415 -12031
rect 6015 -10655 6073 -10643
rect 6015 -12031 6027 -10655
rect 6061 -12031 6073 -10655
rect 6015 -12043 6073 -12031
rect 7673 -10655 7731 -10643
rect 7673 -12031 7685 -10655
rect 7719 -12031 7731 -10655
rect 7673 -12043 7731 -12031
rect 4357 -12165 4415 -12153
rect 4357 -13541 4369 -12165
rect 4403 -13541 4415 -12165
rect 4357 -13553 4415 -13541
rect 6015 -12165 6073 -12153
rect 6015 -13541 6027 -12165
rect 6061 -13541 6073 -12165
rect 6015 -13553 6073 -13541
rect 7673 -12165 7731 -12153
rect 7673 -13541 7685 -12165
rect 7719 -13541 7731 -12165
rect 7673 -13553 7731 -13541
rect 4357 -13675 4415 -13663
rect 4357 -15051 4369 -13675
rect 4403 -15051 4415 -13675
rect 4357 -15063 4415 -15051
rect 6015 -13675 6073 -13663
rect 6015 -15051 6027 -13675
rect 6061 -15051 6073 -13675
rect 6015 -15063 6073 -15051
rect 7673 -13675 7731 -13663
rect 7673 -15051 7685 -13675
rect 7719 -15051 7731 -13675
rect 7673 -15063 7731 -15051
rect 4357 -15185 4415 -15173
rect 4357 -16561 4369 -15185
rect 4403 -16561 4415 -15185
rect 4357 -16573 4415 -16561
rect 6015 -15185 6073 -15173
rect 6015 -16561 6027 -15185
rect 6061 -16561 6073 -15185
rect 6015 -16573 6073 -16561
rect 7673 -15185 7731 -15173
rect 7673 -16561 7685 -15185
rect 7719 -16561 7731 -15185
rect 7673 -16573 7731 -16561
rect 4357 -16695 4415 -16683
rect 4357 -18071 4369 -16695
rect 4403 -18071 4415 -16695
rect 4357 -18083 4415 -18071
rect 6015 -16695 6073 -16683
rect 6015 -18071 6027 -16695
rect 6061 -18071 6073 -16695
rect 6015 -18083 6073 -18071
rect 7673 -16695 7731 -16683
rect 7673 -18071 7685 -16695
rect 7719 -18071 7731 -16695
rect 7673 -18083 7731 -18071
rect 4357 -18205 4415 -18193
rect 4357 -19581 4369 -18205
rect 4403 -19581 4415 -18205
rect 4357 -19593 4415 -19581
rect 6015 -18205 6073 -18193
rect 6015 -19581 6027 -18205
rect 6061 -19581 6073 -18205
rect 6015 -19593 6073 -19581
rect 7673 -18205 7731 -18193
rect 7673 -19581 7685 -18205
rect 7719 -19581 7731 -18205
rect 7673 -19593 7731 -19581
rect 4357 -19715 4415 -19703
rect 4357 -21091 4369 -19715
rect 4403 -21091 4415 -19715
rect 4357 -21103 4415 -21091
rect 6015 -19715 6073 -19703
rect 6015 -21091 6027 -19715
rect 6061 -21091 6073 -19715
rect 6015 -21103 6073 -21091
rect 7673 -19715 7731 -19703
rect 7673 -21091 7685 -19715
rect 7719 -21091 7731 -19715
rect 7673 -21103 7731 -21091
rect 4357 -21225 4415 -21213
rect 4357 -22601 4369 -21225
rect 4403 -22601 4415 -21225
rect 4357 -22613 4415 -22601
rect 6015 -21225 6073 -21213
rect 6015 -22601 6027 -21225
rect 6061 -22601 6073 -21225
rect 6015 -22613 6073 -22601
rect 7673 -21225 7731 -21213
rect 7673 -22601 7685 -21225
rect 7719 -22601 7731 -21225
rect 7673 -22613 7731 -22601
rect 4357 -22735 4415 -22723
rect 4357 -24111 4369 -22735
rect 4403 -24111 4415 -22735
rect 4357 -24123 4415 -24111
rect 6015 -22735 6073 -22723
rect 6015 -24111 6027 -22735
rect 6061 -24111 6073 -22735
rect 6015 -24123 6073 -24111
rect 7673 -22735 7731 -22723
rect 7673 -24111 7685 -22735
rect 7719 -24111 7731 -22735
rect 7673 -24123 7731 -24111
rect 4357 -24245 4415 -24233
rect 4357 -25621 4369 -24245
rect 4403 -25621 4415 -24245
rect 4357 -25633 4415 -25621
rect 6015 -24245 6073 -24233
rect 6015 -25621 6027 -24245
rect 6061 -25621 6073 -24245
rect 6015 -25633 6073 -25621
rect 7673 -24245 7731 -24233
rect 7673 -25621 7685 -24245
rect 7719 -25621 7731 -24245
rect 7673 -25633 7731 -25621
rect 9101 -9648 9159 -9636
rect 9101 -9684 9113 -9648
rect 9147 -9684 9159 -9648
rect 9101 -9718 9159 -9684
rect 9101 -9754 9113 -9718
rect 9147 -9754 9159 -9718
rect 9101 -9788 9159 -9754
rect 9101 -9824 9113 -9788
rect 9147 -9824 9159 -9788
rect 9101 -9836 9159 -9824
rect 9359 -9648 9417 -9636
rect 9359 -9684 9371 -9648
rect 9405 -9684 9417 -9648
rect 9359 -9718 9417 -9684
rect 9359 -9754 9371 -9718
rect 9405 -9754 9417 -9718
rect 9359 -9788 9417 -9754
rect 9359 -9824 9371 -9788
rect 9405 -9824 9417 -9788
rect 9359 -9836 9417 -9824
rect 9617 -9648 9675 -9636
rect 9617 -9684 9629 -9648
rect 9663 -9684 9675 -9648
rect 9617 -9718 9675 -9684
rect 9617 -9754 9629 -9718
rect 9663 -9754 9675 -9718
rect 9617 -9789 9675 -9754
rect 9617 -9825 9629 -9789
rect 9663 -9825 9675 -9789
rect 9617 -9836 9675 -9825
rect 9875 -9648 9933 -9636
rect 9875 -9684 9887 -9648
rect 9921 -9684 9933 -9648
rect 9875 -9718 9933 -9684
rect 9875 -9754 9887 -9718
rect 9921 -9754 9933 -9718
rect 9875 -9788 9933 -9754
rect 9875 -9824 9887 -9788
rect 9921 -9824 9933 -9788
rect 9875 -9836 9933 -9824
rect 10133 -9648 10191 -9636
rect 10133 -9684 10145 -9648
rect 10179 -9684 10191 -9648
rect 10133 -9718 10191 -9684
rect 10133 -9754 10145 -9718
rect 10179 -9754 10191 -9718
rect 10133 -9788 10191 -9754
rect 10133 -9824 10145 -9788
rect 10179 -9824 10191 -9788
rect 10133 -9836 10191 -9824
rect 10391 -9648 10449 -9636
rect 10391 -9684 10403 -9648
rect 10437 -9684 10449 -9648
rect 10391 -9718 10449 -9684
rect 10391 -9754 10403 -9718
rect 10437 -9754 10449 -9718
rect 10391 -9788 10449 -9754
rect 10391 -9824 10403 -9788
rect 10437 -9824 10449 -9788
rect 10391 -9836 10449 -9824
rect 10649 -9648 10707 -9636
rect 10649 -9684 10661 -9648
rect 10695 -9684 10707 -9648
rect 10649 -9718 10707 -9684
rect 10649 -9754 10661 -9718
rect 10695 -9754 10707 -9718
rect 10649 -9788 10707 -9754
rect 10649 -9824 10661 -9788
rect 10695 -9824 10707 -9788
rect 10649 -9836 10707 -9824
rect 10907 -9648 10965 -9636
rect 10907 -9684 10919 -9648
rect 10953 -9684 10965 -9648
rect 10907 -9718 10965 -9684
rect 10907 -9754 10919 -9718
rect 10953 -9754 10965 -9718
rect 10907 -9788 10965 -9754
rect 10907 -9824 10919 -9788
rect 10953 -9824 10965 -9788
rect 10907 -9836 10965 -9824
rect 11165 -9648 11223 -9636
rect 11165 -9684 11177 -9648
rect 11211 -9684 11223 -9648
rect 11165 -9718 11223 -9684
rect 11165 -9754 11177 -9718
rect 11211 -9754 11223 -9718
rect 11165 -9788 11223 -9754
rect 11165 -9824 11177 -9788
rect 11211 -9824 11223 -9788
rect 11165 -9836 11223 -9824
rect 11771 -9648 11829 -9636
rect 11771 -9684 11783 -9648
rect 11817 -9684 11829 -9648
rect 11771 -9718 11829 -9684
rect 11771 -9754 11783 -9718
rect 11817 -9754 11829 -9718
rect 11771 -9788 11829 -9754
rect 11771 -9824 11783 -9788
rect 11817 -9824 11829 -9788
rect 11771 -9836 11829 -9824
rect 12029 -9648 12087 -9636
rect 12029 -9684 12041 -9648
rect 12075 -9684 12087 -9648
rect 12029 -9718 12087 -9684
rect 12029 -9754 12041 -9718
rect 12075 -9754 12087 -9718
rect 12029 -9788 12087 -9754
rect 12029 -9824 12041 -9788
rect 12075 -9824 12087 -9788
rect 12029 -9836 12087 -9824
rect 12287 -9648 12345 -9636
rect 12287 -9684 12299 -9648
rect 12333 -9684 12345 -9648
rect 12287 -9718 12345 -9684
rect 12287 -9754 12299 -9718
rect 12333 -9754 12345 -9718
rect 12287 -9789 12345 -9754
rect 12287 -9825 12299 -9789
rect 12333 -9825 12345 -9789
rect 12287 -9836 12345 -9825
rect 12545 -9648 12603 -9636
rect 12545 -9684 12557 -9648
rect 12591 -9684 12603 -9648
rect 12545 -9718 12603 -9684
rect 12545 -9754 12557 -9718
rect 12591 -9754 12603 -9718
rect 12545 -9788 12603 -9754
rect 12545 -9824 12557 -9788
rect 12591 -9824 12603 -9788
rect 12545 -9836 12603 -9824
rect 12803 -9648 12861 -9636
rect 12803 -9684 12815 -9648
rect 12849 -9684 12861 -9648
rect 12803 -9718 12861 -9684
rect 12803 -9754 12815 -9718
rect 12849 -9754 12861 -9718
rect 12803 -9788 12861 -9754
rect 12803 -9824 12815 -9788
rect 12849 -9824 12861 -9788
rect 12803 -9836 12861 -9824
rect 13061 -9648 13119 -9636
rect 13061 -9684 13073 -9648
rect 13107 -9684 13119 -9648
rect 13061 -9718 13119 -9684
rect 13061 -9754 13073 -9718
rect 13107 -9754 13119 -9718
rect 13061 -9788 13119 -9754
rect 13061 -9824 13073 -9788
rect 13107 -9824 13119 -9788
rect 13061 -9836 13119 -9824
rect 13319 -9648 13377 -9636
rect 13319 -9684 13331 -9648
rect 13365 -9684 13377 -9648
rect 13319 -9718 13377 -9684
rect 13319 -9754 13331 -9718
rect 13365 -9754 13377 -9718
rect 13319 -9788 13377 -9754
rect 13319 -9824 13331 -9788
rect 13365 -9824 13377 -9788
rect 13319 -9836 13377 -9824
rect 13577 -9648 13635 -9636
rect 13577 -9684 13589 -9648
rect 13623 -9684 13635 -9648
rect 13577 -9718 13635 -9684
rect 13577 -9754 13589 -9718
rect 13623 -9754 13635 -9718
rect 13577 -9788 13635 -9754
rect 13577 -9824 13589 -9788
rect 13623 -9824 13635 -9788
rect 13577 -9836 13635 -9824
rect 13835 -9648 13893 -9636
rect 13835 -9684 13847 -9648
rect 13881 -9684 13893 -9648
rect 13835 -9718 13893 -9684
rect 13835 -9754 13847 -9718
rect 13881 -9754 13893 -9718
rect 13835 -9788 13893 -9754
rect 13835 -9824 13847 -9788
rect 13881 -9824 13893 -9788
rect 13835 -9836 13893 -9824
rect 14434 -9647 14492 -9635
rect 14434 -9683 14446 -9647
rect 14480 -9683 14492 -9647
rect 14434 -9717 14492 -9683
rect 14434 -9753 14446 -9717
rect 14480 -9753 14492 -9717
rect 14434 -9787 14492 -9753
rect 14434 -9823 14446 -9787
rect 14480 -9823 14492 -9787
rect 14434 -9835 14492 -9823
rect 14692 -9647 14750 -9635
rect 14692 -9683 14704 -9647
rect 14738 -9683 14750 -9647
rect 14692 -9717 14750 -9683
rect 14692 -9753 14704 -9717
rect 14738 -9753 14750 -9717
rect 14692 -9787 14750 -9753
rect 14692 -9823 14704 -9787
rect 14738 -9823 14750 -9787
rect 14692 -9835 14750 -9823
rect 14950 -9647 15008 -9635
rect 14950 -9683 14962 -9647
rect 14996 -9683 15008 -9647
rect 14950 -9717 15008 -9683
rect 14950 -9753 14962 -9717
rect 14996 -9753 15008 -9717
rect 14950 -9788 15008 -9753
rect 14950 -9824 14962 -9788
rect 14996 -9824 15008 -9788
rect 14950 -9835 15008 -9824
rect 15208 -9647 15266 -9635
rect 15208 -9683 15220 -9647
rect 15254 -9683 15266 -9647
rect 15208 -9717 15266 -9683
rect 15208 -9753 15220 -9717
rect 15254 -9753 15266 -9717
rect 15208 -9787 15266 -9753
rect 15208 -9823 15220 -9787
rect 15254 -9823 15266 -9787
rect 15208 -9835 15266 -9823
rect 15466 -9647 15524 -9635
rect 15466 -9683 15478 -9647
rect 15512 -9683 15524 -9647
rect 15466 -9717 15524 -9683
rect 15466 -9753 15478 -9717
rect 15512 -9753 15524 -9717
rect 15466 -9787 15524 -9753
rect 15466 -9823 15478 -9787
rect 15512 -9823 15524 -9787
rect 15466 -9835 15524 -9823
rect 15724 -9647 15782 -9635
rect 15724 -9683 15736 -9647
rect 15770 -9683 15782 -9647
rect 15724 -9717 15782 -9683
rect 15724 -9753 15736 -9717
rect 15770 -9753 15782 -9717
rect 15724 -9787 15782 -9753
rect 15724 -9823 15736 -9787
rect 15770 -9823 15782 -9787
rect 15724 -9835 15782 -9823
rect 15982 -9647 16040 -9635
rect 15982 -9683 15994 -9647
rect 16028 -9683 16040 -9647
rect 15982 -9717 16040 -9683
rect 15982 -9753 15994 -9717
rect 16028 -9753 16040 -9717
rect 15982 -9787 16040 -9753
rect 15982 -9823 15994 -9787
rect 16028 -9823 16040 -9787
rect 15982 -9835 16040 -9823
rect 16240 -9647 16298 -9635
rect 16240 -9683 16252 -9647
rect 16286 -9683 16298 -9647
rect 16240 -9717 16298 -9683
rect 16240 -9753 16252 -9717
rect 16286 -9753 16298 -9717
rect 16240 -9787 16298 -9753
rect 16240 -9823 16252 -9787
rect 16286 -9823 16298 -9787
rect 16240 -9835 16298 -9823
rect 16498 -9647 16556 -9635
rect 16498 -9683 16510 -9647
rect 16544 -9683 16556 -9647
rect 16498 -9717 16556 -9683
rect 16498 -9753 16510 -9717
rect 16544 -9753 16556 -9717
rect 16498 -9787 16556 -9753
rect 16498 -9823 16510 -9787
rect 16544 -9823 16556 -9787
rect 16498 -9835 16556 -9823
rect 9101 -10066 9159 -10054
rect 9101 -10102 9113 -10066
rect 9147 -10102 9159 -10066
rect 9101 -10136 9159 -10102
rect 9101 -10172 9113 -10136
rect 9147 -10172 9159 -10136
rect 9101 -10206 9159 -10172
rect 9101 -10242 9113 -10206
rect 9147 -10242 9159 -10206
rect 9101 -10254 9159 -10242
rect 9359 -10066 9417 -10054
rect 9359 -10102 9371 -10066
rect 9405 -10102 9417 -10066
rect 9359 -10136 9417 -10102
rect 9359 -10172 9371 -10136
rect 9405 -10172 9417 -10136
rect 9359 -10206 9417 -10172
rect 9359 -10242 9371 -10206
rect 9405 -10242 9417 -10206
rect 9359 -10254 9417 -10242
rect 9617 -10066 9675 -10054
rect 9617 -10102 9629 -10066
rect 9663 -10102 9675 -10066
rect 9617 -10136 9675 -10102
rect 9617 -10172 9629 -10136
rect 9663 -10172 9675 -10136
rect 9617 -10207 9675 -10172
rect 9617 -10243 9629 -10207
rect 9663 -10243 9675 -10207
rect 9617 -10254 9675 -10243
rect 9875 -10066 9933 -10054
rect 9875 -10102 9887 -10066
rect 9921 -10102 9933 -10066
rect 9875 -10136 9933 -10102
rect 9875 -10172 9887 -10136
rect 9921 -10172 9933 -10136
rect 9875 -10206 9933 -10172
rect 9875 -10242 9887 -10206
rect 9921 -10242 9933 -10206
rect 9875 -10254 9933 -10242
rect 10133 -10066 10191 -10054
rect 10133 -10102 10145 -10066
rect 10179 -10102 10191 -10066
rect 10133 -10136 10191 -10102
rect 10133 -10172 10145 -10136
rect 10179 -10172 10191 -10136
rect 10133 -10206 10191 -10172
rect 10133 -10242 10145 -10206
rect 10179 -10242 10191 -10206
rect 10133 -10254 10191 -10242
rect 10391 -10066 10449 -10054
rect 10391 -10102 10403 -10066
rect 10437 -10102 10449 -10066
rect 10391 -10136 10449 -10102
rect 10391 -10172 10403 -10136
rect 10437 -10172 10449 -10136
rect 10391 -10206 10449 -10172
rect 10391 -10242 10403 -10206
rect 10437 -10242 10449 -10206
rect 10391 -10254 10449 -10242
rect 10649 -10066 10707 -10054
rect 10649 -10102 10661 -10066
rect 10695 -10102 10707 -10066
rect 10649 -10136 10707 -10102
rect 10649 -10172 10661 -10136
rect 10695 -10172 10707 -10136
rect 10649 -10206 10707 -10172
rect 10649 -10242 10661 -10206
rect 10695 -10242 10707 -10206
rect 10649 -10254 10707 -10242
rect 10907 -10066 10965 -10054
rect 10907 -10102 10919 -10066
rect 10953 -10102 10965 -10066
rect 10907 -10136 10965 -10102
rect 10907 -10172 10919 -10136
rect 10953 -10172 10965 -10136
rect 10907 -10206 10965 -10172
rect 10907 -10242 10919 -10206
rect 10953 -10242 10965 -10206
rect 10907 -10254 10965 -10242
rect 11165 -10066 11223 -10054
rect 11165 -10102 11177 -10066
rect 11211 -10102 11223 -10066
rect 11165 -10136 11223 -10102
rect 11165 -10172 11177 -10136
rect 11211 -10172 11223 -10136
rect 11165 -10206 11223 -10172
rect 11165 -10242 11177 -10206
rect 11211 -10242 11223 -10206
rect 11165 -10254 11223 -10242
rect 11771 -10066 11829 -10054
rect 11771 -10102 11783 -10066
rect 11817 -10102 11829 -10066
rect 11771 -10136 11829 -10102
rect 11771 -10172 11783 -10136
rect 11817 -10172 11829 -10136
rect 11771 -10206 11829 -10172
rect 11771 -10242 11783 -10206
rect 11817 -10242 11829 -10206
rect 11771 -10254 11829 -10242
rect 12029 -10066 12087 -10054
rect 12029 -10102 12041 -10066
rect 12075 -10102 12087 -10066
rect 12029 -10136 12087 -10102
rect 12029 -10172 12041 -10136
rect 12075 -10172 12087 -10136
rect 12029 -10206 12087 -10172
rect 12029 -10242 12041 -10206
rect 12075 -10242 12087 -10206
rect 12029 -10254 12087 -10242
rect 12287 -10066 12345 -10054
rect 12287 -10102 12299 -10066
rect 12333 -10102 12345 -10066
rect 12287 -10136 12345 -10102
rect 12287 -10172 12299 -10136
rect 12333 -10172 12345 -10136
rect 12287 -10207 12345 -10172
rect 12287 -10243 12299 -10207
rect 12333 -10243 12345 -10207
rect 12287 -10254 12345 -10243
rect 12545 -10066 12603 -10054
rect 12545 -10102 12557 -10066
rect 12591 -10102 12603 -10066
rect 12545 -10136 12603 -10102
rect 12545 -10172 12557 -10136
rect 12591 -10172 12603 -10136
rect 12545 -10206 12603 -10172
rect 12545 -10242 12557 -10206
rect 12591 -10242 12603 -10206
rect 12545 -10254 12603 -10242
rect 12803 -10066 12861 -10054
rect 12803 -10102 12815 -10066
rect 12849 -10102 12861 -10066
rect 12803 -10136 12861 -10102
rect 12803 -10172 12815 -10136
rect 12849 -10172 12861 -10136
rect 12803 -10206 12861 -10172
rect 12803 -10242 12815 -10206
rect 12849 -10242 12861 -10206
rect 12803 -10254 12861 -10242
rect 13061 -10066 13119 -10054
rect 13061 -10102 13073 -10066
rect 13107 -10102 13119 -10066
rect 13061 -10136 13119 -10102
rect 13061 -10172 13073 -10136
rect 13107 -10172 13119 -10136
rect 13061 -10206 13119 -10172
rect 13061 -10242 13073 -10206
rect 13107 -10242 13119 -10206
rect 13061 -10254 13119 -10242
rect 13319 -10066 13377 -10054
rect 13319 -10102 13331 -10066
rect 13365 -10102 13377 -10066
rect 13319 -10136 13377 -10102
rect 13319 -10172 13331 -10136
rect 13365 -10172 13377 -10136
rect 13319 -10206 13377 -10172
rect 13319 -10242 13331 -10206
rect 13365 -10242 13377 -10206
rect 13319 -10254 13377 -10242
rect 13577 -10066 13635 -10054
rect 13577 -10102 13589 -10066
rect 13623 -10102 13635 -10066
rect 13577 -10136 13635 -10102
rect 13577 -10172 13589 -10136
rect 13623 -10172 13635 -10136
rect 13577 -10206 13635 -10172
rect 13577 -10242 13589 -10206
rect 13623 -10242 13635 -10206
rect 13577 -10254 13635 -10242
rect 13835 -10066 13893 -10054
rect 13835 -10102 13847 -10066
rect 13881 -10102 13893 -10066
rect 13835 -10136 13893 -10102
rect 13835 -10172 13847 -10136
rect 13881 -10172 13893 -10136
rect 13835 -10206 13893 -10172
rect 13835 -10242 13847 -10206
rect 13881 -10242 13893 -10206
rect 13835 -10254 13893 -10242
rect 14434 -10065 14492 -10053
rect 14434 -10101 14446 -10065
rect 14480 -10101 14492 -10065
rect 14434 -10135 14492 -10101
rect 14434 -10171 14446 -10135
rect 14480 -10171 14492 -10135
rect 14434 -10205 14492 -10171
rect 14434 -10241 14446 -10205
rect 14480 -10241 14492 -10205
rect 14434 -10253 14492 -10241
rect 14692 -10065 14750 -10053
rect 14692 -10101 14704 -10065
rect 14738 -10101 14750 -10065
rect 14692 -10135 14750 -10101
rect 14692 -10171 14704 -10135
rect 14738 -10171 14750 -10135
rect 14692 -10205 14750 -10171
rect 14692 -10241 14704 -10205
rect 14738 -10241 14750 -10205
rect 14692 -10253 14750 -10241
rect 14950 -10065 15008 -10053
rect 14950 -10101 14962 -10065
rect 14996 -10101 15008 -10065
rect 14950 -10135 15008 -10101
rect 14950 -10171 14962 -10135
rect 14996 -10171 15008 -10135
rect 14950 -10206 15008 -10171
rect 14950 -10242 14962 -10206
rect 14996 -10242 15008 -10206
rect 14950 -10253 15008 -10242
rect 15208 -10065 15266 -10053
rect 15208 -10101 15220 -10065
rect 15254 -10101 15266 -10065
rect 15208 -10135 15266 -10101
rect 15208 -10171 15220 -10135
rect 15254 -10171 15266 -10135
rect 15208 -10205 15266 -10171
rect 15208 -10241 15220 -10205
rect 15254 -10241 15266 -10205
rect 15208 -10253 15266 -10241
rect 15466 -10065 15524 -10053
rect 15466 -10101 15478 -10065
rect 15512 -10101 15524 -10065
rect 15466 -10135 15524 -10101
rect 15466 -10171 15478 -10135
rect 15512 -10171 15524 -10135
rect 15466 -10205 15524 -10171
rect 15466 -10241 15478 -10205
rect 15512 -10241 15524 -10205
rect 15466 -10253 15524 -10241
rect 15724 -10065 15782 -10053
rect 15724 -10101 15736 -10065
rect 15770 -10101 15782 -10065
rect 15724 -10135 15782 -10101
rect 15724 -10171 15736 -10135
rect 15770 -10171 15782 -10135
rect 15724 -10205 15782 -10171
rect 15724 -10241 15736 -10205
rect 15770 -10241 15782 -10205
rect 15724 -10253 15782 -10241
rect 15982 -10065 16040 -10053
rect 15982 -10101 15994 -10065
rect 16028 -10101 16040 -10065
rect 15982 -10135 16040 -10101
rect 15982 -10171 15994 -10135
rect 16028 -10171 16040 -10135
rect 15982 -10205 16040 -10171
rect 15982 -10241 15994 -10205
rect 16028 -10241 16040 -10205
rect 15982 -10253 16040 -10241
rect 16240 -10065 16298 -10053
rect 16240 -10101 16252 -10065
rect 16286 -10101 16298 -10065
rect 16240 -10135 16298 -10101
rect 16240 -10171 16252 -10135
rect 16286 -10171 16298 -10135
rect 16240 -10205 16298 -10171
rect 16240 -10241 16252 -10205
rect 16286 -10241 16298 -10205
rect 16240 -10253 16298 -10241
rect 16498 -10065 16556 -10053
rect 16498 -10101 16510 -10065
rect 16544 -10101 16556 -10065
rect 16498 -10135 16556 -10101
rect 16498 -10171 16510 -10135
rect 16544 -10171 16556 -10135
rect 16498 -10205 16556 -10171
rect 16498 -10241 16510 -10205
rect 16544 -10241 16556 -10205
rect 16498 -10253 16556 -10241
rect 9101 -10484 9159 -10472
rect 9101 -10520 9113 -10484
rect 9147 -10520 9159 -10484
rect 9101 -10554 9159 -10520
rect 9101 -10590 9113 -10554
rect 9147 -10590 9159 -10554
rect 9101 -10624 9159 -10590
rect 9101 -10660 9113 -10624
rect 9147 -10660 9159 -10624
rect 9101 -10672 9159 -10660
rect 9359 -10484 9417 -10472
rect 9359 -10520 9371 -10484
rect 9405 -10520 9417 -10484
rect 9359 -10554 9417 -10520
rect 9359 -10590 9371 -10554
rect 9405 -10590 9417 -10554
rect 9359 -10624 9417 -10590
rect 9359 -10660 9371 -10624
rect 9405 -10660 9417 -10624
rect 9359 -10672 9417 -10660
rect 9617 -10484 9675 -10472
rect 9617 -10520 9629 -10484
rect 9663 -10520 9675 -10484
rect 9617 -10554 9675 -10520
rect 9617 -10590 9629 -10554
rect 9663 -10590 9675 -10554
rect 9617 -10625 9675 -10590
rect 9617 -10661 9629 -10625
rect 9663 -10661 9675 -10625
rect 9617 -10672 9675 -10661
rect 9875 -10484 9933 -10472
rect 9875 -10520 9887 -10484
rect 9921 -10520 9933 -10484
rect 9875 -10554 9933 -10520
rect 9875 -10590 9887 -10554
rect 9921 -10590 9933 -10554
rect 9875 -10624 9933 -10590
rect 9875 -10660 9887 -10624
rect 9921 -10660 9933 -10624
rect 9875 -10672 9933 -10660
rect 10133 -10484 10191 -10472
rect 10133 -10520 10145 -10484
rect 10179 -10520 10191 -10484
rect 10133 -10554 10191 -10520
rect 10133 -10590 10145 -10554
rect 10179 -10590 10191 -10554
rect 10133 -10624 10191 -10590
rect 10133 -10660 10145 -10624
rect 10179 -10660 10191 -10624
rect 10133 -10672 10191 -10660
rect 10391 -10484 10449 -10472
rect 10391 -10520 10403 -10484
rect 10437 -10520 10449 -10484
rect 10391 -10554 10449 -10520
rect 10391 -10590 10403 -10554
rect 10437 -10590 10449 -10554
rect 10391 -10624 10449 -10590
rect 10391 -10660 10403 -10624
rect 10437 -10660 10449 -10624
rect 10391 -10672 10449 -10660
rect 10649 -10484 10707 -10472
rect 10649 -10520 10661 -10484
rect 10695 -10520 10707 -10484
rect 10649 -10554 10707 -10520
rect 10649 -10590 10661 -10554
rect 10695 -10590 10707 -10554
rect 10649 -10624 10707 -10590
rect 10649 -10660 10661 -10624
rect 10695 -10660 10707 -10624
rect 10649 -10672 10707 -10660
rect 10907 -10484 10965 -10472
rect 10907 -10520 10919 -10484
rect 10953 -10520 10965 -10484
rect 10907 -10554 10965 -10520
rect 10907 -10590 10919 -10554
rect 10953 -10590 10965 -10554
rect 10907 -10624 10965 -10590
rect 10907 -10660 10919 -10624
rect 10953 -10660 10965 -10624
rect 10907 -10672 10965 -10660
rect 11165 -10484 11223 -10472
rect 11165 -10520 11177 -10484
rect 11211 -10520 11223 -10484
rect 11165 -10554 11223 -10520
rect 11165 -10590 11177 -10554
rect 11211 -10590 11223 -10554
rect 11165 -10624 11223 -10590
rect 11165 -10660 11177 -10624
rect 11211 -10660 11223 -10624
rect 11165 -10672 11223 -10660
rect 11771 -10484 11829 -10472
rect 11771 -10520 11783 -10484
rect 11817 -10520 11829 -10484
rect 11771 -10554 11829 -10520
rect 11771 -10590 11783 -10554
rect 11817 -10590 11829 -10554
rect 11771 -10624 11829 -10590
rect 11771 -10660 11783 -10624
rect 11817 -10660 11829 -10624
rect 11771 -10672 11829 -10660
rect 12029 -10484 12087 -10472
rect 12029 -10520 12041 -10484
rect 12075 -10520 12087 -10484
rect 12029 -10554 12087 -10520
rect 12029 -10590 12041 -10554
rect 12075 -10590 12087 -10554
rect 12029 -10624 12087 -10590
rect 12029 -10660 12041 -10624
rect 12075 -10660 12087 -10624
rect 12029 -10672 12087 -10660
rect 12287 -10484 12345 -10472
rect 12287 -10520 12299 -10484
rect 12333 -10520 12345 -10484
rect 12287 -10554 12345 -10520
rect 12287 -10590 12299 -10554
rect 12333 -10590 12345 -10554
rect 12287 -10625 12345 -10590
rect 12287 -10661 12299 -10625
rect 12333 -10661 12345 -10625
rect 12287 -10672 12345 -10661
rect 12545 -10484 12603 -10472
rect 12545 -10520 12557 -10484
rect 12591 -10520 12603 -10484
rect 12545 -10554 12603 -10520
rect 12545 -10590 12557 -10554
rect 12591 -10590 12603 -10554
rect 12545 -10624 12603 -10590
rect 12545 -10660 12557 -10624
rect 12591 -10660 12603 -10624
rect 12545 -10672 12603 -10660
rect 12803 -10484 12861 -10472
rect 12803 -10520 12815 -10484
rect 12849 -10520 12861 -10484
rect 12803 -10554 12861 -10520
rect 12803 -10590 12815 -10554
rect 12849 -10590 12861 -10554
rect 12803 -10624 12861 -10590
rect 12803 -10660 12815 -10624
rect 12849 -10660 12861 -10624
rect 12803 -10672 12861 -10660
rect 13061 -10484 13119 -10472
rect 13061 -10520 13073 -10484
rect 13107 -10520 13119 -10484
rect 13061 -10554 13119 -10520
rect 13061 -10590 13073 -10554
rect 13107 -10590 13119 -10554
rect 13061 -10624 13119 -10590
rect 13061 -10660 13073 -10624
rect 13107 -10660 13119 -10624
rect 13061 -10672 13119 -10660
rect 13319 -10484 13377 -10472
rect 13319 -10520 13331 -10484
rect 13365 -10520 13377 -10484
rect 13319 -10554 13377 -10520
rect 13319 -10590 13331 -10554
rect 13365 -10590 13377 -10554
rect 13319 -10624 13377 -10590
rect 13319 -10660 13331 -10624
rect 13365 -10660 13377 -10624
rect 13319 -10672 13377 -10660
rect 13577 -10484 13635 -10472
rect 13577 -10520 13589 -10484
rect 13623 -10520 13635 -10484
rect 13577 -10554 13635 -10520
rect 13577 -10590 13589 -10554
rect 13623 -10590 13635 -10554
rect 13577 -10624 13635 -10590
rect 13577 -10660 13589 -10624
rect 13623 -10660 13635 -10624
rect 13577 -10672 13635 -10660
rect 13835 -10484 13893 -10472
rect 13835 -10520 13847 -10484
rect 13881 -10520 13893 -10484
rect 13835 -10554 13893 -10520
rect 13835 -10590 13847 -10554
rect 13881 -10590 13893 -10554
rect 13835 -10624 13893 -10590
rect 13835 -10660 13847 -10624
rect 13881 -10660 13893 -10624
rect 13835 -10672 13893 -10660
rect 14434 -10483 14492 -10471
rect 14434 -10519 14446 -10483
rect 14480 -10519 14492 -10483
rect 14434 -10553 14492 -10519
rect 14434 -10589 14446 -10553
rect 14480 -10589 14492 -10553
rect 14434 -10623 14492 -10589
rect 14434 -10659 14446 -10623
rect 14480 -10659 14492 -10623
rect 14434 -10671 14492 -10659
rect 14692 -10483 14750 -10471
rect 14692 -10519 14704 -10483
rect 14738 -10519 14750 -10483
rect 14692 -10553 14750 -10519
rect 14692 -10589 14704 -10553
rect 14738 -10589 14750 -10553
rect 14692 -10623 14750 -10589
rect 14692 -10659 14704 -10623
rect 14738 -10659 14750 -10623
rect 14692 -10671 14750 -10659
rect 14950 -10483 15008 -10471
rect 14950 -10519 14962 -10483
rect 14996 -10519 15008 -10483
rect 14950 -10553 15008 -10519
rect 14950 -10589 14962 -10553
rect 14996 -10589 15008 -10553
rect 14950 -10624 15008 -10589
rect 14950 -10660 14962 -10624
rect 14996 -10660 15008 -10624
rect 14950 -10671 15008 -10660
rect 15208 -10483 15266 -10471
rect 15208 -10519 15220 -10483
rect 15254 -10519 15266 -10483
rect 15208 -10553 15266 -10519
rect 15208 -10589 15220 -10553
rect 15254 -10589 15266 -10553
rect 15208 -10623 15266 -10589
rect 15208 -10659 15220 -10623
rect 15254 -10659 15266 -10623
rect 15208 -10671 15266 -10659
rect 15466 -10483 15524 -10471
rect 15466 -10519 15478 -10483
rect 15512 -10519 15524 -10483
rect 15466 -10553 15524 -10519
rect 15466 -10589 15478 -10553
rect 15512 -10589 15524 -10553
rect 15466 -10623 15524 -10589
rect 15466 -10659 15478 -10623
rect 15512 -10659 15524 -10623
rect 15466 -10671 15524 -10659
rect 15724 -10483 15782 -10471
rect 15724 -10519 15736 -10483
rect 15770 -10519 15782 -10483
rect 15724 -10553 15782 -10519
rect 15724 -10589 15736 -10553
rect 15770 -10589 15782 -10553
rect 15724 -10623 15782 -10589
rect 15724 -10659 15736 -10623
rect 15770 -10659 15782 -10623
rect 15724 -10671 15782 -10659
rect 15982 -10483 16040 -10471
rect 15982 -10519 15994 -10483
rect 16028 -10519 16040 -10483
rect 15982 -10553 16040 -10519
rect 15982 -10589 15994 -10553
rect 16028 -10589 16040 -10553
rect 15982 -10623 16040 -10589
rect 15982 -10659 15994 -10623
rect 16028 -10659 16040 -10623
rect 15982 -10671 16040 -10659
rect 16240 -10483 16298 -10471
rect 16240 -10519 16252 -10483
rect 16286 -10519 16298 -10483
rect 16240 -10553 16298 -10519
rect 16240 -10589 16252 -10553
rect 16286 -10589 16298 -10553
rect 16240 -10623 16298 -10589
rect 16240 -10659 16252 -10623
rect 16286 -10659 16298 -10623
rect 16240 -10671 16298 -10659
rect 16498 -10483 16556 -10471
rect 16498 -10519 16510 -10483
rect 16544 -10519 16556 -10483
rect 16498 -10553 16556 -10519
rect 16498 -10589 16510 -10553
rect 16544 -10589 16556 -10553
rect 16498 -10623 16556 -10589
rect 16498 -10659 16510 -10623
rect 16544 -10659 16556 -10623
rect 16498 -10671 16556 -10659
rect 9101 -10902 9159 -10890
rect 9101 -10938 9113 -10902
rect 9147 -10938 9159 -10902
rect 9101 -10972 9159 -10938
rect 9101 -11008 9113 -10972
rect 9147 -11008 9159 -10972
rect 9101 -11042 9159 -11008
rect 9101 -11078 9113 -11042
rect 9147 -11078 9159 -11042
rect 9101 -11090 9159 -11078
rect 9359 -10902 9417 -10890
rect 9359 -10938 9371 -10902
rect 9405 -10938 9417 -10902
rect 9359 -10972 9417 -10938
rect 9359 -11008 9371 -10972
rect 9405 -11008 9417 -10972
rect 9359 -11042 9417 -11008
rect 9359 -11078 9371 -11042
rect 9405 -11078 9417 -11042
rect 9359 -11090 9417 -11078
rect 9617 -10902 9675 -10890
rect 9617 -10938 9629 -10902
rect 9663 -10938 9675 -10902
rect 9617 -10972 9675 -10938
rect 9617 -11008 9629 -10972
rect 9663 -11008 9675 -10972
rect 9617 -11043 9675 -11008
rect 9617 -11079 9629 -11043
rect 9663 -11079 9675 -11043
rect 9617 -11090 9675 -11079
rect 9875 -10902 9933 -10890
rect 9875 -10938 9887 -10902
rect 9921 -10938 9933 -10902
rect 9875 -10972 9933 -10938
rect 9875 -11008 9887 -10972
rect 9921 -11008 9933 -10972
rect 9875 -11042 9933 -11008
rect 9875 -11078 9887 -11042
rect 9921 -11078 9933 -11042
rect 9875 -11090 9933 -11078
rect 10133 -10902 10191 -10890
rect 10133 -10938 10145 -10902
rect 10179 -10938 10191 -10902
rect 10133 -10972 10191 -10938
rect 10133 -11008 10145 -10972
rect 10179 -11008 10191 -10972
rect 10133 -11042 10191 -11008
rect 10133 -11078 10145 -11042
rect 10179 -11078 10191 -11042
rect 10133 -11090 10191 -11078
rect 10391 -10902 10449 -10890
rect 10391 -10938 10403 -10902
rect 10437 -10938 10449 -10902
rect 10391 -10972 10449 -10938
rect 10391 -11008 10403 -10972
rect 10437 -11008 10449 -10972
rect 10391 -11042 10449 -11008
rect 10391 -11078 10403 -11042
rect 10437 -11078 10449 -11042
rect 10391 -11090 10449 -11078
rect 10649 -10902 10707 -10890
rect 10649 -10938 10661 -10902
rect 10695 -10938 10707 -10902
rect 10649 -10972 10707 -10938
rect 10649 -11008 10661 -10972
rect 10695 -11008 10707 -10972
rect 10649 -11042 10707 -11008
rect 10649 -11078 10661 -11042
rect 10695 -11078 10707 -11042
rect 10649 -11090 10707 -11078
rect 10907 -10902 10965 -10890
rect 10907 -10938 10919 -10902
rect 10953 -10938 10965 -10902
rect 10907 -10972 10965 -10938
rect 10907 -11008 10919 -10972
rect 10953 -11008 10965 -10972
rect 10907 -11042 10965 -11008
rect 10907 -11078 10919 -11042
rect 10953 -11078 10965 -11042
rect 10907 -11090 10965 -11078
rect 11165 -10902 11223 -10890
rect 11165 -10938 11177 -10902
rect 11211 -10938 11223 -10902
rect 11165 -10972 11223 -10938
rect 11165 -11008 11177 -10972
rect 11211 -11008 11223 -10972
rect 11165 -11042 11223 -11008
rect 11165 -11078 11177 -11042
rect 11211 -11078 11223 -11042
rect 11165 -11090 11223 -11078
rect 11771 -10902 11829 -10890
rect 11771 -10938 11783 -10902
rect 11817 -10938 11829 -10902
rect 11771 -10972 11829 -10938
rect 11771 -11008 11783 -10972
rect 11817 -11008 11829 -10972
rect 11771 -11042 11829 -11008
rect 11771 -11078 11783 -11042
rect 11817 -11078 11829 -11042
rect 11771 -11090 11829 -11078
rect 12029 -10902 12087 -10890
rect 12029 -10938 12041 -10902
rect 12075 -10938 12087 -10902
rect 12029 -10972 12087 -10938
rect 12029 -11008 12041 -10972
rect 12075 -11008 12087 -10972
rect 12029 -11042 12087 -11008
rect 12029 -11078 12041 -11042
rect 12075 -11078 12087 -11042
rect 12029 -11090 12087 -11078
rect 12287 -10902 12345 -10890
rect 12287 -10938 12299 -10902
rect 12333 -10938 12345 -10902
rect 12287 -10972 12345 -10938
rect 12287 -11008 12299 -10972
rect 12333 -11008 12345 -10972
rect 12287 -11043 12345 -11008
rect 12287 -11079 12299 -11043
rect 12333 -11079 12345 -11043
rect 12287 -11090 12345 -11079
rect 12545 -10902 12603 -10890
rect 12545 -10938 12557 -10902
rect 12591 -10938 12603 -10902
rect 12545 -10972 12603 -10938
rect 12545 -11008 12557 -10972
rect 12591 -11008 12603 -10972
rect 12545 -11042 12603 -11008
rect 12545 -11078 12557 -11042
rect 12591 -11078 12603 -11042
rect 12545 -11090 12603 -11078
rect 12803 -10902 12861 -10890
rect 12803 -10938 12815 -10902
rect 12849 -10938 12861 -10902
rect 12803 -10972 12861 -10938
rect 12803 -11008 12815 -10972
rect 12849 -11008 12861 -10972
rect 12803 -11042 12861 -11008
rect 12803 -11078 12815 -11042
rect 12849 -11078 12861 -11042
rect 12803 -11090 12861 -11078
rect 13061 -10902 13119 -10890
rect 13061 -10938 13073 -10902
rect 13107 -10938 13119 -10902
rect 13061 -10972 13119 -10938
rect 13061 -11008 13073 -10972
rect 13107 -11008 13119 -10972
rect 13061 -11042 13119 -11008
rect 13061 -11078 13073 -11042
rect 13107 -11078 13119 -11042
rect 13061 -11090 13119 -11078
rect 13319 -10902 13377 -10890
rect 13319 -10938 13331 -10902
rect 13365 -10938 13377 -10902
rect 13319 -10972 13377 -10938
rect 13319 -11008 13331 -10972
rect 13365 -11008 13377 -10972
rect 13319 -11042 13377 -11008
rect 13319 -11078 13331 -11042
rect 13365 -11078 13377 -11042
rect 13319 -11090 13377 -11078
rect 13577 -10902 13635 -10890
rect 13577 -10938 13589 -10902
rect 13623 -10938 13635 -10902
rect 13577 -10972 13635 -10938
rect 13577 -11008 13589 -10972
rect 13623 -11008 13635 -10972
rect 13577 -11042 13635 -11008
rect 13577 -11078 13589 -11042
rect 13623 -11078 13635 -11042
rect 13577 -11090 13635 -11078
rect 13835 -10902 13893 -10890
rect 13835 -10938 13847 -10902
rect 13881 -10938 13893 -10902
rect 13835 -10972 13893 -10938
rect 13835 -11008 13847 -10972
rect 13881 -11008 13893 -10972
rect 13835 -11042 13893 -11008
rect 13835 -11078 13847 -11042
rect 13881 -11078 13893 -11042
rect 13835 -11090 13893 -11078
rect 14434 -10901 14492 -10889
rect 14434 -10937 14446 -10901
rect 14480 -10937 14492 -10901
rect 14434 -10971 14492 -10937
rect 14434 -11007 14446 -10971
rect 14480 -11007 14492 -10971
rect 14434 -11041 14492 -11007
rect 14434 -11077 14446 -11041
rect 14480 -11077 14492 -11041
rect 14434 -11089 14492 -11077
rect 14692 -10901 14750 -10889
rect 14692 -10937 14704 -10901
rect 14738 -10937 14750 -10901
rect 14692 -10971 14750 -10937
rect 14692 -11007 14704 -10971
rect 14738 -11007 14750 -10971
rect 14692 -11041 14750 -11007
rect 14692 -11077 14704 -11041
rect 14738 -11077 14750 -11041
rect 14692 -11089 14750 -11077
rect 14950 -10901 15008 -10889
rect 14950 -10937 14962 -10901
rect 14996 -10937 15008 -10901
rect 14950 -10971 15008 -10937
rect 14950 -11007 14962 -10971
rect 14996 -11007 15008 -10971
rect 14950 -11042 15008 -11007
rect 14950 -11078 14962 -11042
rect 14996 -11078 15008 -11042
rect 14950 -11089 15008 -11078
rect 15208 -10901 15266 -10889
rect 15208 -10937 15220 -10901
rect 15254 -10937 15266 -10901
rect 15208 -10971 15266 -10937
rect 15208 -11007 15220 -10971
rect 15254 -11007 15266 -10971
rect 15208 -11041 15266 -11007
rect 15208 -11077 15220 -11041
rect 15254 -11077 15266 -11041
rect 15208 -11089 15266 -11077
rect 15466 -10901 15524 -10889
rect 15466 -10937 15478 -10901
rect 15512 -10937 15524 -10901
rect 15466 -10971 15524 -10937
rect 15466 -11007 15478 -10971
rect 15512 -11007 15524 -10971
rect 15466 -11041 15524 -11007
rect 15466 -11077 15478 -11041
rect 15512 -11077 15524 -11041
rect 15466 -11089 15524 -11077
rect 15724 -10901 15782 -10889
rect 15724 -10937 15736 -10901
rect 15770 -10937 15782 -10901
rect 15724 -10971 15782 -10937
rect 15724 -11007 15736 -10971
rect 15770 -11007 15782 -10971
rect 15724 -11041 15782 -11007
rect 15724 -11077 15736 -11041
rect 15770 -11077 15782 -11041
rect 15724 -11089 15782 -11077
rect 15982 -10901 16040 -10889
rect 15982 -10937 15994 -10901
rect 16028 -10937 16040 -10901
rect 15982 -10971 16040 -10937
rect 15982 -11007 15994 -10971
rect 16028 -11007 16040 -10971
rect 15982 -11041 16040 -11007
rect 15982 -11077 15994 -11041
rect 16028 -11077 16040 -11041
rect 15982 -11089 16040 -11077
rect 16240 -10901 16298 -10889
rect 16240 -10937 16252 -10901
rect 16286 -10937 16298 -10901
rect 16240 -10971 16298 -10937
rect 16240 -11007 16252 -10971
rect 16286 -11007 16298 -10971
rect 16240 -11041 16298 -11007
rect 16240 -11077 16252 -11041
rect 16286 -11077 16298 -11041
rect 16240 -11089 16298 -11077
rect 16498 -10901 16556 -10889
rect 16498 -10937 16510 -10901
rect 16544 -10937 16556 -10901
rect 16498 -10971 16556 -10937
rect 16498 -11007 16510 -10971
rect 16544 -11007 16556 -10971
rect 16498 -11041 16556 -11007
rect 16498 -11077 16510 -11041
rect 16544 -11077 16556 -11041
rect 16498 -11089 16556 -11077
rect 9101 -11320 9159 -11308
rect 9101 -11356 9113 -11320
rect 9147 -11356 9159 -11320
rect 9101 -11390 9159 -11356
rect 9101 -11426 9113 -11390
rect 9147 -11426 9159 -11390
rect 9101 -11460 9159 -11426
rect 9101 -11496 9113 -11460
rect 9147 -11496 9159 -11460
rect 9101 -11508 9159 -11496
rect 9359 -11320 9417 -11308
rect 9359 -11356 9371 -11320
rect 9405 -11356 9417 -11320
rect 9359 -11390 9417 -11356
rect 9359 -11426 9371 -11390
rect 9405 -11426 9417 -11390
rect 9359 -11460 9417 -11426
rect 9359 -11496 9371 -11460
rect 9405 -11496 9417 -11460
rect 9359 -11508 9417 -11496
rect 9617 -11320 9675 -11308
rect 9617 -11356 9629 -11320
rect 9663 -11356 9675 -11320
rect 9617 -11390 9675 -11356
rect 9617 -11426 9629 -11390
rect 9663 -11426 9675 -11390
rect 9617 -11461 9675 -11426
rect 9617 -11497 9629 -11461
rect 9663 -11497 9675 -11461
rect 9617 -11508 9675 -11497
rect 9875 -11320 9933 -11308
rect 9875 -11356 9887 -11320
rect 9921 -11356 9933 -11320
rect 9875 -11390 9933 -11356
rect 9875 -11426 9887 -11390
rect 9921 -11426 9933 -11390
rect 9875 -11460 9933 -11426
rect 9875 -11496 9887 -11460
rect 9921 -11496 9933 -11460
rect 9875 -11508 9933 -11496
rect 10133 -11320 10191 -11308
rect 10133 -11356 10145 -11320
rect 10179 -11356 10191 -11320
rect 10133 -11390 10191 -11356
rect 10133 -11426 10145 -11390
rect 10179 -11426 10191 -11390
rect 10133 -11460 10191 -11426
rect 10133 -11496 10145 -11460
rect 10179 -11496 10191 -11460
rect 10133 -11508 10191 -11496
rect 10391 -11320 10449 -11308
rect 10391 -11356 10403 -11320
rect 10437 -11356 10449 -11320
rect 10391 -11390 10449 -11356
rect 10391 -11426 10403 -11390
rect 10437 -11426 10449 -11390
rect 10391 -11460 10449 -11426
rect 10391 -11496 10403 -11460
rect 10437 -11496 10449 -11460
rect 10391 -11508 10449 -11496
rect 10649 -11320 10707 -11308
rect 10649 -11356 10661 -11320
rect 10695 -11356 10707 -11320
rect 10649 -11390 10707 -11356
rect 10649 -11426 10661 -11390
rect 10695 -11426 10707 -11390
rect 10649 -11460 10707 -11426
rect 10649 -11496 10661 -11460
rect 10695 -11496 10707 -11460
rect 10649 -11508 10707 -11496
rect 10907 -11320 10965 -11308
rect 10907 -11356 10919 -11320
rect 10953 -11356 10965 -11320
rect 10907 -11390 10965 -11356
rect 10907 -11426 10919 -11390
rect 10953 -11426 10965 -11390
rect 10907 -11460 10965 -11426
rect 10907 -11496 10919 -11460
rect 10953 -11496 10965 -11460
rect 10907 -11508 10965 -11496
rect 11165 -11320 11223 -11308
rect 11165 -11356 11177 -11320
rect 11211 -11356 11223 -11320
rect 11165 -11390 11223 -11356
rect 11165 -11426 11177 -11390
rect 11211 -11426 11223 -11390
rect 11165 -11460 11223 -11426
rect 11165 -11496 11177 -11460
rect 11211 -11496 11223 -11460
rect 11165 -11508 11223 -11496
rect 11771 -11320 11829 -11308
rect 11771 -11356 11783 -11320
rect 11817 -11356 11829 -11320
rect 11771 -11390 11829 -11356
rect 11771 -11426 11783 -11390
rect 11817 -11426 11829 -11390
rect 11771 -11460 11829 -11426
rect 11771 -11496 11783 -11460
rect 11817 -11496 11829 -11460
rect 11771 -11508 11829 -11496
rect 12029 -11320 12087 -11308
rect 12029 -11356 12041 -11320
rect 12075 -11356 12087 -11320
rect 12029 -11390 12087 -11356
rect 12029 -11426 12041 -11390
rect 12075 -11426 12087 -11390
rect 12029 -11460 12087 -11426
rect 12029 -11496 12041 -11460
rect 12075 -11496 12087 -11460
rect 12029 -11508 12087 -11496
rect 12287 -11320 12345 -11308
rect 12287 -11356 12299 -11320
rect 12333 -11356 12345 -11320
rect 12287 -11390 12345 -11356
rect 12287 -11426 12299 -11390
rect 12333 -11426 12345 -11390
rect 12287 -11461 12345 -11426
rect 12287 -11497 12299 -11461
rect 12333 -11497 12345 -11461
rect 12287 -11508 12345 -11497
rect 12545 -11320 12603 -11308
rect 12545 -11356 12557 -11320
rect 12591 -11356 12603 -11320
rect 12545 -11390 12603 -11356
rect 12545 -11426 12557 -11390
rect 12591 -11426 12603 -11390
rect 12545 -11460 12603 -11426
rect 12545 -11496 12557 -11460
rect 12591 -11496 12603 -11460
rect 12545 -11508 12603 -11496
rect 12803 -11320 12861 -11308
rect 12803 -11356 12815 -11320
rect 12849 -11356 12861 -11320
rect 12803 -11390 12861 -11356
rect 12803 -11426 12815 -11390
rect 12849 -11426 12861 -11390
rect 12803 -11460 12861 -11426
rect 12803 -11496 12815 -11460
rect 12849 -11496 12861 -11460
rect 12803 -11508 12861 -11496
rect 13061 -11320 13119 -11308
rect 13061 -11356 13073 -11320
rect 13107 -11356 13119 -11320
rect 13061 -11390 13119 -11356
rect 13061 -11426 13073 -11390
rect 13107 -11426 13119 -11390
rect 13061 -11460 13119 -11426
rect 13061 -11496 13073 -11460
rect 13107 -11496 13119 -11460
rect 13061 -11508 13119 -11496
rect 13319 -11320 13377 -11308
rect 13319 -11356 13331 -11320
rect 13365 -11356 13377 -11320
rect 13319 -11390 13377 -11356
rect 13319 -11426 13331 -11390
rect 13365 -11426 13377 -11390
rect 13319 -11460 13377 -11426
rect 13319 -11496 13331 -11460
rect 13365 -11496 13377 -11460
rect 13319 -11508 13377 -11496
rect 13577 -11320 13635 -11308
rect 13577 -11356 13589 -11320
rect 13623 -11356 13635 -11320
rect 13577 -11390 13635 -11356
rect 13577 -11426 13589 -11390
rect 13623 -11426 13635 -11390
rect 13577 -11460 13635 -11426
rect 13577 -11496 13589 -11460
rect 13623 -11496 13635 -11460
rect 13577 -11508 13635 -11496
rect 13835 -11320 13893 -11308
rect 13835 -11356 13847 -11320
rect 13881 -11356 13893 -11320
rect 13835 -11390 13893 -11356
rect 13835 -11426 13847 -11390
rect 13881 -11426 13893 -11390
rect 13835 -11460 13893 -11426
rect 13835 -11496 13847 -11460
rect 13881 -11496 13893 -11460
rect 13835 -11508 13893 -11496
rect 14434 -11319 14492 -11307
rect 14434 -11355 14446 -11319
rect 14480 -11355 14492 -11319
rect 14434 -11389 14492 -11355
rect 14434 -11425 14446 -11389
rect 14480 -11425 14492 -11389
rect 14434 -11459 14492 -11425
rect 14434 -11495 14446 -11459
rect 14480 -11495 14492 -11459
rect 14434 -11507 14492 -11495
rect 14692 -11319 14750 -11307
rect 14692 -11355 14704 -11319
rect 14738 -11355 14750 -11319
rect 14692 -11389 14750 -11355
rect 14692 -11425 14704 -11389
rect 14738 -11425 14750 -11389
rect 14692 -11459 14750 -11425
rect 14692 -11495 14704 -11459
rect 14738 -11495 14750 -11459
rect 14692 -11507 14750 -11495
rect 14950 -11319 15008 -11307
rect 14950 -11355 14962 -11319
rect 14996 -11355 15008 -11319
rect 14950 -11389 15008 -11355
rect 14950 -11425 14962 -11389
rect 14996 -11425 15008 -11389
rect 14950 -11460 15008 -11425
rect 14950 -11496 14962 -11460
rect 14996 -11496 15008 -11460
rect 14950 -11507 15008 -11496
rect 15208 -11319 15266 -11307
rect 15208 -11355 15220 -11319
rect 15254 -11355 15266 -11319
rect 15208 -11389 15266 -11355
rect 15208 -11425 15220 -11389
rect 15254 -11425 15266 -11389
rect 15208 -11459 15266 -11425
rect 15208 -11495 15220 -11459
rect 15254 -11495 15266 -11459
rect 15208 -11507 15266 -11495
rect 15466 -11319 15524 -11307
rect 15466 -11355 15478 -11319
rect 15512 -11355 15524 -11319
rect 15466 -11389 15524 -11355
rect 15466 -11425 15478 -11389
rect 15512 -11425 15524 -11389
rect 15466 -11459 15524 -11425
rect 15466 -11495 15478 -11459
rect 15512 -11495 15524 -11459
rect 15466 -11507 15524 -11495
rect 15724 -11319 15782 -11307
rect 15724 -11355 15736 -11319
rect 15770 -11355 15782 -11319
rect 15724 -11389 15782 -11355
rect 15724 -11425 15736 -11389
rect 15770 -11425 15782 -11389
rect 15724 -11459 15782 -11425
rect 15724 -11495 15736 -11459
rect 15770 -11495 15782 -11459
rect 15724 -11507 15782 -11495
rect 15982 -11319 16040 -11307
rect 15982 -11355 15994 -11319
rect 16028 -11355 16040 -11319
rect 15982 -11389 16040 -11355
rect 15982 -11425 15994 -11389
rect 16028 -11425 16040 -11389
rect 15982 -11459 16040 -11425
rect 15982 -11495 15994 -11459
rect 16028 -11495 16040 -11459
rect 15982 -11507 16040 -11495
rect 16240 -11319 16298 -11307
rect 16240 -11355 16252 -11319
rect 16286 -11355 16298 -11319
rect 16240 -11389 16298 -11355
rect 16240 -11425 16252 -11389
rect 16286 -11425 16298 -11389
rect 16240 -11459 16298 -11425
rect 16240 -11495 16252 -11459
rect 16286 -11495 16298 -11459
rect 16240 -11507 16298 -11495
rect 16498 -11319 16556 -11307
rect 16498 -11355 16510 -11319
rect 16544 -11355 16556 -11319
rect 16498 -11389 16556 -11355
rect 16498 -11425 16510 -11389
rect 16544 -11425 16556 -11389
rect 16498 -11459 16556 -11425
rect 16498 -11495 16510 -11459
rect 16544 -11495 16556 -11459
rect 16498 -11507 16556 -11495
rect 9101 -11738 9159 -11726
rect 9101 -11774 9113 -11738
rect 9147 -11774 9159 -11738
rect 9101 -11808 9159 -11774
rect 9101 -11844 9113 -11808
rect 9147 -11844 9159 -11808
rect 9101 -11878 9159 -11844
rect 9101 -11914 9113 -11878
rect 9147 -11914 9159 -11878
rect 9101 -11926 9159 -11914
rect 9359 -11738 9417 -11726
rect 9359 -11774 9371 -11738
rect 9405 -11774 9417 -11738
rect 9359 -11808 9417 -11774
rect 9359 -11844 9371 -11808
rect 9405 -11844 9417 -11808
rect 9359 -11878 9417 -11844
rect 9359 -11914 9371 -11878
rect 9405 -11914 9417 -11878
rect 9359 -11926 9417 -11914
rect 9617 -11738 9675 -11726
rect 9617 -11774 9629 -11738
rect 9663 -11774 9675 -11738
rect 9617 -11808 9675 -11774
rect 9617 -11844 9629 -11808
rect 9663 -11844 9675 -11808
rect 9617 -11879 9675 -11844
rect 9617 -11915 9629 -11879
rect 9663 -11915 9675 -11879
rect 9617 -11926 9675 -11915
rect 9875 -11738 9933 -11726
rect 9875 -11774 9887 -11738
rect 9921 -11774 9933 -11738
rect 9875 -11808 9933 -11774
rect 9875 -11844 9887 -11808
rect 9921 -11844 9933 -11808
rect 9875 -11878 9933 -11844
rect 9875 -11914 9887 -11878
rect 9921 -11914 9933 -11878
rect 9875 -11926 9933 -11914
rect 10133 -11738 10191 -11726
rect 10133 -11774 10145 -11738
rect 10179 -11774 10191 -11738
rect 10133 -11808 10191 -11774
rect 10133 -11844 10145 -11808
rect 10179 -11844 10191 -11808
rect 10133 -11878 10191 -11844
rect 10133 -11914 10145 -11878
rect 10179 -11914 10191 -11878
rect 10133 -11926 10191 -11914
rect 10391 -11738 10449 -11726
rect 10391 -11774 10403 -11738
rect 10437 -11774 10449 -11738
rect 10391 -11808 10449 -11774
rect 10391 -11844 10403 -11808
rect 10437 -11844 10449 -11808
rect 10391 -11878 10449 -11844
rect 10391 -11914 10403 -11878
rect 10437 -11914 10449 -11878
rect 10391 -11926 10449 -11914
rect 10649 -11738 10707 -11726
rect 10649 -11774 10661 -11738
rect 10695 -11774 10707 -11738
rect 10649 -11808 10707 -11774
rect 10649 -11844 10661 -11808
rect 10695 -11844 10707 -11808
rect 10649 -11878 10707 -11844
rect 10649 -11914 10661 -11878
rect 10695 -11914 10707 -11878
rect 10649 -11926 10707 -11914
rect 10907 -11738 10965 -11726
rect 10907 -11774 10919 -11738
rect 10953 -11774 10965 -11738
rect 10907 -11808 10965 -11774
rect 10907 -11844 10919 -11808
rect 10953 -11844 10965 -11808
rect 10907 -11878 10965 -11844
rect 10907 -11914 10919 -11878
rect 10953 -11914 10965 -11878
rect 10907 -11926 10965 -11914
rect 11165 -11738 11223 -11726
rect 11165 -11774 11177 -11738
rect 11211 -11774 11223 -11738
rect 11165 -11808 11223 -11774
rect 11165 -11844 11177 -11808
rect 11211 -11844 11223 -11808
rect 11165 -11878 11223 -11844
rect 11165 -11914 11177 -11878
rect 11211 -11914 11223 -11878
rect 11165 -11926 11223 -11914
rect 11771 -11738 11829 -11726
rect 11771 -11774 11783 -11738
rect 11817 -11774 11829 -11738
rect 11771 -11808 11829 -11774
rect 11771 -11844 11783 -11808
rect 11817 -11844 11829 -11808
rect 11771 -11878 11829 -11844
rect 11771 -11914 11783 -11878
rect 11817 -11914 11829 -11878
rect 11771 -11926 11829 -11914
rect 12029 -11738 12087 -11726
rect 12029 -11774 12041 -11738
rect 12075 -11774 12087 -11738
rect 12029 -11808 12087 -11774
rect 12029 -11844 12041 -11808
rect 12075 -11844 12087 -11808
rect 12029 -11878 12087 -11844
rect 12029 -11914 12041 -11878
rect 12075 -11914 12087 -11878
rect 12029 -11926 12087 -11914
rect 12287 -11738 12345 -11726
rect 12287 -11774 12299 -11738
rect 12333 -11774 12345 -11738
rect 12287 -11808 12345 -11774
rect 12287 -11844 12299 -11808
rect 12333 -11844 12345 -11808
rect 12287 -11879 12345 -11844
rect 12287 -11915 12299 -11879
rect 12333 -11915 12345 -11879
rect 12287 -11926 12345 -11915
rect 12545 -11738 12603 -11726
rect 12545 -11774 12557 -11738
rect 12591 -11774 12603 -11738
rect 12545 -11808 12603 -11774
rect 12545 -11844 12557 -11808
rect 12591 -11844 12603 -11808
rect 12545 -11878 12603 -11844
rect 12545 -11914 12557 -11878
rect 12591 -11914 12603 -11878
rect 12545 -11926 12603 -11914
rect 12803 -11738 12861 -11726
rect 12803 -11774 12815 -11738
rect 12849 -11774 12861 -11738
rect 12803 -11808 12861 -11774
rect 12803 -11844 12815 -11808
rect 12849 -11844 12861 -11808
rect 12803 -11878 12861 -11844
rect 12803 -11914 12815 -11878
rect 12849 -11914 12861 -11878
rect 12803 -11926 12861 -11914
rect 13061 -11738 13119 -11726
rect 13061 -11774 13073 -11738
rect 13107 -11774 13119 -11738
rect 13061 -11808 13119 -11774
rect 13061 -11844 13073 -11808
rect 13107 -11844 13119 -11808
rect 13061 -11878 13119 -11844
rect 13061 -11914 13073 -11878
rect 13107 -11914 13119 -11878
rect 13061 -11926 13119 -11914
rect 13319 -11738 13377 -11726
rect 13319 -11774 13331 -11738
rect 13365 -11774 13377 -11738
rect 13319 -11808 13377 -11774
rect 13319 -11844 13331 -11808
rect 13365 -11844 13377 -11808
rect 13319 -11878 13377 -11844
rect 13319 -11914 13331 -11878
rect 13365 -11914 13377 -11878
rect 13319 -11926 13377 -11914
rect 13577 -11738 13635 -11726
rect 13577 -11774 13589 -11738
rect 13623 -11774 13635 -11738
rect 13577 -11808 13635 -11774
rect 13577 -11844 13589 -11808
rect 13623 -11844 13635 -11808
rect 13577 -11878 13635 -11844
rect 13577 -11914 13589 -11878
rect 13623 -11914 13635 -11878
rect 13577 -11926 13635 -11914
rect 13835 -11738 13893 -11726
rect 13835 -11774 13847 -11738
rect 13881 -11774 13893 -11738
rect 13835 -11808 13893 -11774
rect 13835 -11844 13847 -11808
rect 13881 -11844 13893 -11808
rect 13835 -11878 13893 -11844
rect 13835 -11914 13847 -11878
rect 13881 -11914 13893 -11878
rect 13835 -11926 13893 -11914
rect 14434 -11737 14492 -11725
rect 14434 -11773 14446 -11737
rect 14480 -11773 14492 -11737
rect 14434 -11807 14492 -11773
rect 14434 -11843 14446 -11807
rect 14480 -11843 14492 -11807
rect 14434 -11877 14492 -11843
rect 14434 -11913 14446 -11877
rect 14480 -11913 14492 -11877
rect 14434 -11925 14492 -11913
rect 14692 -11737 14750 -11725
rect 14692 -11773 14704 -11737
rect 14738 -11773 14750 -11737
rect 14692 -11807 14750 -11773
rect 14692 -11843 14704 -11807
rect 14738 -11843 14750 -11807
rect 14692 -11877 14750 -11843
rect 14692 -11913 14704 -11877
rect 14738 -11913 14750 -11877
rect 14692 -11925 14750 -11913
rect 14950 -11737 15008 -11725
rect 14950 -11773 14962 -11737
rect 14996 -11773 15008 -11737
rect 14950 -11807 15008 -11773
rect 14950 -11843 14962 -11807
rect 14996 -11843 15008 -11807
rect 14950 -11878 15008 -11843
rect 14950 -11914 14962 -11878
rect 14996 -11914 15008 -11878
rect 14950 -11925 15008 -11914
rect 15208 -11737 15266 -11725
rect 15208 -11773 15220 -11737
rect 15254 -11773 15266 -11737
rect 15208 -11807 15266 -11773
rect 15208 -11843 15220 -11807
rect 15254 -11843 15266 -11807
rect 15208 -11877 15266 -11843
rect 15208 -11913 15220 -11877
rect 15254 -11913 15266 -11877
rect 15208 -11925 15266 -11913
rect 15466 -11737 15524 -11725
rect 15466 -11773 15478 -11737
rect 15512 -11773 15524 -11737
rect 15466 -11807 15524 -11773
rect 15466 -11843 15478 -11807
rect 15512 -11843 15524 -11807
rect 15466 -11877 15524 -11843
rect 15466 -11913 15478 -11877
rect 15512 -11913 15524 -11877
rect 15466 -11925 15524 -11913
rect 15724 -11737 15782 -11725
rect 15724 -11773 15736 -11737
rect 15770 -11773 15782 -11737
rect 15724 -11807 15782 -11773
rect 15724 -11843 15736 -11807
rect 15770 -11843 15782 -11807
rect 15724 -11877 15782 -11843
rect 15724 -11913 15736 -11877
rect 15770 -11913 15782 -11877
rect 15724 -11925 15782 -11913
rect 15982 -11737 16040 -11725
rect 15982 -11773 15994 -11737
rect 16028 -11773 16040 -11737
rect 15982 -11807 16040 -11773
rect 15982 -11843 15994 -11807
rect 16028 -11843 16040 -11807
rect 15982 -11877 16040 -11843
rect 15982 -11913 15994 -11877
rect 16028 -11913 16040 -11877
rect 15982 -11925 16040 -11913
rect 16240 -11737 16298 -11725
rect 16240 -11773 16252 -11737
rect 16286 -11773 16298 -11737
rect 16240 -11807 16298 -11773
rect 16240 -11843 16252 -11807
rect 16286 -11843 16298 -11807
rect 16240 -11877 16298 -11843
rect 16240 -11913 16252 -11877
rect 16286 -11913 16298 -11877
rect 16240 -11925 16298 -11913
rect 16498 -11737 16556 -11725
rect 16498 -11773 16510 -11737
rect 16544 -11773 16556 -11737
rect 16498 -11807 16556 -11773
rect 16498 -11843 16510 -11807
rect 16544 -11843 16556 -11807
rect 16498 -11877 16556 -11843
rect 16498 -11913 16510 -11877
rect 16544 -11913 16556 -11877
rect 16498 -11925 16556 -11913
rect 9101 -12156 9159 -12144
rect 9101 -12192 9113 -12156
rect 9147 -12192 9159 -12156
rect 9101 -12226 9159 -12192
rect 9101 -12262 9113 -12226
rect 9147 -12262 9159 -12226
rect 9101 -12296 9159 -12262
rect 9101 -12332 9113 -12296
rect 9147 -12332 9159 -12296
rect 9101 -12344 9159 -12332
rect 9359 -12156 9417 -12144
rect 9359 -12192 9371 -12156
rect 9405 -12192 9417 -12156
rect 9359 -12226 9417 -12192
rect 9359 -12262 9371 -12226
rect 9405 -12262 9417 -12226
rect 9359 -12296 9417 -12262
rect 9359 -12332 9371 -12296
rect 9405 -12332 9417 -12296
rect 9359 -12344 9417 -12332
rect 9617 -12156 9675 -12144
rect 9617 -12192 9629 -12156
rect 9663 -12192 9675 -12156
rect 9617 -12226 9675 -12192
rect 9617 -12262 9629 -12226
rect 9663 -12262 9675 -12226
rect 9617 -12297 9675 -12262
rect 9617 -12333 9629 -12297
rect 9663 -12333 9675 -12297
rect 9617 -12344 9675 -12333
rect 9875 -12156 9933 -12144
rect 9875 -12192 9887 -12156
rect 9921 -12192 9933 -12156
rect 9875 -12226 9933 -12192
rect 9875 -12262 9887 -12226
rect 9921 -12262 9933 -12226
rect 9875 -12296 9933 -12262
rect 9875 -12332 9887 -12296
rect 9921 -12332 9933 -12296
rect 9875 -12344 9933 -12332
rect 10133 -12156 10191 -12144
rect 10133 -12192 10145 -12156
rect 10179 -12192 10191 -12156
rect 10133 -12226 10191 -12192
rect 10133 -12262 10145 -12226
rect 10179 -12262 10191 -12226
rect 10133 -12296 10191 -12262
rect 10133 -12332 10145 -12296
rect 10179 -12332 10191 -12296
rect 10133 -12344 10191 -12332
rect 10391 -12156 10449 -12144
rect 10391 -12192 10403 -12156
rect 10437 -12192 10449 -12156
rect 10391 -12226 10449 -12192
rect 10391 -12262 10403 -12226
rect 10437 -12262 10449 -12226
rect 10391 -12296 10449 -12262
rect 10391 -12332 10403 -12296
rect 10437 -12332 10449 -12296
rect 10391 -12344 10449 -12332
rect 10649 -12156 10707 -12144
rect 10649 -12192 10661 -12156
rect 10695 -12192 10707 -12156
rect 10649 -12226 10707 -12192
rect 10649 -12262 10661 -12226
rect 10695 -12262 10707 -12226
rect 10649 -12296 10707 -12262
rect 10649 -12332 10661 -12296
rect 10695 -12332 10707 -12296
rect 10649 -12344 10707 -12332
rect 10907 -12156 10965 -12144
rect 10907 -12192 10919 -12156
rect 10953 -12192 10965 -12156
rect 10907 -12226 10965 -12192
rect 10907 -12262 10919 -12226
rect 10953 -12262 10965 -12226
rect 10907 -12296 10965 -12262
rect 10907 -12332 10919 -12296
rect 10953 -12332 10965 -12296
rect 10907 -12344 10965 -12332
rect 11165 -12156 11223 -12144
rect 11165 -12192 11177 -12156
rect 11211 -12192 11223 -12156
rect 11165 -12226 11223 -12192
rect 11165 -12262 11177 -12226
rect 11211 -12262 11223 -12226
rect 11165 -12296 11223 -12262
rect 11165 -12332 11177 -12296
rect 11211 -12332 11223 -12296
rect 11165 -12344 11223 -12332
rect 11771 -12156 11829 -12144
rect 11771 -12192 11783 -12156
rect 11817 -12192 11829 -12156
rect 11771 -12226 11829 -12192
rect 11771 -12262 11783 -12226
rect 11817 -12262 11829 -12226
rect 11771 -12296 11829 -12262
rect 11771 -12332 11783 -12296
rect 11817 -12332 11829 -12296
rect 11771 -12344 11829 -12332
rect 12029 -12156 12087 -12144
rect 12029 -12192 12041 -12156
rect 12075 -12192 12087 -12156
rect 12029 -12226 12087 -12192
rect 12029 -12262 12041 -12226
rect 12075 -12262 12087 -12226
rect 12029 -12296 12087 -12262
rect 12029 -12332 12041 -12296
rect 12075 -12332 12087 -12296
rect 12029 -12344 12087 -12332
rect 12287 -12156 12345 -12144
rect 12287 -12192 12299 -12156
rect 12333 -12192 12345 -12156
rect 12287 -12226 12345 -12192
rect 12287 -12262 12299 -12226
rect 12333 -12262 12345 -12226
rect 12287 -12297 12345 -12262
rect 12287 -12333 12299 -12297
rect 12333 -12333 12345 -12297
rect 12287 -12344 12345 -12333
rect 12545 -12156 12603 -12144
rect 12545 -12192 12557 -12156
rect 12591 -12192 12603 -12156
rect 12545 -12226 12603 -12192
rect 12545 -12262 12557 -12226
rect 12591 -12262 12603 -12226
rect 12545 -12296 12603 -12262
rect 12545 -12332 12557 -12296
rect 12591 -12332 12603 -12296
rect 12545 -12344 12603 -12332
rect 12803 -12156 12861 -12144
rect 12803 -12192 12815 -12156
rect 12849 -12192 12861 -12156
rect 12803 -12226 12861 -12192
rect 12803 -12262 12815 -12226
rect 12849 -12262 12861 -12226
rect 12803 -12296 12861 -12262
rect 12803 -12332 12815 -12296
rect 12849 -12332 12861 -12296
rect 12803 -12344 12861 -12332
rect 13061 -12156 13119 -12144
rect 13061 -12192 13073 -12156
rect 13107 -12192 13119 -12156
rect 13061 -12226 13119 -12192
rect 13061 -12262 13073 -12226
rect 13107 -12262 13119 -12226
rect 13061 -12296 13119 -12262
rect 13061 -12332 13073 -12296
rect 13107 -12332 13119 -12296
rect 13061 -12344 13119 -12332
rect 13319 -12156 13377 -12144
rect 13319 -12192 13331 -12156
rect 13365 -12192 13377 -12156
rect 13319 -12226 13377 -12192
rect 13319 -12262 13331 -12226
rect 13365 -12262 13377 -12226
rect 13319 -12296 13377 -12262
rect 13319 -12332 13331 -12296
rect 13365 -12332 13377 -12296
rect 13319 -12344 13377 -12332
rect 13577 -12156 13635 -12144
rect 13577 -12192 13589 -12156
rect 13623 -12192 13635 -12156
rect 13577 -12226 13635 -12192
rect 13577 -12262 13589 -12226
rect 13623 -12262 13635 -12226
rect 13577 -12296 13635 -12262
rect 13577 -12332 13589 -12296
rect 13623 -12332 13635 -12296
rect 13577 -12344 13635 -12332
rect 13835 -12156 13893 -12144
rect 13835 -12192 13847 -12156
rect 13881 -12192 13893 -12156
rect 13835 -12226 13893 -12192
rect 13835 -12262 13847 -12226
rect 13881 -12262 13893 -12226
rect 13835 -12296 13893 -12262
rect 13835 -12332 13847 -12296
rect 13881 -12332 13893 -12296
rect 13835 -12344 13893 -12332
rect 14434 -12155 14492 -12143
rect 14434 -12191 14446 -12155
rect 14480 -12191 14492 -12155
rect 14434 -12225 14492 -12191
rect 14434 -12261 14446 -12225
rect 14480 -12261 14492 -12225
rect 14434 -12295 14492 -12261
rect 14434 -12331 14446 -12295
rect 14480 -12331 14492 -12295
rect 14434 -12343 14492 -12331
rect 14692 -12155 14750 -12143
rect 14692 -12191 14704 -12155
rect 14738 -12191 14750 -12155
rect 14692 -12225 14750 -12191
rect 14692 -12261 14704 -12225
rect 14738 -12261 14750 -12225
rect 14692 -12295 14750 -12261
rect 14692 -12331 14704 -12295
rect 14738 -12331 14750 -12295
rect 14692 -12343 14750 -12331
rect 14950 -12155 15008 -12143
rect 14950 -12191 14962 -12155
rect 14996 -12191 15008 -12155
rect 14950 -12225 15008 -12191
rect 14950 -12261 14962 -12225
rect 14996 -12261 15008 -12225
rect 14950 -12296 15008 -12261
rect 14950 -12332 14962 -12296
rect 14996 -12332 15008 -12296
rect 14950 -12343 15008 -12332
rect 15208 -12155 15266 -12143
rect 15208 -12191 15220 -12155
rect 15254 -12191 15266 -12155
rect 15208 -12225 15266 -12191
rect 15208 -12261 15220 -12225
rect 15254 -12261 15266 -12225
rect 15208 -12295 15266 -12261
rect 15208 -12331 15220 -12295
rect 15254 -12331 15266 -12295
rect 15208 -12343 15266 -12331
rect 15466 -12155 15524 -12143
rect 15466 -12191 15478 -12155
rect 15512 -12191 15524 -12155
rect 15466 -12225 15524 -12191
rect 15466 -12261 15478 -12225
rect 15512 -12261 15524 -12225
rect 15466 -12295 15524 -12261
rect 15466 -12331 15478 -12295
rect 15512 -12331 15524 -12295
rect 15466 -12343 15524 -12331
rect 15724 -12155 15782 -12143
rect 15724 -12191 15736 -12155
rect 15770 -12191 15782 -12155
rect 15724 -12225 15782 -12191
rect 15724 -12261 15736 -12225
rect 15770 -12261 15782 -12225
rect 15724 -12295 15782 -12261
rect 15724 -12331 15736 -12295
rect 15770 -12331 15782 -12295
rect 15724 -12343 15782 -12331
rect 15982 -12155 16040 -12143
rect 15982 -12191 15994 -12155
rect 16028 -12191 16040 -12155
rect 15982 -12225 16040 -12191
rect 15982 -12261 15994 -12225
rect 16028 -12261 16040 -12225
rect 15982 -12295 16040 -12261
rect 15982 -12331 15994 -12295
rect 16028 -12331 16040 -12295
rect 15982 -12343 16040 -12331
rect 16240 -12155 16298 -12143
rect 16240 -12191 16252 -12155
rect 16286 -12191 16298 -12155
rect 16240 -12225 16298 -12191
rect 16240 -12261 16252 -12225
rect 16286 -12261 16298 -12225
rect 16240 -12295 16298 -12261
rect 16240 -12331 16252 -12295
rect 16286 -12331 16298 -12295
rect 16240 -12343 16298 -12331
rect 16498 -12155 16556 -12143
rect 16498 -12191 16510 -12155
rect 16544 -12191 16556 -12155
rect 16498 -12225 16556 -12191
rect 16498 -12261 16510 -12225
rect 16544 -12261 16556 -12225
rect 16498 -12295 16556 -12261
rect 16498 -12331 16510 -12295
rect 16544 -12331 16556 -12295
rect 16498 -12343 16556 -12331
rect 8981 -12810 9039 -12796
rect 8981 -12844 8993 -12810
rect 9027 -12844 9039 -12810
rect 8981 -12878 9039 -12844
rect 8981 -12914 8993 -12878
rect 9027 -12914 9039 -12878
rect 8981 -12948 9039 -12914
rect 8981 -12982 8993 -12948
rect 9027 -12982 9039 -12948
rect 8981 -12996 9039 -12982
rect 9239 -12810 9297 -12796
rect 9239 -12844 9251 -12810
rect 9285 -12844 9297 -12810
rect 9239 -12878 9297 -12844
rect 9239 -12914 9251 -12878
rect 9285 -12914 9297 -12878
rect 9239 -12948 9297 -12914
rect 9239 -12982 9251 -12948
rect 9285 -12982 9297 -12948
rect 9239 -12996 9297 -12982
rect 9521 -12810 9579 -12796
rect 9521 -12844 9533 -12810
rect 9567 -12844 9579 -12810
rect 9521 -12878 9579 -12844
rect 9521 -12914 9533 -12878
rect 9567 -12914 9579 -12878
rect 9521 -12948 9579 -12914
rect 9521 -12982 9533 -12948
rect 9567 -12982 9579 -12948
rect 9521 -12996 9579 -12982
rect 9779 -12810 9837 -12796
rect 9779 -12844 9791 -12810
rect 9825 -12844 9837 -12810
rect 9779 -12878 9837 -12844
rect 9779 -12914 9791 -12878
rect 9825 -12914 9837 -12878
rect 9779 -12948 9837 -12914
rect 9779 -12982 9791 -12948
rect 9825 -12982 9837 -12948
rect 9779 -12996 9837 -12982
rect 10001 -12810 10059 -12796
rect 10001 -12844 10013 -12810
rect 10047 -12844 10059 -12810
rect 10001 -12878 10059 -12844
rect 10001 -12914 10013 -12878
rect 10047 -12914 10059 -12878
rect 10001 -12948 10059 -12914
rect 10001 -12982 10013 -12948
rect 10047 -12982 10059 -12948
rect 10001 -12996 10059 -12982
rect 10259 -12810 10317 -12796
rect 10259 -12844 10271 -12810
rect 10305 -12844 10317 -12810
rect 10259 -12878 10317 -12844
rect 10259 -12914 10271 -12878
rect 10305 -12914 10317 -12878
rect 10259 -12948 10317 -12914
rect 10259 -12982 10271 -12948
rect 10305 -12982 10317 -12948
rect 10259 -12996 10317 -12982
rect 10504 -12808 10562 -12794
rect 10504 -12842 10516 -12808
rect 10550 -12842 10562 -12808
rect 10504 -12876 10562 -12842
rect 10504 -12912 10516 -12876
rect 10550 -12912 10562 -12876
rect 10504 -12946 10562 -12912
rect 10504 -12980 10516 -12946
rect 10550 -12980 10562 -12946
rect 10504 -12994 10562 -12980
rect 10762 -12808 10820 -12794
rect 10762 -12842 10774 -12808
rect 10808 -12842 10820 -12808
rect 10762 -12876 10820 -12842
rect 10762 -12912 10774 -12876
rect 10808 -12912 10820 -12876
rect 10762 -12946 10820 -12912
rect 10762 -12980 10774 -12946
rect 10808 -12980 10820 -12946
rect 10762 -12994 10820 -12980
rect 11014 -12798 11072 -12784
rect 11014 -12832 11026 -12798
rect 11060 -12832 11072 -12798
rect 11014 -12866 11072 -12832
rect 11014 -12902 11026 -12866
rect 11060 -12902 11072 -12866
rect 11014 -12936 11072 -12902
rect 11014 -12970 11026 -12936
rect 11060 -12970 11072 -12936
rect 11014 -12984 11072 -12970
rect 11272 -12798 11330 -12784
rect 11272 -12832 11284 -12798
rect 11318 -12832 11330 -12798
rect 11272 -12866 11330 -12832
rect 11272 -12902 11284 -12866
rect 11318 -12902 11330 -12866
rect 11272 -12936 11330 -12902
rect 11272 -12970 11284 -12936
rect 11318 -12970 11330 -12936
rect 11272 -12984 11330 -12970
rect 11651 -12810 11709 -12796
rect 11651 -12844 11663 -12810
rect 11697 -12844 11709 -12810
rect 11651 -12878 11709 -12844
rect 11651 -12914 11663 -12878
rect 11697 -12914 11709 -12878
rect 11651 -12948 11709 -12914
rect 11651 -12982 11663 -12948
rect 11697 -12982 11709 -12948
rect 11651 -12996 11709 -12982
rect 11909 -12810 11967 -12796
rect 11909 -12844 11921 -12810
rect 11955 -12844 11967 -12810
rect 11909 -12878 11967 -12844
rect 11909 -12914 11921 -12878
rect 11955 -12914 11967 -12878
rect 11909 -12948 11967 -12914
rect 11909 -12982 11921 -12948
rect 11955 -12982 11967 -12948
rect 11909 -12996 11967 -12982
rect 12191 -12810 12249 -12796
rect 12191 -12844 12203 -12810
rect 12237 -12844 12249 -12810
rect 12191 -12878 12249 -12844
rect 12191 -12914 12203 -12878
rect 12237 -12914 12249 -12878
rect 12191 -12948 12249 -12914
rect 12191 -12982 12203 -12948
rect 12237 -12982 12249 -12948
rect 12191 -12996 12249 -12982
rect 12449 -12810 12507 -12796
rect 12449 -12844 12461 -12810
rect 12495 -12844 12507 -12810
rect 12449 -12878 12507 -12844
rect 12449 -12914 12461 -12878
rect 12495 -12914 12507 -12878
rect 12449 -12948 12507 -12914
rect 12449 -12982 12461 -12948
rect 12495 -12982 12507 -12948
rect 12449 -12996 12507 -12982
rect 12671 -12810 12729 -12796
rect 12671 -12844 12683 -12810
rect 12717 -12844 12729 -12810
rect 12671 -12878 12729 -12844
rect 12671 -12914 12683 -12878
rect 12717 -12914 12729 -12878
rect 12671 -12948 12729 -12914
rect 12671 -12982 12683 -12948
rect 12717 -12982 12729 -12948
rect 12671 -12996 12729 -12982
rect 12929 -12810 12987 -12796
rect 12929 -12844 12941 -12810
rect 12975 -12844 12987 -12810
rect 12929 -12878 12987 -12844
rect 12929 -12914 12941 -12878
rect 12975 -12914 12987 -12878
rect 12929 -12948 12987 -12914
rect 12929 -12982 12941 -12948
rect 12975 -12982 12987 -12948
rect 12929 -12996 12987 -12982
rect 13174 -12808 13232 -12794
rect 13174 -12842 13186 -12808
rect 13220 -12842 13232 -12808
rect 13174 -12876 13232 -12842
rect 13174 -12912 13186 -12876
rect 13220 -12912 13232 -12876
rect 13174 -12946 13232 -12912
rect 13174 -12980 13186 -12946
rect 13220 -12980 13232 -12946
rect 13174 -12994 13232 -12980
rect 13432 -12808 13490 -12794
rect 13432 -12842 13444 -12808
rect 13478 -12842 13490 -12808
rect 13432 -12876 13490 -12842
rect 13432 -12912 13444 -12876
rect 13478 -12912 13490 -12876
rect 13432 -12946 13490 -12912
rect 13432 -12980 13444 -12946
rect 13478 -12980 13490 -12946
rect 13432 -12994 13490 -12980
rect 13684 -12798 13742 -12784
rect 13684 -12832 13696 -12798
rect 13730 -12832 13742 -12798
rect 13684 -12866 13742 -12832
rect 13684 -12902 13696 -12866
rect 13730 -12902 13742 -12866
rect 13684 -12936 13742 -12902
rect 13684 -12970 13696 -12936
rect 13730 -12970 13742 -12936
rect 13684 -12984 13742 -12970
rect 13942 -12798 14000 -12784
rect 13942 -12832 13954 -12798
rect 13988 -12832 14000 -12798
rect 13942 -12866 14000 -12832
rect 13942 -12902 13954 -12866
rect 13988 -12902 14000 -12866
rect 13942 -12936 14000 -12902
rect 13942 -12970 13954 -12936
rect 13988 -12970 14000 -12936
rect 13942 -12984 14000 -12970
rect 14314 -12809 14372 -12795
rect 14314 -12843 14326 -12809
rect 14360 -12843 14372 -12809
rect 14314 -12877 14372 -12843
rect 14314 -12913 14326 -12877
rect 14360 -12913 14372 -12877
rect 14314 -12947 14372 -12913
rect 14314 -12981 14326 -12947
rect 14360 -12981 14372 -12947
rect 14314 -12995 14372 -12981
rect 14572 -12809 14630 -12795
rect 14572 -12843 14584 -12809
rect 14618 -12843 14630 -12809
rect 14572 -12877 14630 -12843
rect 14572 -12913 14584 -12877
rect 14618 -12913 14630 -12877
rect 14572 -12947 14630 -12913
rect 14572 -12981 14584 -12947
rect 14618 -12981 14630 -12947
rect 14572 -12995 14630 -12981
rect 14854 -12809 14912 -12795
rect 14854 -12843 14866 -12809
rect 14900 -12843 14912 -12809
rect 14854 -12877 14912 -12843
rect 14854 -12913 14866 -12877
rect 14900 -12913 14912 -12877
rect 14854 -12947 14912 -12913
rect 14854 -12981 14866 -12947
rect 14900 -12981 14912 -12947
rect 14854 -12995 14912 -12981
rect 15112 -12809 15170 -12795
rect 15112 -12843 15124 -12809
rect 15158 -12843 15170 -12809
rect 15112 -12877 15170 -12843
rect 15112 -12913 15124 -12877
rect 15158 -12913 15170 -12877
rect 15112 -12947 15170 -12913
rect 15112 -12981 15124 -12947
rect 15158 -12981 15170 -12947
rect 15112 -12995 15170 -12981
rect 15334 -12809 15392 -12795
rect 15334 -12843 15346 -12809
rect 15380 -12843 15392 -12809
rect 15334 -12877 15392 -12843
rect 15334 -12913 15346 -12877
rect 15380 -12913 15392 -12877
rect 15334 -12947 15392 -12913
rect 15334 -12981 15346 -12947
rect 15380 -12981 15392 -12947
rect 15334 -12995 15392 -12981
rect 15592 -12809 15650 -12795
rect 15592 -12843 15604 -12809
rect 15638 -12843 15650 -12809
rect 15592 -12877 15650 -12843
rect 15592 -12913 15604 -12877
rect 15638 -12913 15650 -12877
rect 15592 -12947 15650 -12913
rect 15592 -12981 15604 -12947
rect 15638 -12981 15650 -12947
rect 15592 -12995 15650 -12981
rect 15837 -12807 15895 -12793
rect 15837 -12841 15849 -12807
rect 15883 -12841 15895 -12807
rect 15837 -12875 15895 -12841
rect 15837 -12911 15849 -12875
rect 15883 -12911 15895 -12875
rect 15837 -12945 15895 -12911
rect 15837 -12979 15849 -12945
rect 15883 -12979 15895 -12945
rect 15837 -12993 15895 -12979
rect 16095 -12807 16153 -12793
rect 16095 -12841 16107 -12807
rect 16141 -12841 16153 -12807
rect 16095 -12875 16153 -12841
rect 16095 -12911 16107 -12875
rect 16141 -12911 16153 -12875
rect 16095 -12945 16153 -12911
rect 16095 -12979 16107 -12945
rect 16141 -12979 16153 -12945
rect 16095 -12993 16153 -12979
rect 16347 -12797 16405 -12783
rect 16347 -12831 16359 -12797
rect 16393 -12831 16405 -12797
rect 16347 -12865 16405 -12831
rect 16347 -12901 16359 -12865
rect 16393 -12901 16405 -12865
rect 16347 -12935 16405 -12901
rect 16347 -12969 16359 -12935
rect 16393 -12969 16405 -12935
rect 16347 -12983 16405 -12969
rect 16605 -12797 16663 -12783
rect 16605 -12831 16617 -12797
rect 16651 -12831 16663 -12797
rect 16605 -12865 16663 -12831
rect 16605 -12901 16617 -12865
rect 16651 -12901 16663 -12865
rect 16605 -12935 16663 -12901
rect 16605 -12969 16617 -12935
rect 16651 -12969 16663 -12935
rect 16605 -12983 16663 -12969
rect 9101 -15365 9159 -15353
rect 9101 -15401 9113 -15365
rect 9147 -15401 9159 -15365
rect 9101 -15435 9159 -15401
rect 9101 -15471 9113 -15435
rect 9147 -15471 9159 -15435
rect 9101 -15505 9159 -15471
rect 9101 -15541 9113 -15505
rect 9147 -15541 9159 -15505
rect 9101 -15553 9159 -15541
rect 9359 -15365 9417 -15353
rect 9359 -15401 9371 -15365
rect 9405 -15401 9417 -15365
rect 9359 -15435 9417 -15401
rect 9359 -15471 9371 -15435
rect 9405 -15471 9417 -15435
rect 9359 -15505 9417 -15471
rect 9359 -15541 9371 -15505
rect 9405 -15541 9417 -15505
rect 9359 -15553 9417 -15541
rect 9617 -15365 9675 -15353
rect 9617 -15401 9629 -15365
rect 9663 -15401 9675 -15365
rect 9617 -15435 9675 -15401
rect 9617 -15471 9629 -15435
rect 9663 -15471 9675 -15435
rect 9617 -15506 9675 -15471
rect 9617 -15542 9629 -15506
rect 9663 -15542 9675 -15506
rect 9617 -15553 9675 -15542
rect 9875 -15365 9933 -15353
rect 9875 -15401 9887 -15365
rect 9921 -15401 9933 -15365
rect 9875 -15435 9933 -15401
rect 9875 -15471 9887 -15435
rect 9921 -15471 9933 -15435
rect 9875 -15505 9933 -15471
rect 9875 -15541 9887 -15505
rect 9921 -15541 9933 -15505
rect 9875 -15553 9933 -15541
rect 10133 -15365 10191 -15353
rect 10133 -15401 10145 -15365
rect 10179 -15401 10191 -15365
rect 10133 -15435 10191 -15401
rect 10133 -15471 10145 -15435
rect 10179 -15471 10191 -15435
rect 10133 -15505 10191 -15471
rect 10133 -15541 10145 -15505
rect 10179 -15541 10191 -15505
rect 10133 -15553 10191 -15541
rect 10391 -15365 10449 -15353
rect 10391 -15401 10403 -15365
rect 10437 -15401 10449 -15365
rect 10391 -15435 10449 -15401
rect 10391 -15471 10403 -15435
rect 10437 -15471 10449 -15435
rect 10391 -15505 10449 -15471
rect 10391 -15541 10403 -15505
rect 10437 -15541 10449 -15505
rect 10391 -15553 10449 -15541
rect 10649 -15365 10707 -15353
rect 10649 -15401 10661 -15365
rect 10695 -15401 10707 -15365
rect 10649 -15435 10707 -15401
rect 10649 -15471 10661 -15435
rect 10695 -15471 10707 -15435
rect 10649 -15505 10707 -15471
rect 10649 -15541 10661 -15505
rect 10695 -15541 10707 -15505
rect 10649 -15553 10707 -15541
rect 10907 -15365 10965 -15353
rect 10907 -15401 10919 -15365
rect 10953 -15401 10965 -15365
rect 10907 -15435 10965 -15401
rect 10907 -15471 10919 -15435
rect 10953 -15471 10965 -15435
rect 10907 -15505 10965 -15471
rect 10907 -15541 10919 -15505
rect 10953 -15541 10965 -15505
rect 10907 -15553 10965 -15541
rect 11165 -15365 11223 -15353
rect 11165 -15401 11177 -15365
rect 11211 -15401 11223 -15365
rect 11165 -15435 11223 -15401
rect 11165 -15471 11177 -15435
rect 11211 -15471 11223 -15435
rect 11165 -15505 11223 -15471
rect 11165 -15541 11177 -15505
rect 11211 -15541 11223 -15505
rect 11165 -15553 11223 -15541
rect 11771 -15365 11829 -15353
rect 11771 -15401 11783 -15365
rect 11817 -15401 11829 -15365
rect 11771 -15435 11829 -15401
rect 11771 -15471 11783 -15435
rect 11817 -15471 11829 -15435
rect 11771 -15505 11829 -15471
rect 11771 -15541 11783 -15505
rect 11817 -15541 11829 -15505
rect 11771 -15553 11829 -15541
rect 12029 -15365 12087 -15353
rect 12029 -15401 12041 -15365
rect 12075 -15401 12087 -15365
rect 12029 -15435 12087 -15401
rect 12029 -15471 12041 -15435
rect 12075 -15471 12087 -15435
rect 12029 -15505 12087 -15471
rect 12029 -15541 12041 -15505
rect 12075 -15541 12087 -15505
rect 12029 -15553 12087 -15541
rect 12287 -15365 12345 -15353
rect 12287 -15401 12299 -15365
rect 12333 -15401 12345 -15365
rect 12287 -15435 12345 -15401
rect 12287 -15471 12299 -15435
rect 12333 -15471 12345 -15435
rect 12287 -15506 12345 -15471
rect 12287 -15542 12299 -15506
rect 12333 -15542 12345 -15506
rect 12287 -15553 12345 -15542
rect 12545 -15365 12603 -15353
rect 12545 -15401 12557 -15365
rect 12591 -15401 12603 -15365
rect 12545 -15435 12603 -15401
rect 12545 -15471 12557 -15435
rect 12591 -15471 12603 -15435
rect 12545 -15505 12603 -15471
rect 12545 -15541 12557 -15505
rect 12591 -15541 12603 -15505
rect 12545 -15553 12603 -15541
rect 12803 -15365 12861 -15353
rect 12803 -15401 12815 -15365
rect 12849 -15401 12861 -15365
rect 12803 -15435 12861 -15401
rect 12803 -15471 12815 -15435
rect 12849 -15471 12861 -15435
rect 12803 -15505 12861 -15471
rect 12803 -15541 12815 -15505
rect 12849 -15541 12861 -15505
rect 12803 -15553 12861 -15541
rect 13061 -15365 13119 -15353
rect 13061 -15401 13073 -15365
rect 13107 -15401 13119 -15365
rect 13061 -15435 13119 -15401
rect 13061 -15471 13073 -15435
rect 13107 -15471 13119 -15435
rect 13061 -15505 13119 -15471
rect 13061 -15541 13073 -15505
rect 13107 -15541 13119 -15505
rect 13061 -15553 13119 -15541
rect 13319 -15365 13377 -15353
rect 13319 -15401 13331 -15365
rect 13365 -15401 13377 -15365
rect 13319 -15435 13377 -15401
rect 13319 -15471 13331 -15435
rect 13365 -15471 13377 -15435
rect 13319 -15505 13377 -15471
rect 13319 -15541 13331 -15505
rect 13365 -15541 13377 -15505
rect 13319 -15553 13377 -15541
rect 13577 -15365 13635 -15353
rect 13577 -15401 13589 -15365
rect 13623 -15401 13635 -15365
rect 13577 -15435 13635 -15401
rect 13577 -15471 13589 -15435
rect 13623 -15471 13635 -15435
rect 13577 -15505 13635 -15471
rect 13577 -15541 13589 -15505
rect 13623 -15541 13635 -15505
rect 13577 -15553 13635 -15541
rect 13835 -15365 13893 -15353
rect 13835 -15401 13847 -15365
rect 13881 -15401 13893 -15365
rect 13835 -15435 13893 -15401
rect 13835 -15471 13847 -15435
rect 13881 -15471 13893 -15435
rect 13835 -15505 13893 -15471
rect 13835 -15541 13847 -15505
rect 13881 -15541 13893 -15505
rect 13835 -15553 13893 -15541
rect 14434 -15364 14492 -15352
rect 14434 -15400 14446 -15364
rect 14480 -15400 14492 -15364
rect 14434 -15434 14492 -15400
rect 14434 -15470 14446 -15434
rect 14480 -15470 14492 -15434
rect 14434 -15504 14492 -15470
rect 14434 -15540 14446 -15504
rect 14480 -15540 14492 -15504
rect 14434 -15552 14492 -15540
rect 14692 -15364 14750 -15352
rect 14692 -15400 14704 -15364
rect 14738 -15400 14750 -15364
rect 14692 -15434 14750 -15400
rect 14692 -15470 14704 -15434
rect 14738 -15470 14750 -15434
rect 14692 -15504 14750 -15470
rect 14692 -15540 14704 -15504
rect 14738 -15540 14750 -15504
rect 14692 -15552 14750 -15540
rect 14950 -15364 15008 -15352
rect 14950 -15400 14962 -15364
rect 14996 -15400 15008 -15364
rect 14950 -15434 15008 -15400
rect 14950 -15470 14962 -15434
rect 14996 -15470 15008 -15434
rect 14950 -15505 15008 -15470
rect 14950 -15541 14962 -15505
rect 14996 -15541 15008 -15505
rect 14950 -15552 15008 -15541
rect 15208 -15364 15266 -15352
rect 15208 -15400 15220 -15364
rect 15254 -15400 15266 -15364
rect 15208 -15434 15266 -15400
rect 15208 -15470 15220 -15434
rect 15254 -15470 15266 -15434
rect 15208 -15504 15266 -15470
rect 15208 -15540 15220 -15504
rect 15254 -15540 15266 -15504
rect 15208 -15552 15266 -15540
rect 15466 -15364 15524 -15352
rect 15466 -15400 15478 -15364
rect 15512 -15400 15524 -15364
rect 15466 -15434 15524 -15400
rect 15466 -15470 15478 -15434
rect 15512 -15470 15524 -15434
rect 15466 -15504 15524 -15470
rect 15466 -15540 15478 -15504
rect 15512 -15540 15524 -15504
rect 15466 -15552 15524 -15540
rect 15724 -15364 15782 -15352
rect 15724 -15400 15736 -15364
rect 15770 -15400 15782 -15364
rect 15724 -15434 15782 -15400
rect 15724 -15470 15736 -15434
rect 15770 -15470 15782 -15434
rect 15724 -15504 15782 -15470
rect 15724 -15540 15736 -15504
rect 15770 -15540 15782 -15504
rect 15724 -15552 15782 -15540
rect 15982 -15364 16040 -15352
rect 15982 -15400 15994 -15364
rect 16028 -15400 16040 -15364
rect 15982 -15434 16040 -15400
rect 15982 -15470 15994 -15434
rect 16028 -15470 16040 -15434
rect 15982 -15504 16040 -15470
rect 15982 -15540 15994 -15504
rect 16028 -15540 16040 -15504
rect 15982 -15552 16040 -15540
rect 16240 -15364 16298 -15352
rect 16240 -15400 16252 -15364
rect 16286 -15400 16298 -15364
rect 16240 -15434 16298 -15400
rect 16240 -15470 16252 -15434
rect 16286 -15470 16298 -15434
rect 16240 -15504 16298 -15470
rect 16240 -15540 16252 -15504
rect 16286 -15540 16298 -15504
rect 16240 -15552 16298 -15540
rect 16498 -15364 16556 -15352
rect 16498 -15400 16510 -15364
rect 16544 -15400 16556 -15364
rect 16498 -15434 16556 -15400
rect 16498 -15470 16510 -15434
rect 16544 -15470 16556 -15434
rect 16498 -15504 16556 -15470
rect 16498 -15540 16510 -15504
rect 16544 -15540 16556 -15504
rect 16498 -15552 16556 -15540
rect 9101 -15783 9159 -15771
rect 9101 -15819 9113 -15783
rect 9147 -15819 9159 -15783
rect 9101 -15853 9159 -15819
rect 9101 -15889 9113 -15853
rect 9147 -15889 9159 -15853
rect 9101 -15923 9159 -15889
rect 9101 -15959 9113 -15923
rect 9147 -15959 9159 -15923
rect 9101 -15971 9159 -15959
rect 9359 -15783 9417 -15771
rect 9359 -15819 9371 -15783
rect 9405 -15819 9417 -15783
rect 9359 -15853 9417 -15819
rect 9359 -15889 9371 -15853
rect 9405 -15889 9417 -15853
rect 9359 -15923 9417 -15889
rect 9359 -15959 9371 -15923
rect 9405 -15959 9417 -15923
rect 9359 -15971 9417 -15959
rect 9617 -15783 9675 -15771
rect 9617 -15819 9629 -15783
rect 9663 -15819 9675 -15783
rect 9617 -15853 9675 -15819
rect 9617 -15889 9629 -15853
rect 9663 -15889 9675 -15853
rect 9617 -15924 9675 -15889
rect 9617 -15960 9629 -15924
rect 9663 -15960 9675 -15924
rect 9617 -15971 9675 -15960
rect 9875 -15783 9933 -15771
rect 9875 -15819 9887 -15783
rect 9921 -15819 9933 -15783
rect 9875 -15853 9933 -15819
rect 9875 -15889 9887 -15853
rect 9921 -15889 9933 -15853
rect 9875 -15923 9933 -15889
rect 9875 -15959 9887 -15923
rect 9921 -15959 9933 -15923
rect 9875 -15971 9933 -15959
rect 10133 -15783 10191 -15771
rect 10133 -15819 10145 -15783
rect 10179 -15819 10191 -15783
rect 10133 -15853 10191 -15819
rect 10133 -15889 10145 -15853
rect 10179 -15889 10191 -15853
rect 10133 -15923 10191 -15889
rect 10133 -15959 10145 -15923
rect 10179 -15959 10191 -15923
rect 10133 -15971 10191 -15959
rect 10391 -15783 10449 -15771
rect 10391 -15819 10403 -15783
rect 10437 -15819 10449 -15783
rect 10391 -15853 10449 -15819
rect 10391 -15889 10403 -15853
rect 10437 -15889 10449 -15853
rect 10391 -15923 10449 -15889
rect 10391 -15959 10403 -15923
rect 10437 -15959 10449 -15923
rect 10391 -15971 10449 -15959
rect 10649 -15783 10707 -15771
rect 10649 -15819 10661 -15783
rect 10695 -15819 10707 -15783
rect 10649 -15853 10707 -15819
rect 10649 -15889 10661 -15853
rect 10695 -15889 10707 -15853
rect 10649 -15923 10707 -15889
rect 10649 -15959 10661 -15923
rect 10695 -15959 10707 -15923
rect 10649 -15971 10707 -15959
rect 10907 -15783 10965 -15771
rect 10907 -15819 10919 -15783
rect 10953 -15819 10965 -15783
rect 10907 -15853 10965 -15819
rect 10907 -15889 10919 -15853
rect 10953 -15889 10965 -15853
rect 10907 -15923 10965 -15889
rect 10907 -15959 10919 -15923
rect 10953 -15959 10965 -15923
rect 10907 -15971 10965 -15959
rect 11165 -15783 11223 -15771
rect 11165 -15819 11177 -15783
rect 11211 -15819 11223 -15783
rect 11165 -15853 11223 -15819
rect 11165 -15889 11177 -15853
rect 11211 -15889 11223 -15853
rect 11165 -15923 11223 -15889
rect 11165 -15959 11177 -15923
rect 11211 -15959 11223 -15923
rect 11165 -15971 11223 -15959
rect 11771 -15783 11829 -15771
rect 11771 -15819 11783 -15783
rect 11817 -15819 11829 -15783
rect 11771 -15853 11829 -15819
rect 11771 -15889 11783 -15853
rect 11817 -15889 11829 -15853
rect 11771 -15923 11829 -15889
rect 11771 -15959 11783 -15923
rect 11817 -15959 11829 -15923
rect 11771 -15971 11829 -15959
rect 12029 -15783 12087 -15771
rect 12029 -15819 12041 -15783
rect 12075 -15819 12087 -15783
rect 12029 -15853 12087 -15819
rect 12029 -15889 12041 -15853
rect 12075 -15889 12087 -15853
rect 12029 -15923 12087 -15889
rect 12029 -15959 12041 -15923
rect 12075 -15959 12087 -15923
rect 12029 -15971 12087 -15959
rect 12287 -15783 12345 -15771
rect 12287 -15819 12299 -15783
rect 12333 -15819 12345 -15783
rect 12287 -15853 12345 -15819
rect 12287 -15889 12299 -15853
rect 12333 -15889 12345 -15853
rect 12287 -15924 12345 -15889
rect 12287 -15960 12299 -15924
rect 12333 -15960 12345 -15924
rect 12287 -15971 12345 -15960
rect 12545 -15783 12603 -15771
rect 12545 -15819 12557 -15783
rect 12591 -15819 12603 -15783
rect 12545 -15853 12603 -15819
rect 12545 -15889 12557 -15853
rect 12591 -15889 12603 -15853
rect 12545 -15923 12603 -15889
rect 12545 -15959 12557 -15923
rect 12591 -15959 12603 -15923
rect 12545 -15971 12603 -15959
rect 12803 -15783 12861 -15771
rect 12803 -15819 12815 -15783
rect 12849 -15819 12861 -15783
rect 12803 -15853 12861 -15819
rect 12803 -15889 12815 -15853
rect 12849 -15889 12861 -15853
rect 12803 -15923 12861 -15889
rect 12803 -15959 12815 -15923
rect 12849 -15959 12861 -15923
rect 12803 -15971 12861 -15959
rect 13061 -15783 13119 -15771
rect 13061 -15819 13073 -15783
rect 13107 -15819 13119 -15783
rect 13061 -15853 13119 -15819
rect 13061 -15889 13073 -15853
rect 13107 -15889 13119 -15853
rect 13061 -15923 13119 -15889
rect 13061 -15959 13073 -15923
rect 13107 -15959 13119 -15923
rect 13061 -15971 13119 -15959
rect 13319 -15783 13377 -15771
rect 13319 -15819 13331 -15783
rect 13365 -15819 13377 -15783
rect 13319 -15853 13377 -15819
rect 13319 -15889 13331 -15853
rect 13365 -15889 13377 -15853
rect 13319 -15923 13377 -15889
rect 13319 -15959 13331 -15923
rect 13365 -15959 13377 -15923
rect 13319 -15971 13377 -15959
rect 13577 -15783 13635 -15771
rect 13577 -15819 13589 -15783
rect 13623 -15819 13635 -15783
rect 13577 -15853 13635 -15819
rect 13577 -15889 13589 -15853
rect 13623 -15889 13635 -15853
rect 13577 -15923 13635 -15889
rect 13577 -15959 13589 -15923
rect 13623 -15959 13635 -15923
rect 13577 -15971 13635 -15959
rect 13835 -15783 13893 -15771
rect 13835 -15819 13847 -15783
rect 13881 -15819 13893 -15783
rect 13835 -15853 13893 -15819
rect 13835 -15889 13847 -15853
rect 13881 -15889 13893 -15853
rect 13835 -15923 13893 -15889
rect 13835 -15959 13847 -15923
rect 13881 -15959 13893 -15923
rect 13835 -15971 13893 -15959
rect 14434 -15782 14492 -15770
rect 14434 -15818 14446 -15782
rect 14480 -15818 14492 -15782
rect 14434 -15852 14492 -15818
rect 14434 -15888 14446 -15852
rect 14480 -15888 14492 -15852
rect 14434 -15922 14492 -15888
rect 14434 -15958 14446 -15922
rect 14480 -15958 14492 -15922
rect 14434 -15970 14492 -15958
rect 14692 -15782 14750 -15770
rect 14692 -15818 14704 -15782
rect 14738 -15818 14750 -15782
rect 14692 -15852 14750 -15818
rect 14692 -15888 14704 -15852
rect 14738 -15888 14750 -15852
rect 14692 -15922 14750 -15888
rect 14692 -15958 14704 -15922
rect 14738 -15958 14750 -15922
rect 14692 -15970 14750 -15958
rect 14950 -15782 15008 -15770
rect 14950 -15818 14962 -15782
rect 14996 -15818 15008 -15782
rect 14950 -15852 15008 -15818
rect 14950 -15888 14962 -15852
rect 14996 -15888 15008 -15852
rect 14950 -15923 15008 -15888
rect 14950 -15959 14962 -15923
rect 14996 -15959 15008 -15923
rect 14950 -15970 15008 -15959
rect 15208 -15782 15266 -15770
rect 15208 -15818 15220 -15782
rect 15254 -15818 15266 -15782
rect 15208 -15852 15266 -15818
rect 15208 -15888 15220 -15852
rect 15254 -15888 15266 -15852
rect 15208 -15922 15266 -15888
rect 15208 -15958 15220 -15922
rect 15254 -15958 15266 -15922
rect 15208 -15970 15266 -15958
rect 15466 -15782 15524 -15770
rect 15466 -15818 15478 -15782
rect 15512 -15818 15524 -15782
rect 15466 -15852 15524 -15818
rect 15466 -15888 15478 -15852
rect 15512 -15888 15524 -15852
rect 15466 -15922 15524 -15888
rect 15466 -15958 15478 -15922
rect 15512 -15958 15524 -15922
rect 15466 -15970 15524 -15958
rect 15724 -15782 15782 -15770
rect 15724 -15818 15736 -15782
rect 15770 -15818 15782 -15782
rect 15724 -15852 15782 -15818
rect 15724 -15888 15736 -15852
rect 15770 -15888 15782 -15852
rect 15724 -15922 15782 -15888
rect 15724 -15958 15736 -15922
rect 15770 -15958 15782 -15922
rect 15724 -15970 15782 -15958
rect 15982 -15782 16040 -15770
rect 15982 -15818 15994 -15782
rect 16028 -15818 16040 -15782
rect 15982 -15852 16040 -15818
rect 15982 -15888 15994 -15852
rect 16028 -15888 16040 -15852
rect 15982 -15922 16040 -15888
rect 15982 -15958 15994 -15922
rect 16028 -15958 16040 -15922
rect 15982 -15970 16040 -15958
rect 16240 -15782 16298 -15770
rect 16240 -15818 16252 -15782
rect 16286 -15818 16298 -15782
rect 16240 -15852 16298 -15818
rect 16240 -15888 16252 -15852
rect 16286 -15888 16298 -15852
rect 16240 -15922 16298 -15888
rect 16240 -15958 16252 -15922
rect 16286 -15958 16298 -15922
rect 16240 -15970 16298 -15958
rect 16498 -15782 16556 -15770
rect 16498 -15818 16510 -15782
rect 16544 -15818 16556 -15782
rect 16498 -15852 16556 -15818
rect 16498 -15888 16510 -15852
rect 16544 -15888 16556 -15852
rect 16498 -15922 16556 -15888
rect 16498 -15958 16510 -15922
rect 16544 -15958 16556 -15922
rect 16498 -15970 16556 -15958
rect 9101 -16201 9159 -16189
rect 9101 -16237 9113 -16201
rect 9147 -16237 9159 -16201
rect 9101 -16271 9159 -16237
rect 9101 -16307 9113 -16271
rect 9147 -16307 9159 -16271
rect 9101 -16341 9159 -16307
rect 9101 -16377 9113 -16341
rect 9147 -16377 9159 -16341
rect 9101 -16389 9159 -16377
rect 9359 -16201 9417 -16189
rect 9359 -16237 9371 -16201
rect 9405 -16237 9417 -16201
rect 9359 -16271 9417 -16237
rect 9359 -16307 9371 -16271
rect 9405 -16307 9417 -16271
rect 9359 -16341 9417 -16307
rect 9359 -16377 9371 -16341
rect 9405 -16377 9417 -16341
rect 9359 -16389 9417 -16377
rect 9617 -16201 9675 -16189
rect 9617 -16237 9629 -16201
rect 9663 -16237 9675 -16201
rect 9617 -16271 9675 -16237
rect 9617 -16307 9629 -16271
rect 9663 -16307 9675 -16271
rect 9617 -16342 9675 -16307
rect 9617 -16378 9629 -16342
rect 9663 -16378 9675 -16342
rect 9617 -16389 9675 -16378
rect 9875 -16201 9933 -16189
rect 9875 -16237 9887 -16201
rect 9921 -16237 9933 -16201
rect 9875 -16271 9933 -16237
rect 9875 -16307 9887 -16271
rect 9921 -16307 9933 -16271
rect 9875 -16341 9933 -16307
rect 9875 -16377 9887 -16341
rect 9921 -16377 9933 -16341
rect 9875 -16389 9933 -16377
rect 10133 -16201 10191 -16189
rect 10133 -16237 10145 -16201
rect 10179 -16237 10191 -16201
rect 10133 -16271 10191 -16237
rect 10133 -16307 10145 -16271
rect 10179 -16307 10191 -16271
rect 10133 -16341 10191 -16307
rect 10133 -16377 10145 -16341
rect 10179 -16377 10191 -16341
rect 10133 -16389 10191 -16377
rect 10391 -16201 10449 -16189
rect 10391 -16237 10403 -16201
rect 10437 -16237 10449 -16201
rect 10391 -16271 10449 -16237
rect 10391 -16307 10403 -16271
rect 10437 -16307 10449 -16271
rect 10391 -16341 10449 -16307
rect 10391 -16377 10403 -16341
rect 10437 -16377 10449 -16341
rect 10391 -16389 10449 -16377
rect 10649 -16201 10707 -16189
rect 10649 -16237 10661 -16201
rect 10695 -16237 10707 -16201
rect 10649 -16271 10707 -16237
rect 10649 -16307 10661 -16271
rect 10695 -16307 10707 -16271
rect 10649 -16341 10707 -16307
rect 10649 -16377 10661 -16341
rect 10695 -16377 10707 -16341
rect 10649 -16389 10707 -16377
rect 10907 -16201 10965 -16189
rect 10907 -16237 10919 -16201
rect 10953 -16237 10965 -16201
rect 10907 -16271 10965 -16237
rect 10907 -16307 10919 -16271
rect 10953 -16307 10965 -16271
rect 10907 -16341 10965 -16307
rect 10907 -16377 10919 -16341
rect 10953 -16377 10965 -16341
rect 10907 -16389 10965 -16377
rect 11165 -16201 11223 -16189
rect 11165 -16237 11177 -16201
rect 11211 -16237 11223 -16201
rect 11165 -16271 11223 -16237
rect 11165 -16307 11177 -16271
rect 11211 -16307 11223 -16271
rect 11165 -16341 11223 -16307
rect 11165 -16377 11177 -16341
rect 11211 -16377 11223 -16341
rect 11165 -16389 11223 -16377
rect 11771 -16201 11829 -16189
rect 11771 -16237 11783 -16201
rect 11817 -16237 11829 -16201
rect 11771 -16271 11829 -16237
rect 11771 -16307 11783 -16271
rect 11817 -16307 11829 -16271
rect 11771 -16341 11829 -16307
rect 11771 -16377 11783 -16341
rect 11817 -16377 11829 -16341
rect 11771 -16389 11829 -16377
rect 12029 -16201 12087 -16189
rect 12029 -16237 12041 -16201
rect 12075 -16237 12087 -16201
rect 12029 -16271 12087 -16237
rect 12029 -16307 12041 -16271
rect 12075 -16307 12087 -16271
rect 12029 -16341 12087 -16307
rect 12029 -16377 12041 -16341
rect 12075 -16377 12087 -16341
rect 12029 -16389 12087 -16377
rect 12287 -16201 12345 -16189
rect 12287 -16237 12299 -16201
rect 12333 -16237 12345 -16201
rect 12287 -16271 12345 -16237
rect 12287 -16307 12299 -16271
rect 12333 -16307 12345 -16271
rect 12287 -16342 12345 -16307
rect 12287 -16378 12299 -16342
rect 12333 -16378 12345 -16342
rect 12287 -16389 12345 -16378
rect 12545 -16201 12603 -16189
rect 12545 -16237 12557 -16201
rect 12591 -16237 12603 -16201
rect 12545 -16271 12603 -16237
rect 12545 -16307 12557 -16271
rect 12591 -16307 12603 -16271
rect 12545 -16341 12603 -16307
rect 12545 -16377 12557 -16341
rect 12591 -16377 12603 -16341
rect 12545 -16389 12603 -16377
rect 12803 -16201 12861 -16189
rect 12803 -16237 12815 -16201
rect 12849 -16237 12861 -16201
rect 12803 -16271 12861 -16237
rect 12803 -16307 12815 -16271
rect 12849 -16307 12861 -16271
rect 12803 -16341 12861 -16307
rect 12803 -16377 12815 -16341
rect 12849 -16377 12861 -16341
rect 12803 -16389 12861 -16377
rect 13061 -16201 13119 -16189
rect 13061 -16237 13073 -16201
rect 13107 -16237 13119 -16201
rect 13061 -16271 13119 -16237
rect 13061 -16307 13073 -16271
rect 13107 -16307 13119 -16271
rect 13061 -16341 13119 -16307
rect 13061 -16377 13073 -16341
rect 13107 -16377 13119 -16341
rect 13061 -16389 13119 -16377
rect 13319 -16201 13377 -16189
rect 13319 -16237 13331 -16201
rect 13365 -16237 13377 -16201
rect 13319 -16271 13377 -16237
rect 13319 -16307 13331 -16271
rect 13365 -16307 13377 -16271
rect 13319 -16341 13377 -16307
rect 13319 -16377 13331 -16341
rect 13365 -16377 13377 -16341
rect 13319 -16389 13377 -16377
rect 13577 -16201 13635 -16189
rect 13577 -16237 13589 -16201
rect 13623 -16237 13635 -16201
rect 13577 -16271 13635 -16237
rect 13577 -16307 13589 -16271
rect 13623 -16307 13635 -16271
rect 13577 -16341 13635 -16307
rect 13577 -16377 13589 -16341
rect 13623 -16377 13635 -16341
rect 13577 -16389 13635 -16377
rect 13835 -16201 13893 -16189
rect 13835 -16237 13847 -16201
rect 13881 -16237 13893 -16201
rect 13835 -16271 13893 -16237
rect 13835 -16307 13847 -16271
rect 13881 -16307 13893 -16271
rect 13835 -16341 13893 -16307
rect 13835 -16377 13847 -16341
rect 13881 -16377 13893 -16341
rect 13835 -16389 13893 -16377
rect 14434 -16200 14492 -16188
rect 14434 -16236 14446 -16200
rect 14480 -16236 14492 -16200
rect 14434 -16270 14492 -16236
rect 14434 -16306 14446 -16270
rect 14480 -16306 14492 -16270
rect 14434 -16340 14492 -16306
rect 14434 -16376 14446 -16340
rect 14480 -16376 14492 -16340
rect 14434 -16388 14492 -16376
rect 14692 -16200 14750 -16188
rect 14692 -16236 14704 -16200
rect 14738 -16236 14750 -16200
rect 14692 -16270 14750 -16236
rect 14692 -16306 14704 -16270
rect 14738 -16306 14750 -16270
rect 14692 -16340 14750 -16306
rect 14692 -16376 14704 -16340
rect 14738 -16376 14750 -16340
rect 14692 -16388 14750 -16376
rect 14950 -16200 15008 -16188
rect 14950 -16236 14962 -16200
rect 14996 -16236 15008 -16200
rect 14950 -16270 15008 -16236
rect 14950 -16306 14962 -16270
rect 14996 -16306 15008 -16270
rect 14950 -16341 15008 -16306
rect 14950 -16377 14962 -16341
rect 14996 -16377 15008 -16341
rect 14950 -16388 15008 -16377
rect 15208 -16200 15266 -16188
rect 15208 -16236 15220 -16200
rect 15254 -16236 15266 -16200
rect 15208 -16270 15266 -16236
rect 15208 -16306 15220 -16270
rect 15254 -16306 15266 -16270
rect 15208 -16340 15266 -16306
rect 15208 -16376 15220 -16340
rect 15254 -16376 15266 -16340
rect 15208 -16388 15266 -16376
rect 15466 -16200 15524 -16188
rect 15466 -16236 15478 -16200
rect 15512 -16236 15524 -16200
rect 15466 -16270 15524 -16236
rect 15466 -16306 15478 -16270
rect 15512 -16306 15524 -16270
rect 15466 -16340 15524 -16306
rect 15466 -16376 15478 -16340
rect 15512 -16376 15524 -16340
rect 15466 -16388 15524 -16376
rect 15724 -16200 15782 -16188
rect 15724 -16236 15736 -16200
rect 15770 -16236 15782 -16200
rect 15724 -16270 15782 -16236
rect 15724 -16306 15736 -16270
rect 15770 -16306 15782 -16270
rect 15724 -16340 15782 -16306
rect 15724 -16376 15736 -16340
rect 15770 -16376 15782 -16340
rect 15724 -16388 15782 -16376
rect 15982 -16200 16040 -16188
rect 15982 -16236 15994 -16200
rect 16028 -16236 16040 -16200
rect 15982 -16270 16040 -16236
rect 15982 -16306 15994 -16270
rect 16028 -16306 16040 -16270
rect 15982 -16340 16040 -16306
rect 15982 -16376 15994 -16340
rect 16028 -16376 16040 -16340
rect 15982 -16388 16040 -16376
rect 16240 -16200 16298 -16188
rect 16240 -16236 16252 -16200
rect 16286 -16236 16298 -16200
rect 16240 -16270 16298 -16236
rect 16240 -16306 16252 -16270
rect 16286 -16306 16298 -16270
rect 16240 -16340 16298 -16306
rect 16240 -16376 16252 -16340
rect 16286 -16376 16298 -16340
rect 16240 -16388 16298 -16376
rect 16498 -16200 16556 -16188
rect 16498 -16236 16510 -16200
rect 16544 -16236 16556 -16200
rect 16498 -16270 16556 -16236
rect 16498 -16306 16510 -16270
rect 16544 -16306 16556 -16270
rect 16498 -16340 16556 -16306
rect 16498 -16376 16510 -16340
rect 16544 -16376 16556 -16340
rect 16498 -16388 16556 -16376
rect 9101 -16619 9159 -16607
rect 9101 -16655 9113 -16619
rect 9147 -16655 9159 -16619
rect 9101 -16689 9159 -16655
rect 9101 -16725 9113 -16689
rect 9147 -16725 9159 -16689
rect 9101 -16759 9159 -16725
rect 9101 -16795 9113 -16759
rect 9147 -16795 9159 -16759
rect 9101 -16807 9159 -16795
rect 9359 -16619 9417 -16607
rect 9359 -16655 9371 -16619
rect 9405 -16655 9417 -16619
rect 9359 -16689 9417 -16655
rect 9359 -16725 9371 -16689
rect 9405 -16725 9417 -16689
rect 9359 -16759 9417 -16725
rect 9359 -16795 9371 -16759
rect 9405 -16795 9417 -16759
rect 9359 -16807 9417 -16795
rect 9617 -16619 9675 -16607
rect 9617 -16655 9629 -16619
rect 9663 -16655 9675 -16619
rect 9617 -16689 9675 -16655
rect 9617 -16725 9629 -16689
rect 9663 -16725 9675 -16689
rect 9617 -16760 9675 -16725
rect 9617 -16796 9629 -16760
rect 9663 -16796 9675 -16760
rect 9617 -16807 9675 -16796
rect 9875 -16619 9933 -16607
rect 9875 -16655 9887 -16619
rect 9921 -16655 9933 -16619
rect 9875 -16689 9933 -16655
rect 9875 -16725 9887 -16689
rect 9921 -16725 9933 -16689
rect 9875 -16759 9933 -16725
rect 9875 -16795 9887 -16759
rect 9921 -16795 9933 -16759
rect 9875 -16807 9933 -16795
rect 10133 -16619 10191 -16607
rect 10133 -16655 10145 -16619
rect 10179 -16655 10191 -16619
rect 10133 -16689 10191 -16655
rect 10133 -16725 10145 -16689
rect 10179 -16725 10191 -16689
rect 10133 -16759 10191 -16725
rect 10133 -16795 10145 -16759
rect 10179 -16795 10191 -16759
rect 10133 -16807 10191 -16795
rect 10391 -16619 10449 -16607
rect 10391 -16655 10403 -16619
rect 10437 -16655 10449 -16619
rect 10391 -16689 10449 -16655
rect 10391 -16725 10403 -16689
rect 10437 -16725 10449 -16689
rect 10391 -16759 10449 -16725
rect 10391 -16795 10403 -16759
rect 10437 -16795 10449 -16759
rect 10391 -16807 10449 -16795
rect 10649 -16619 10707 -16607
rect 10649 -16655 10661 -16619
rect 10695 -16655 10707 -16619
rect 10649 -16689 10707 -16655
rect 10649 -16725 10661 -16689
rect 10695 -16725 10707 -16689
rect 10649 -16759 10707 -16725
rect 10649 -16795 10661 -16759
rect 10695 -16795 10707 -16759
rect 10649 -16807 10707 -16795
rect 10907 -16619 10965 -16607
rect 10907 -16655 10919 -16619
rect 10953 -16655 10965 -16619
rect 10907 -16689 10965 -16655
rect 10907 -16725 10919 -16689
rect 10953 -16725 10965 -16689
rect 10907 -16759 10965 -16725
rect 10907 -16795 10919 -16759
rect 10953 -16795 10965 -16759
rect 10907 -16807 10965 -16795
rect 11165 -16619 11223 -16607
rect 11165 -16655 11177 -16619
rect 11211 -16655 11223 -16619
rect 11165 -16689 11223 -16655
rect 11165 -16725 11177 -16689
rect 11211 -16725 11223 -16689
rect 11165 -16759 11223 -16725
rect 11165 -16795 11177 -16759
rect 11211 -16795 11223 -16759
rect 11165 -16807 11223 -16795
rect 11771 -16619 11829 -16607
rect 11771 -16655 11783 -16619
rect 11817 -16655 11829 -16619
rect 11771 -16689 11829 -16655
rect 11771 -16725 11783 -16689
rect 11817 -16725 11829 -16689
rect 11771 -16759 11829 -16725
rect 11771 -16795 11783 -16759
rect 11817 -16795 11829 -16759
rect 11771 -16807 11829 -16795
rect 12029 -16619 12087 -16607
rect 12029 -16655 12041 -16619
rect 12075 -16655 12087 -16619
rect 12029 -16689 12087 -16655
rect 12029 -16725 12041 -16689
rect 12075 -16725 12087 -16689
rect 12029 -16759 12087 -16725
rect 12029 -16795 12041 -16759
rect 12075 -16795 12087 -16759
rect 12029 -16807 12087 -16795
rect 12287 -16619 12345 -16607
rect 12287 -16655 12299 -16619
rect 12333 -16655 12345 -16619
rect 12287 -16689 12345 -16655
rect 12287 -16725 12299 -16689
rect 12333 -16725 12345 -16689
rect 12287 -16760 12345 -16725
rect 12287 -16796 12299 -16760
rect 12333 -16796 12345 -16760
rect 12287 -16807 12345 -16796
rect 12545 -16619 12603 -16607
rect 12545 -16655 12557 -16619
rect 12591 -16655 12603 -16619
rect 12545 -16689 12603 -16655
rect 12545 -16725 12557 -16689
rect 12591 -16725 12603 -16689
rect 12545 -16759 12603 -16725
rect 12545 -16795 12557 -16759
rect 12591 -16795 12603 -16759
rect 12545 -16807 12603 -16795
rect 12803 -16619 12861 -16607
rect 12803 -16655 12815 -16619
rect 12849 -16655 12861 -16619
rect 12803 -16689 12861 -16655
rect 12803 -16725 12815 -16689
rect 12849 -16725 12861 -16689
rect 12803 -16759 12861 -16725
rect 12803 -16795 12815 -16759
rect 12849 -16795 12861 -16759
rect 12803 -16807 12861 -16795
rect 13061 -16619 13119 -16607
rect 13061 -16655 13073 -16619
rect 13107 -16655 13119 -16619
rect 13061 -16689 13119 -16655
rect 13061 -16725 13073 -16689
rect 13107 -16725 13119 -16689
rect 13061 -16759 13119 -16725
rect 13061 -16795 13073 -16759
rect 13107 -16795 13119 -16759
rect 13061 -16807 13119 -16795
rect 13319 -16619 13377 -16607
rect 13319 -16655 13331 -16619
rect 13365 -16655 13377 -16619
rect 13319 -16689 13377 -16655
rect 13319 -16725 13331 -16689
rect 13365 -16725 13377 -16689
rect 13319 -16759 13377 -16725
rect 13319 -16795 13331 -16759
rect 13365 -16795 13377 -16759
rect 13319 -16807 13377 -16795
rect 13577 -16619 13635 -16607
rect 13577 -16655 13589 -16619
rect 13623 -16655 13635 -16619
rect 13577 -16689 13635 -16655
rect 13577 -16725 13589 -16689
rect 13623 -16725 13635 -16689
rect 13577 -16759 13635 -16725
rect 13577 -16795 13589 -16759
rect 13623 -16795 13635 -16759
rect 13577 -16807 13635 -16795
rect 13835 -16619 13893 -16607
rect 13835 -16655 13847 -16619
rect 13881 -16655 13893 -16619
rect 13835 -16689 13893 -16655
rect 13835 -16725 13847 -16689
rect 13881 -16725 13893 -16689
rect 13835 -16759 13893 -16725
rect 13835 -16795 13847 -16759
rect 13881 -16795 13893 -16759
rect 13835 -16807 13893 -16795
rect 14434 -16618 14492 -16606
rect 14434 -16654 14446 -16618
rect 14480 -16654 14492 -16618
rect 14434 -16688 14492 -16654
rect 14434 -16724 14446 -16688
rect 14480 -16724 14492 -16688
rect 14434 -16758 14492 -16724
rect 14434 -16794 14446 -16758
rect 14480 -16794 14492 -16758
rect 14434 -16806 14492 -16794
rect 14692 -16618 14750 -16606
rect 14692 -16654 14704 -16618
rect 14738 -16654 14750 -16618
rect 14692 -16688 14750 -16654
rect 14692 -16724 14704 -16688
rect 14738 -16724 14750 -16688
rect 14692 -16758 14750 -16724
rect 14692 -16794 14704 -16758
rect 14738 -16794 14750 -16758
rect 14692 -16806 14750 -16794
rect 14950 -16618 15008 -16606
rect 14950 -16654 14962 -16618
rect 14996 -16654 15008 -16618
rect 14950 -16688 15008 -16654
rect 14950 -16724 14962 -16688
rect 14996 -16724 15008 -16688
rect 14950 -16759 15008 -16724
rect 14950 -16795 14962 -16759
rect 14996 -16795 15008 -16759
rect 14950 -16806 15008 -16795
rect 15208 -16618 15266 -16606
rect 15208 -16654 15220 -16618
rect 15254 -16654 15266 -16618
rect 15208 -16688 15266 -16654
rect 15208 -16724 15220 -16688
rect 15254 -16724 15266 -16688
rect 15208 -16758 15266 -16724
rect 15208 -16794 15220 -16758
rect 15254 -16794 15266 -16758
rect 15208 -16806 15266 -16794
rect 15466 -16618 15524 -16606
rect 15466 -16654 15478 -16618
rect 15512 -16654 15524 -16618
rect 15466 -16688 15524 -16654
rect 15466 -16724 15478 -16688
rect 15512 -16724 15524 -16688
rect 15466 -16758 15524 -16724
rect 15466 -16794 15478 -16758
rect 15512 -16794 15524 -16758
rect 15466 -16806 15524 -16794
rect 15724 -16618 15782 -16606
rect 15724 -16654 15736 -16618
rect 15770 -16654 15782 -16618
rect 15724 -16688 15782 -16654
rect 15724 -16724 15736 -16688
rect 15770 -16724 15782 -16688
rect 15724 -16758 15782 -16724
rect 15724 -16794 15736 -16758
rect 15770 -16794 15782 -16758
rect 15724 -16806 15782 -16794
rect 15982 -16618 16040 -16606
rect 15982 -16654 15994 -16618
rect 16028 -16654 16040 -16618
rect 15982 -16688 16040 -16654
rect 15982 -16724 15994 -16688
rect 16028 -16724 16040 -16688
rect 15982 -16758 16040 -16724
rect 15982 -16794 15994 -16758
rect 16028 -16794 16040 -16758
rect 15982 -16806 16040 -16794
rect 16240 -16618 16298 -16606
rect 16240 -16654 16252 -16618
rect 16286 -16654 16298 -16618
rect 16240 -16688 16298 -16654
rect 16240 -16724 16252 -16688
rect 16286 -16724 16298 -16688
rect 16240 -16758 16298 -16724
rect 16240 -16794 16252 -16758
rect 16286 -16794 16298 -16758
rect 16240 -16806 16298 -16794
rect 16498 -16618 16556 -16606
rect 16498 -16654 16510 -16618
rect 16544 -16654 16556 -16618
rect 16498 -16688 16556 -16654
rect 16498 -16724 16510 -16688
rect 16544 -16724 16556 -16688
rect 16498 -16758 16556 -16724
rect 16498 -16794 16510 -16758
rect 16544 -16794 16556 -16758
rect 16498 -16806 16556 -16794
rect 9101 -17037 9159 -17025
rect 9101 -17073 9113 -17037
rect 9147 -17073 9159 -17037
rect 9101 -17107 9159 -17073
rect 9101 -17143 9113 -17107
rect 9147 -17143 9159 -17107
rect 9101 -17177 9159 -17143
rect 9101 -17213 9113 -17177
rect 9147 -17213 9159 -17177
rect 9101 -17225 9159 -17213
rect 9359 -17037 9417 -17025
rect 9359 -17073 9371 -17037
rect 9405 -17073 9417 -17037
rect 9359 -17107 9417 -17073
rect 9359 -17143 9371 -17107
rect 9405 -17143 9417 -17107
rect 9359 -17177 9417 -17143
rect 9359 -17213 9371 -17177
rect 9405 -17213 9417 -17177
rect 9359 -17225 9417 -17213
rect 9617 -17037 9675 -17025
rect 9617 -17073 9629 -17037
rect 9663 -17073 9675 -17037
rect 9617 -17107 9675 -17073
rect 9617 -17143 9629 -17107
rect 9663 -17143 9675 -17107
rect 9617 -17178 9675 -17143
rect 9617 -17214 9629 -17178
rect 9663 -17214 9675 -17178
rect 9617 -17225 9675 -17214
rect 9875 -17037 9933 -17025
rect 9875 -17073 9887 -17037
rect 9921 -17073 9933 -17037
rect 9875 -17107 9933 -17073
rect 9875 -17143 9887 -17107
rect 9921 -17143 9933 -17107
rect 9875 -17177 9933 -17143
rect 9875 -17213 9887 -17177
rect 9921 -17213 9933 -17177
rect 9875 -17225 9933 -17213
rect 10133 -17037 10191 -17025
rect 10133 -17073 10145 -17037
rect 10179 -17073 10191 -17037
rect 10133 -17107 10191 -17073
rect 10133 -17143 10145 -17107
rect 10179 -17143 10191 -17107
rect 10133 -17177 10191 -17143
rect 10133 -17213 10145 -17177
rect 10179 -17213 10191 -17177
rect 10133 -17225 10191 -17213
rect 10391 -17037 10449 -17025
rect 10391 -17073 10403 -17037
rect 10437 -17073 10449 -17037
rect 10391 -17107 10449 -17073
rect 10391 -17143 10403 -17107
rect 10437 -17143 10449 -17107
rect 10391 -17177 10449 -17143
rect 10391 -17213 10403 -17177
rect 10437 -17213 10449 -17177
rect 10391 -17225 10449 -17213
rect 10649 -17037 10707 -17025
rect 10649 -17073 10661 -17037
rect 10695 -17073 10707 -17037
rect 10649 -17107 10707 -17073
rect 10649 -17143 10661 -17107
rect 10695 -17143 10707 -17107
rect 10649 -17177 10707 -17143
rect 10649 -17213 10661 -17177
rect 10695 -17213 10707 -17177
rect 10649 -17225 10707 -17213
rect 10907 -17037 10965 -17025
rect 10907 -17073 10919 -17037
rect 10953 -17073 10965 -17037
rect 10907 -17107 10965 -17073
rect 10907 -17143 10919 -17107
rect 10953 -17143 10965 -17107
rect 10907 -17177 10965 -17143
rect 10907 -17213 10919 -17177
rect 10953 -17213 10965 -17177
rect 10907 -17225 10965 -17213
rect 11165 -17037 11223 -17025
rect 11165 -17073 11177 -17037
rect 11211 -17073 11223 -17037
rect 11165 -17107 11223 -17073
rect 11165 -17143 11177 -17107
rect 11211 -17143 11223 -17107
rect 11165 -17177 11223 -17143
rect 11165 -17213 11177 -17177
rect 11211 -17213 11223 -17177
rect 11165 -17225 11223 -17213
rect 11771 -17037 11829 -17025
rect 11771 -17073 11783 -17037
rect 11817 -17073 11829 -17037
rect 11771 -17107 11829 -17073
rect 11771 -17143 11783 -17107
rect 11817 -17143 11829 -17107
rect 11771 -17177 11829 -17143
rect 11771 -17213 11783 -17177
rect 11817 -17213 11829 -17177
rect 11771 -17225 11829 -17213
rect 12029 -17037 12087 -17025
rect 12029 -17073 12041 -17037
rect 12075 -17073 12087 -17037
rect 12029 -17107 12087 -17073
rect 12029 -17143 12041 -17107
rect 12075 -17143 12087 -17107
rect 12029 -17177 12087 -17143
rect 12029 -17213 12041 -17177
rect 12075 -17213 12087 -17177
rect 12029 -17225 12087 -17213
rect 12287 -17037 12345 -17025
rect 12287 -17073 12299 -17037
rect 12333 -17073 12345 -17037
rect 12287 -17107 12345 -17073
rect 12287 -17143 12299 -17107
rect 12333 -17143 12345 -17107
rect 12287 -17178 12345 -17143
rect 12287 -17214 12299 -17178
rect 12333 -17214 12345 -17178
rect 12287 -17225 12345 -17214
rect 12545 -17037 12603 -17025
rect 12545 -17073 12557 -17037
rect 12591 -17073 12603 -17037
rect 12545 -17107 12603 -17073
rect 12545 -17143 12557 -17107
rect 12591 -17143 12603 -17107
rect 12545 -17177 12603 -17143
rect 12545 -17213 12557 -17177
rect 12591 -17213 12603 -17177
rect 12545 -17225 12603 -17213
rect 12803 -17037 12861 -17025
rect 12803 -17073 12815 -17037
rect 12849 -17073 12861 -17037
rect 12803 -17107 12861 -17073
rect 12803 -17143 12815 -17107
rect 12849 -17143 12861 -17107
rect 12803 -17177 12861 -17143
rect 12803 -17213 12815 -17177
rect 12849 -17213 12861 -17177
rect 12803 -17225 12861 -17213
rect 13061 -17037 13119 -17025
rect 13061 -17073 13073 -17037
rect 13107 -17073 13119 -17037
rect 13061 -17107 13119 -17073
rect 13061 -17143 13073 -17107
rect 13107 -17143 13119 -17107
rect 13061 -17177 13119 -17143
rect 13061 -17213 13073 -17177
rect 13107 -17213 13119 -17177
rect 13061 -17225 13119 -17213
rect 13319 -17037 13377 -17025
rect 13319 -17073 13331 -17037
rect 13365 -17073 13377 -17037
rect 13319 -17107 13377 -17073
rect 13319 -17143 13331 -17107
rect 13365 -17143 13377 -17107
rect 13319 -17177 13377 -17143
rect 13319 -17213 13331 -17177
rect 13365 -17213 13377 -17177
rect 13319 -17225 13377 -17213
rect 13577 -17037 13635 -17025
rect 13577 -17073 13589 -17037
rect 13623 -17073 13635 -17037
rect 13577 -17107 13635 -17073
rect 13577 -17143 13589 -17107
rect 13623 -17143 13635 -17107
rect 13577 -17177 13635 -17143
rect 13577 -17213 13589 -17177
rect 13623 -17213 13635 -17177
rect 13577 -17225 13635 -17213
rect 13835 -17037 13893 -17025
rect 13835 -17073 13847 -17037
rect 13881 -17073 13893 -17037
rect 13835 -17107 13893 -17073
rect 13835 -17143 13847 -17107
rect 13881 -17143 13893 -17107
rect 13835 -17177 13893 -17143
rect 13835 -17213 13847 -17177
rect 13881 -17213 13893 -17177
rect 13835 -17225 13893 -17213
rect 14434 -17036 14492 -17024
rect 14434 -17072 14446 -17036
rect 14480 -17072 14492 -17036
rect 14434 -17106 14492 -17072
rect 14434 -17142 14446 -17106
rect 14480 -17142 14492 -17106
rect 14434 -17176 14492 -17142
rect 14434 -17212 14446 -17176
rect 14480 -17212 14492 -17176
rect 14434 -17224 14492 -17212
rect 14692 -17036 14750 -17024
rect 14692 -17072 14704 -17036
rect 14738 -17072 14750 -17036
rect 14692 -17106 14750 -17072
rect 14692 -17142 14704 -17106
rect 14738 -17142 14750 -17106
rect 14692 -17176 14750 -17142
rect 14692 -17212 14704 -17176
rect 14738 -17212 14750 -17176
rect 14692 -17224 14750 -17212
rect 14950 -17036 15008 -17024
rect 14950 -17072 14962 -17036
rect 14996 -17072 15008 -17036
rect 14950 -17106 15008 -17072
rect 14950 -17142 14962 -17106
rect 14996 -17142 15008 -17106
rect 14950 -17177 15008 -17142
rect 14950 -17213 14962 -17177
rect 14996 -17213 15008 -17177
rect 14950 -17224 15008 -17213
rect 15208 -17036 15266 -17024
rect 15208 -17072 15220 -17036
rect 15254 -17072 15266 -17036
rect 15208 -17106 15266 -17072
rect 15208 -17142 15220 -17106
rect 15254 -17142 15266 -17106
rect 15208 -17176 15266 -17142
rect 15208 -17212 15220 -17176
rect 15254 -17212 15266 -17176
rect 15208 -17224 15266 -17212
rect 15466 -17036 15524 -17024
rect 15466 -17072 15478 -17036
rect 15512 -17072 15524 -17036
rect 15466 -17106 15524 -17072
rect 15466 -17142 15478 -17106
rect 15512 -17142 15524 -17106
rect 15466 -17176 15524 -17142
rect 15466 -17212 15478 -17176
rect 15512 -17212 15524 -17176
rect 15466 -17224 15524 -17212
rect 15724 -17036 15782 -17024
rect 15724 -17072 15736 -17036
rect 15770 -17072 15782 -17036
rect 15724 -17106 15782 -17072
rect 15724 -17142 15736 -17106
rect 15770 -17142 15782 -17106
rect 15724 -17176 15782 -17142
rect 15724 -17212 15736 -17176
rect 15770 -17212 15782 -17176
rect 15724 -17224 15782 -17212
rect 15982 -17036 16040 -17024
rect 15982 -17072 15994 -17036
rect 16028 -17072 16040 -17036
rect 15982 -17106 16040 -17072
rect 15982 -17142 15994 -17106
rect 16028 -17142 16040 -17106
rect 15982 -17176 16040 -17142
rect 15982 -17212 15994 -17176
rect 16028 -17212 16040 -17176
rect 15982 -17224 16040 -17212
rect 16240 -17036 16298 -17024
rect 16240 -17072 16252 -17036
rect 16286 -17072 16298 -17036
rect 16240 -17106 16298 -17072
rect 16240 -17142 16252 -17106
rect 16286 -17142 16298 -17106
rect 16240 -17176 16298 -17142
rect 16240 -17212 16252 -17176
rect 16286 -17212 16298 -17176
rect 16240 -17224 16298 -17212
rect 16498 -17036 16556 -17024
rect 16498 -17072 16510 -17036
rect 16544 -17072 16556 -17036
rect 16498 -17106 16556 -17072
rect 16498 -17142 16510 -17106
rect 16544 -17142 16556 -17106
rect 16498 -17176 16556 -17142
rect 16498 -17212 16510 -17176
rect 16544 -17212 16556 -17176
rect 16498 -17224 16556 -17212
rect 9101 -17455 9159 -17443
rect 9101 -17491 9113 -17455
rect 9147 -17491 9159 -17455
rect 9101 -17525 9159 -17491
rect 9101 -17561 9113 -17525
rect 9147 -17561 9159 -17525
rect 9101 -17595 9159 -17561
rect 9101 -17631 9113 -17595
rect 9147 -17631 9159 -17595
rect 9101 -17643 9159 -17631
rect 9359 -17455 9417 -17443
rect 9359 -17491 9371 -17455
rect 9405 -17491 9417 -17455
rect 9359 -17525 9417 -17491
rect 9359 -17561 9371 -17525
rect 9405 -17561 9417 -17525
rect 9359 -17595 9417 -17561
rect 9359 -17631 9371 -17595
rect 9405 -17631 9417 -17595
rect 9359 -17643 9417 -17631
rect 9617 -17455 9675 -17443
rect 9617 -17491 9629 -17455
rect 9663 -17491 9675 -17455
rect 9617 -17525 9675 -17491
rect 9617 -17561 9629 -17525
rect 9663 -17561 9675 -17525
rect 9617 -17596 9675 -17561
rect 9617 -17632 9629 -17596
rect 9663 -17632 9675 -17596
rect 9617 -17643 9675 -17632
rect 9875 -17455 9933 -17443
rect 9875 -17491 9887 -17455
rect 9921 -17491 9933 -17455
rect 9875 -17525 9933 -17491
rect 9875 -17561 9887 -17525
rect 9921 -17561 9933 -17525
rect 9875 -17595 9933 -17561
rect 9875 -17631 9887 -17595
rect 9921 -17631 9933 -17595
rect 9875 -17643 9933 -17631
rect 10133 -17455 10191 -17443
rect 10133 -17491 10145 -17455
rect 10179 -17491 10191 -17455
rect 10133 -17525 10191 -17491
rect 10133 -17561 10145 -17525
rect 10179 -17561 10191 -17525
rect 10133 -17595 10191 -17561
rect 10133 -17631 10145 -17595
rect 10179 -17631 10191 -17595
rect 10133 -17643 10191 -17631
rect 10391 -17455 10449 -17443
rect 10391 -17491 10403 -17455
rect 10437 -17491 10449 -17455
rect 10391 -17525 10449 -17491
rect 10391 -17561 10403 -17525
rect 10437 -17561 10449 -17525
rect 10391 -17595 10449 -17561
rect 10391 -17631 10403 -17595
rect 10437 -17631 10449 -17595
rect 10391 -17643 10449 -17631
rect 10649 -17455 10707 -17443
rect 10649 -17491 10661 -17455
rect 10695 -17491 10707 -17455
rect 10649 -17525 10707 -17491
rect 10649 -17561 10661 -17525
rect 10695 -17561 10707 -17525
rect 10649 -17595 10707 -17561
rect 10649 -17631 10661 -17595
rect 10695 -17631 10707 -17595
rect 10649 -17643 10707 -17631
rect 10907 -17455 10965 -17443
rect 10907 -17491 10919 -17455
rect 10953 -17491 10965 -17455
rect 10907 -17525 10965 -17491
rect 10907 -17561 10919 -17525
rect 10953 -17561 10965 -17525
rect 10907 -17595 10965 -17561
rect 10907 -17631 10919 -17595
rect 10953 -17631 10965 -17595
rect 10907 -17643 10965 -17631
rect 11165 -17455 11223 -17443
rect 11165 -17491 11177 -17455
rect 11211 -17491 11223 -17455
rect 11165 -17525 11223 -17491
rect 11165 -17561 11177 -17525
rect 11211 -17561 11223 -17525
rect 11165 -17595 11223 -17561
rect 11165 -17631 11177 -17595
rect 11211 -17631 11223 -17595
rect 11165 -17643 11223 -17631
rect 11771 -17455 11829 -17443
rect 11771 -17491 11783 -17455
rect 11817 -17491 11829 -17455
rect 11771 -17525 11829 -17491
rect 11771 -17561 11783 -17525
rect 11817 -17561 11829 -17525
rect 11771 -17595 11829 -17561
rect 11771 -17631 11783 -17595
rect 11817 -17631 11829 -17595
rect 11771 -17643 11829 -17631
rect 12029 -17455 12087 -17443
rect 12029 -17491 12041 -17455
rect 12075 -17491 12087 -17455
rect 12029 -17525 12087 -17491
rect 12029 -17561 12041 -17525
rect 12075 -17561 12087 -17525
rect 12029 -17595 12087 -17561
rect 12029 -17631 12041 -17595
rect 12075 -17631 12087 -17595
rect 12029 -17643 12087 -17631
rect 12287 -17455 12345 -17443
rect 12287 -17491 12299 -17455
rect 12333 -17491 12345 -17455
rect 12287 -17525 12345 -17491
rect 12287 -17561 12299 -17525
rect 12333 -17561 12345 -17525
rect 12287 -17596 12345 -17561
rect 12287 -17632 12299 -17596
rect 12333 -17632 12345 -17596
rect 12287 -17643 12345 -17632
rect 12545 -17455 12603 -17443
rect 12545 -17491 12557 -17455
rect 12591 -17491 12603 -17455
rect 12545 -17525 12603 -17491
rect 12545 -17561 12557 -17525
rect 12591 -17561 12603 -17525
rect 12545 -17595 12603 -17561
rect 12545 -17631 12557 -17595
rect 12591 -17631 12603 -17595
rect 12545 -17643 12603 -17631
rect 12803 -17455 12861 -17443
rect 12803 -17491 12815 -17455
rect 12849 -17491 12861 -17455
rect 12803 -17525 12861 -17491
rect 12803 -17561 12815 -17525
rect 12849 -17561 12861 -17525
rect 12803 -17595 12861 -17561
rect 12803 -17631 12815 -17595
rect 12849 -17631 12861 -17595
rect 12803 -17643 12861 -17631
rect 13061 -17455 13119 -17443
rect 13061 -17491 13073 -17455
rect 13107 -17491 13119 -17455
rect 13061 -17525 13119 -17491
rect 13061 -17561 13073 -17525
rect 13107 -17561 13119 -17525
rect 13061 -17595 13119 -17561
rect 13061 -17631 13073 -17595
rect 13107 -17631 13119 -17595
rect 13061 -17643 13119 -17631
rect 13319 -17455 13377 -17443
rect 13319 -17491 13331 -17455
rect 13365 -17491 13377 -17455
rect 13319 -17525 13377 -17491
rect 13319 -17561 13331 -17525
rect 13365 -17561 13377 -17525
rect 13319 -17595 13377 -17561
rect 13319 -17631 13331 -17595
rect 13365 -17631 13377 -17595
rect 13319 -17643 13377 -17631
rect 13577 -17455 13635 -17443
rect 13577 -17491 13589 -17455
rect 13623 -17491 13635 -17455
rect 13577 -17525 13635 -17491
rect 13577 -17561 13589 -17525
rect 13623 -17561 13635 -17525
rect 13577 -17595 13635 -17561
rect 13577 -17631 13589 -17595
rect 13623 -17631 13635 -17595
rect 13577 -17643 13635 -17631
rect 13835 -17455 13893 -17443
rect 13835 -17491 13847 -17455
rect 13881 -17491 13893 -17455
rect 13835 -17525 13893 -17491
rect 13835 -17561 13847 -17525
rect 13881 -17561 13893 -17525
rect 13835 -17595 13893 -17561
rect 13835 -17631 13847 -17595
rect 13881 -17631 13893 -17595
rect 13835 -17643 13893 -17631
rect 14434 -17454 14492 -17442
rect 14434 -17490 14446 -17454
rect 14480 -17490 14492 -17454
rect 14434 -17524 14492 -17490
rect 14434 -17560 14446 -17524
rect 14480 -17560 14492 -17524
rect 14434 -17594 14492 -17560
rect 14434 -17630 14446 -17594
rect 14480 -17630 14492 -17594
rect 14434 -17642 14492 -17630
rect 14692 -17454 14750 -17442
rect 14692 -17490 14704 -17454
rect 14738 -17490 14750 -17454
rect 14692 -17524 14750 -17490
rect 14692 -17560 14704 -17524
rect 14738 -17560 14750 -17524
rect 14692 -17594 14750 -17560
rect 14692 -17630 14704 -17594
rect 14738 -17630 14750 -17594
rect 14692 -17642 14750 -17630
rect 14950 -17454 15008 -17442
rect 14950 -17490 14962 -17454
rect 14996 -17490 15008 -17454
rect 14950 -17524 15008 -17490
rect 14950 -17560 14962 -17524
rect 14996 -17560 15008 -17524
rect 14950 -17595 15008 -17560
rect 14950 -17631 14962 -17595
rect 14996 -17631 15008 -17595
rect 14950 -17642 15008 -17631
rect 15208 -17454 15266 -17442
rect 15208 -17490 15220 -17454
rect 15254 -17490 15266 -17454
rect 15208 -17524 15266 -17490
rect 15208 -17560 15220 -17524
rect 15254 -17560 15266 -17524
rect 15208 -17594 15266 -17560
rect 15208 -17630 15220 -17594
rect 15254 -17630 15266 -17594
rect 15208 -17642 15266 -17630
rect 15466 -17454 15524 -17442
rect 15466 -17490 15478 -17454
rect 15512 -17490 15524 -17454
rect 15466 -17524 15524 -17490
rect 15466 -17560 15478 -17524
rect 15512 -17560 15524 -17524
rect 15466 -17594 15524 -17560
rect 15466 -17630 15478 -17594
rect 15512 -17630 15524 -17594
rect 15466 -17642 15524 -17630
rect 15724 -17454 15782 -17442
rect 15724 -17490 15736 -17454
rect 15770 -17490 15782 -17454
rect 15724 -17524 15782 -17490
rect 15724 -17560 15736 -17524
rect 15770 -17560 15782 -17524
rect 15724 -17594 15782 -17560
rect 15724 -17630 15736 -17594
rect 15770 -17630 15782 -17594
rect 15724 -17642 15782 -17630
rect 15982 -17454 16040 -17442
rect 15982 -17490 15994 -17454
rect 16028 -17490 16040 -17454
rect 15982 -17524 16040 -17490
rect 15982 -17560 15994 -17524
rect 16028 -17560 16040 -17524
rect 15982 -17594 16040 -17560
rect 15982 -17630 15994 -17594
rect 16028 -17630 16040 -17594
rect 15982 -17642 16040 -17630
rect 16240 -17454 16298 -17442
rect 16240 -17490 16252 -17454
rect 16286 -17490 16298 -17454
rect 16240 -17524 16298 -17490
rect 16240 -17560 16252 -17524
rect 16286 -17560 16298 -17524
rect 16240 -17594 16298 -17560
rect 16240 -17630 16252 -17594
rect 16286 -17630 16298 -17594
rect 16240 -17642 16298 -17630
rect 16498 -17454 16556 -17442
rect 16498 -17490 16510 -17454
rect 16544 -17490 16556 -17454
rect 16498 -17524 16556 -17490
rect 16498 -17560 16510 -17524
rect 16544 -17560 16556 -17524
rect 16498 -17594 16556 -17560
rect 16498 -17630 16510 -17594
rect 16544 -17630 16556 -17594
rect 16498 -17642 16556 -17630
rect 9101 -17873 9159 -17861
rect 9101 -17909 9113 -17873
rect 9147 -17909 9159 -17873
rect 9101 -17943 9159 -17909
rect 9101 -17979 9113 -17943
rect 9147 -17979 9159 -17943
rect 9101 -18013 9159 -17979
rect 9101 -18049 9113 -18013
rect 9147 -18049 9159 -18013
rect 9101 -18061 9159 -18049
rect 9359 -17873 9417 -17861
rect 9359 -17909 9371 -17873
rect 9405 -17909 9417 -17873
rect 9359 -17943 9417 -17909
rect 9359 -17979 9371 -17943
rect 9405 -17979 9417 -17943
rect 9359 -18013 9417 -17979
rect 9359 -18049 9371 -18013
rect 9405 -18049 9417 -18013
rect 9359 -18061 9417 -18049
rect 9617 -17873 9675 -17861
rect 9617 -17909 9629 -17873
rect 9663 -17909 9675 -17873
rect 9617 -17943 9675 -17909
rect 9617 -17979 9629 -17943
rect 9663 -17979 9675 -17943
rect 9617 -18014 9675 -17979
rect 9617 -18050 9629 -18014
rect 9663 -18050 9675 -18014
rect 9617 -18061 9675 -18050
rect 9875 -17873 9933 -17861
rect 9875 -17909 9887 -17873
rect 9921 -17909 9933 -17873
rect 9875 -17943 9933 -17909
rect 9875 -17979 9887 -17943
rect 9921 -17979 9933 -17943
rect 9875 -18013 9933 -17979
rect 9875 -18049 9887 -18013
rect 9921 -18049 9933 -18013
rect 9875 -18061 9933 -18049
rect 10133 -17873 10191 -17861
rect 10133 -17909 10145 -17873
rect 10179 -17909 10191 -17873
rect 10133 -17943 10191 -17909
rect 10133 -17979 10145 -17943
rect 10179 -17979 10191 -17943
rect 10133 -18013 10191 -17979
rect 10133 -18049 10145 -18013
rect 10179 -18049 10191 -18013
rect 10133 -18061 10191 -18049
rect 10391 -17873 10449 -17861
rect 10391 -17909 10403 -17873
rect 10437 -17909 10449 -17873
rect 10391 -17943 10449 -17909
rect 10391 -17979 10403 -17943
rect 10437 -17979 10449 -17943
rect 10391 -18013 10449 -17979
rect 10391 -18049 10403 -18013
rect 10437 -18049 10449 -18013
rect 10391 -18061 10449 -18049
rect 10649 -17873 10707 -17861
rect 10649 -17909 10661 -17873
rect 10695 -17909 10707 -17873
rect 10649 -17943 10707 -17909
rect 10649 -17979 10661 -17943
rect 10695 -17979 10707 -17943
rect 10649 -18013 10707 -17979
rect 10649 -18049 10661 -18013
rect 10695 -18049 10707 -18013
rect 10649 -18061 10707 -18049
rect 10907 -17873 10965 -17861
rect 10907 -17909 10919 -17873
rect 10953 -17909 10965 -17873
rect 10907 -17943 10965 -17909
rect 10907 -17979 10919 -17943
rect 10953 -17979 10965 -17943
rect 10907 -18013 10965 -17979
rect 10907 -18049 10919 -18013
rect 10953 -18049 10965 -18013
rect 10907 -18061 10965 -18049
rect 11165 -17873 11223 -17861
rect 11165 -17909 11177 -17873
rect 11211 -17909 11223 -17873
rect 11165 -17943 11223 -17909
rect 11165 -17979 11177 -17943
rect 11211 -17979 11223 -17943
rect 11165 -18013 11223 -17979
rect 11165 -18049 11177 -18013
rect 11211 -18049 11223 -18013
rect 11165 -18061 11223 -18049
rect 11771 -17873 11829 -17861
rect 11771 -17909 11783 -17873
rect 11817 -17909 11829 -17873
rect 11771 -17943 11829 -17909
rect 11771 -17979 11783 -17943
rect 11817 -17979 11829 -17943
rect 11771 -18013 11829 -17979
rect 11771 -18049 11783 -18013
rect 11817 -18049 11829 -18013
rect 11771 -18061 11829 -18049
rect 12029 -17873 12087 -17861
rect 12029 -17909 12041 -17873
rect 12075 -17909 12087 -17873
rect 12029 -17943 12087 -17909
rect 12029 -17979 12041 -17943
rect 12075 -17979 12087 -17943
rect 12029 -18013 12087 -17979
rect 12029 -18049 12041 -18013
rect 12075 -18049 12087 -18013
rect 12029 -18061 12087 -18049
rect 12287 -17873 12345 -17861
rect 12287 -17909 12299 -17873
rect 12333 -17909 12345 -17873
rect 12287 -17943 12345 -17909
rect 12287 -17979 12299 -17943
rect 12333 -17979 12345 -17943
rect 12287 -18014 12345 -17979
rect 12287 -18050 12299 -18014
rect 12333 -18050 12345 -18014
rect 12287 -18061 12345 -18050
rect 12545 -17873 12603 -17861
rect 12545 -17909 12557 -17873
rect 12591 -17909 12603 -17873
rect 12545 -17943 12603 -17909
rect 12545 -17979 12557 -17943
rect 12591 -17979 12603 -17943
rect 12545 -18013 12603 -17979
rect 12545 -18049 12557 -18013
rect 12591 -18049 12603 -18013
rect 12545 -18061 12603 -18049
rect 12803 -17873 12861 -17861
rect 12803 -17909 12815 -17873
rect 12849 -17909 12861 -17873
rect 12803 -17943 12861 -17909
rect 12803 -17979 12815 -17943
rect 12849 -17979 12861 -17943
rect 12803 -18013 12861 -17979
rect 12803 -18049 12815 -18013
rect 12849 -18049 12861 -18013
rect 12803 -18061 12861 -18049
rect 13061 -17873 13119 -17861
rect 13061 -17909 13073 -17873
rect 13107 -17909 13119 -17873
rect 13061 -17943 13119 -17909
rect 13061 -17979 13073 -17943
rect 13107 -17979 13119 -17943
rect 13061 -18013 13119 -17979
rect 13061 -18049 13073 -18013
rect 13107 -18049 13119 -18013
rect 13061 -18061 13119 -18049
rect 13319 -17873 13377 -17861
rect 13319 -17909 13331 -17873
rect 13365 -17909 13377 -17873
rect 13319 -17943 13377 -17909
rect 13319 -17979 13331 -17943
rect 13365 -17979 13377 -17943
rect 13319 -18013 13377 -17979
rect 13319 -18049 13331 -18013
rect 13365 -18049 13377 -18013
rect 13319 -18061 13377 -18049
rect 13577 -17873 13635 -17861
rect 13577 -17909 13589 -17873
rect 13623 -17909 13635 -17873
rect 13577 -17943 13635 -17909
rect 13577 -17979 13589 -17943
rect 13623 -17979 13635 -17943
rect 13577 -18013 13635 -17979
rect 13577 -18049 13589 -18013
rect 13623 -18049 13635 -18013
rect 13577 -18061 13635 -18049
rect 13835 -17873 13893 -17861
rect 13835 -17909 13847 -17873
rect 13881 -17909 13893 -17873
rect 13835 -17943 13893 -17909
rect 13835 -17979 13847 -17943
rect 13881 -17979 13893 -17943
rect 13835 -18013 13893 -17979
rect 13835 -18049 13847 -18013
rect 13881 -18049 13893 -18013
rect 13835 -18061 13893 -18049
rect 14434 -17872 14492 -17860
rect 14434 -17908 14446 -17872
rect 14480 -17908 14492 -17872
rect 14434 -17942 14492 -17908
rect 14434 -17978 14446 -17942
rect 14480 -17978 14492 -17942
rect 14434 -18012 14492 -17978
rect 14434 -18048 14446 -18012
rect 14480 -18048 14492 -18012
rect 14434 -18060 14492 -18048
rect 14692 -17872 14750 -17860
rect 14692 -17908 14704 -17872
rect 14738 -17908 14750 -17872
rect 14692 -17942 14750 -17908
rect 14692 -17978 14704 -17942
rect 14738 -17978 14750 -17942
rect 14692 -18012 14750 -17978
rect 14692 -18048 14704 -18012
rect 14738 -18048 14750 -18012
rect 14692 -18060 14750 -18048
rect 14950 -17872 15008 -17860
rect 14950 -17908 14962 -17872
rect 14996 -17908 15008 -17872
rect 14950 -17942 15008 -17908
rect 14950 -17978 14962 -17942
rect 14996 -17978 15008 -17942
rect 14950 -18013 15008 -17978
rect 14950 -18049 14962 -18013
rect 14996 -18049 15008 -18013
rect 14950 -18060 15008 -18049
rect 15208 -17872 15266 -17860
rect 15208 -17908 15220 -17872
rect 15254 -17908 15266 -17872
rect 15208 -17942 15266 -17908
rect 15208 -17978 15220 -17942
rect 15254 -17978 15266 -17942
rect 15208 -18012 15266 -17978
rect 15208 -18048 15220 -18012
rect 15254 -18048 15266 -18012
rect 15208 -18060 15266 -18048
rect 15466 -17872 15524 -17860
rect 15466 -17908 15478 -17872
rect 15512 -17908 15524 -17872
rect 15466 -17942 15524 -17908
rect 15466 -17978 15478 -17942
rect 15512 -17978 15524 -17942
rect 15466 -18012 15524 -17978
rect 15466 -18048 15478 -18012
rect 15512 -18048 15524 -18012
rect 15466 -18060 15524 -18048
rect 15724 -17872 15782 -17860
rect 15724 -17908 15736 -17872
rect 15770 -17908 15782 -17872
rect 15724 -17942 15782 -17908
rect 15724 -17978 15736 -17942
rect 15770 -17978 15782 -17942
rect 15724 -18012 15782 -17978
rect 15724 -18048 15736 -18012
rect 15770 -18048 15782 -18012
rect 15724 -18060 15782 -18048
rect 15982 -17872 16040 -17860
rect 15982 -17908 15994 -17872
rect 16028 -17908 16040 -17872
rect 15982 -17942 16040 -17908
rect 15982 -17978 15994 -17942
rect 16028 -17978 16040 -17942
rect 15982 -18012 16040 -17978
rect 15982 -18048 15994 -18012
rect 16028 -18048 16040 -18012
rect 15982 -18060 16040 -18048
rect 16240 -17872 16298 -17860
rect 16240 -17908 16252 -17872
rect 16286 -17908 16298 -17872
rect 16240 -17942 16298 -17908
rect 16240 -17978 16252 -17942
rect 16286 -17978 16298 -17942
rect 16240 -18012 16298 -17978
rect 16240 -18048 16252 -18012
rect 16286 -18048 16298 -18012
rect 16240 -18060 16298 -18048
rect 16498 -17872 16556 -17860
rect 16498 -17908 16510 -17872
rect 16544 -17908 16556 -17872
rect 16498 -17942 16556 -17908
rect 16498 -17978 16510 -17942
rect 16544 -17978 16556 -17942
rect 16498 -18012 16556 -17978
rect 16498 -18048 16510 -18012
rect 16544 -18048 16556 -18012
rect 16498 -18060 16556 -18048
rect 8981 -18527 9039 -18513
rect 8981 -18561 8993 -18527
rect 9027 -18561 9039 -18527
rect 8981 -18595 9039 -18561
rect 8981 -18631 8993 -18595
rect 9027 -18631 9039 -18595
rect 8981 -18665 9039 -18631
rect 8981 -18699 8993 -18665
rect 9027 -18699 9039 -18665
rect 8981 -18713 9039 -18699
rect 9239 -18527 9297 -18513
rect 9239 -18561 9251 -18527
rect 9285 -18561 9297 -18527
rect 9239 -18595 9297 -18561
rect 9239 -18631 9251 -18595
rect 9285 -18631 9297 -18595
rect 9239 -18665 9297 -18631
rect 9239 -18699 9251 -18665
rect 9285 -18699 9297 -18665
rect 9239 -18713 9297 -18699
rect 9521 -18527 9579 -18513
rect 9521 -18561 9533 -18527
rect 9567 -18561 9579 -18527
rect 9521 -18595 9579 -18561
rect 9521 -18631 9533 -18595
rect 9567 -18631 9579 -18595
rect 9521 -18665 9579 -18631
rect 9521 -18699 9533 -18665
rect 9567 -18699 9579 -18665
rect 9521 -18713 9579 -18699
rect 9779 -18527 9837 -18513
rect 9779 -18561 9791 -18527
rect 9825 -18561 9837 -18527
rect 9779 -18595 9837 -18561
rect 9779 -18631 9791 -18595
rect 9825 -18631 9837 -18595
rect 9779 -18665 9837 -18631
rect 9779 -18699 9791 -18665
rect 9825 -18699 9837 -18665
rect 9779 -18713 9837 -18699
rect 10001 -18527 10059 -18513
rect 10001 -18561 10013 -18527
rect 10047 -18561 10059 -18527
rect 10001 -18595 10059 -18561
rect 10001 -18631 10013 -18595
rect 10047 -18631 10059 -18595
rect 10001 -18665 10059 -18631
rect 10001 -18699 10013 -18665
rect 10047 -18699 10059 -18665
rect 10001 -18713 10059 -18699
rect 10259 -18527 10317 -18513
rect 10259 -18561 10271 -18527
rect 10305 -18561 10317 -18527
rect 10259 -18595 10317 -18561
rect 10259 -18631 10271 -18595
rect 10305 -18631 10317 -18595
rect 10259 -18665 10317 -18631
rect 10259 -18699 10271 -18665
rect 10305 -18699 10317 -18665
rect 10259 -18713 10317 -18699
rect 10504 -18525 10562 -18511
rect 10504 -18559 10516 -18525
rect 10550 -18559 10562 -18525
rect 10504 -18593 10562 -18559
rect 10504 -18629 10516 -18593
rect 10550 -18629 10562 -18593
rect 10504 -18663 10562 -18629
rect 10504 -18697 10516 -18663
rect 10550 -18697 10562 -18663
rect 10504 -18711 10562 -18697
rect 10762 -18525 10820 -18511
rect 10762 -18559 10774 -18525
rect 10808 -18559 10820 -18525
rect 10762 -18593 10820 -18559
rect 10762 -18629 10774 -18593
rect 10808 -18629 10820 -18593
rect 10762 -18663 10820 -18629
rect 10762 -18697 10774 -18663
rect 10808 -18697 10820 -18663
rect 10762 -18711 10820 -18697
rect 11014 -18515 11072 -18501
rect 11014 -18549 11026 -18515
rect 11060 -18549 11072 -18515
rect 11014 -18583 11072 -18549
rect 11014 -18619 11026 -18583
rect 11060 -18619 11072 -18583
rect 11014 -18653 11072 -18619
rect 11014 -18687 11026 -18653
rect 11060 -18687 11072 -18653
rect 11014 -18701 11072 -18687
rect 11272 -18515 11330 -18501
rect 11272 -18549 11284 -18515
rect 11318 -18549 11330 -18515
rect 11272 -18583 11330 -18549
rect 11272 -18619 11284 -18583
rect 11318 -18619 11330 -18583
rect 11272 -18653 11330 -18619
rect 11272 -18687 11284 -18653
rect 11318 -18687 11330 -18653
rect 11272 -18701 11330 -18687
rect 11651 -18527 11709 -18513
rect 11651 -18561 11663 -18527
rect 11697 -18561 11709 -18527
rect 11651 -18595 11709 -18561
rect 11651 -18631 11663 -18595
rect 11697 -18631 11709 -18595
rect 11651 -18665 11709 -18631
rect 11651 -18699 11663 -18665
rect 11697 -18699 11709 -18665
rect 11651 -18713 11709 -18699
rect 11909 -18527 11967 -18513
rect 11909 -18561 11921 -18527
rect 11955 -18561 11967 -18527
rect 11909 -18595 11967 -18561
rect 11909 -18631 11921 -18595
rect 11955 -18631 11967 -18595
rect 11909 -18665 11967 -18631
rect 11909 -18699 11921 -18665
rect 11955 -18699 11967 -18665
rect 11909 -18713 11967 -18699
rect 12191 -18527 12249 -18513
rect 12191 -18561 12203 -18527
rect 12237 -18561 12249 -18527
rect 12191 -18595 12249 -18561
rect 12191 -18631 12203 -18595
rect 12237 -18631 12249 -18595
rect 12191 -18665 12249 -18631
rect 12191 -18699 12203 -18665
rect 12237 -18699 12249 -18665
rect 12191 -18713 12249 -18699
rect 12449 -18527 12507 -18513
rect 12449 -18561 12461 -18527
rect 12495 -18561 12507 -18527
rect 12449 -18595 12507 -18561
rect 12449 -18631 12461 -18595
rect 12495 -18631 12507 -18595
rect 12449 -18665 12507 -18631
rect 12449 -18699 12461 -18665
rect 12495 -18699 12507 -18665
rect 12449 -18713 12507 -18699
rect 12671 -18527 12729 -18513
rect 12671 -18561 12683 -18527
rect 12717 -18561 12729 -18527
rect 12671 -18595 12729 -18561
rect 12671 -18631 12683 -18595
rect 12717 -18631 12729 -18595
rect 12671 -18665 12729 -18631
rect 12671 -18699 12683 -18665
rect 12717 -18699 12729 -18665
rect 12671 -18713 12729 -18699
rect 12929 -18527 12987 -18513
rect 12929 -18561 12941 -18527
rect 12975 -18561 12987 -18527
rect 12929 -18595 12987 -18561
rect 12929 -18631 12941 -18595
rect 12975 -18631 12987 -18595
rect 12929 -18665 12987 -18631
rect 12929 -18699 12941 -18665
rect 12975 -18699 12987 -18665
rect 12929 -18713 12987 -18699
rect 13174 -18525 13232 -18511
rect 13174 -18559 13186 -18525
rect 13220 -18559 13232 -18525
rect 13174 -18593 13232 -18559
rect 13174 -18629 13186 -18593
rect 13220 -18629 13232 -18593
rect 13174 -18663 13232 -18629
rect 13174 -18697 13186 -18663
rect 13220 -18697 13232 -18663
rect 13174 -18711 13232 -18697
rect 13432 -18525 13490 -18511
rect 13432 -18559 13444 -18525
rect 13478 -18559 13490 -18525
rect 13432 -18593 13490 -18559
rect 13432 -18629 13444 -18593
rect 13478 -18629 13490 -18593
rect 13432 -18663 13490 -18629
rect 13432 -18697 13444 -18663
rect 13478 -18697 13490 -18663
rect 13432 -18711 13490 -18697
rect 13684 -18515 13742 -18501
rect 13684 -18549 13696 -18515
rect 13730 -18549 13742 -18515
rect 13684 -18583 13742 -18549
rect 13684 -18619 13696 -18583
rect 13730 -18619 13742 -18583
rect 13684 -18653 13742 -18619
rect 13684 -18687 13696 -18653
rect 13730 -18687 13742 -18653
rect 13684 -18701 13742 -18687
rect 13942 -18515 14000 -18501
rect 13942 -18549 13954 -18515
rect 13988 -18549 14000 -18515
rect 13942 -18583 14000 -18549
rect 13942 -18619 13954 -18583
rect 13988 -18619 14000 -18583
rect 13942 -18653 14000 -18619
rect 13942 -18687 13954 -18653
rect 13988 -18687 14000 -18653
rect 13942 -18701 14000 -18687
rect 14314 -18526 14372 -18512
rect 14314 -18560 14326 -18526
rect 14360 -18560 14372 -18526
rect 14314 -18594 14372 -18560
rect 14314 -18630 14326 -18594
rect 14360 -18630 14372 -18594
rect 14314 -18664 14372 -18630
rect 14314 -18698 14326 -18664
rect 14360 -18698 14372 -18664
rect 14314 -18712 14372 -18698
rect 14572 -18526 14630 -18512
rect 14572 -18560 14584 -18526
rect 14618 -18560 14630 -18526
rect 14572 -18594 14630 -18560
rect 14572 -18630 14584 -18594
rect 14618 -18630 14630 -18594
rect 14572 -18664 14630 -18630
rect 14572 -18698 14584 -18664
rect 14618 -18698 14630 -18664
rect 14572 -18712 14630 -18698
rect 14854 -18526 14912 -18512
rect 14854 -18560 14866 -18526
rect 14900 -18560 14912 -18526
rect 14854 -18594 14912 -18560
rect 14854 -18630 14866 -18594
rect 14900 -18630 14912 -18594
rect 14854 -18664 14912 -18630
rect 14854 -18698 14866 -18664
rect 14900 -18698 14912 -18664
rect 14854 -18712 14912 -18698
rect 15112 -18526 15170 -18512
rect 15112 -18560 15124 -18526
rect 15158 -18560 15170 -18526
rect 15112 -18594 15170 -18560
rect 15112 -18630 15124 -18594
rect 15158 -18630 15170 -18594
rect 15112 -18664 15170 -18630
rect 15112 -18698 15124 -18664
rect 15158 -18698 15170 -18664
rect 15112 -18712 15170 -18698
rect 15334 -18526 15392 -18512
rect 15334 -18560 15346 -18526
rect 15380 -18560 15392 -18526
rect 15334 -18594 15392 -18560
rect 15334 -18630 15346 -18594
rect 15380 -18630 15392 -18594
rect 15334 -18664 15392 -18630
rect 15334 -18698 15346 -18664
rect 15380 -18698 15392 -18664
rect 15334 -18712 15392 -18698
rect 15592 -18526 15650 -18512
rect 15592 -18560 15604 -18526
rect 15638 -18560 15650 -18526
rect 15592 -18594 15650 -18560
rect 15592 -18630 15604 -18594
rect 15638 -18630 15650 -18594
rect 15592 -18664 15650 -18630
rect 15592 -18698 15604 -18664
rect 15638 -18698 15650 -18664
rect 15592 -18712 15650 -18698
rect 15837 -18524 15895 -18510
rect 15837 -18558 15849 -18524
rect 15883 -18558 15895 -18524
rect 15837 -18592 15895 -18558
rect 15837 -18628 15849 -18592
rect 15883 -18628 15895 -18592
rect 15837 -18662 15895 -18628
rect 15837 -18696 15849 -18662
rect 15883 -18696 15895 -18662
rect 15837 -18710 15895 -18696
rect 16095 -18524 16153 -18510
rect 16095 -18558 16107 -18524
rect 16141 -18558 16153 -18524
rect 16095 -18592 16153 -18558
rect 16095 -18628 16107 -18592
rect 16141 -18628 16153 -18592
rect 16095 -18662 16153 -18628
rect 16095 -18696 16107 -18662
rect 16141 -18696 16153 -18662
rect 16095 -18710 16153 -18696
rect 16347 -18514 16405 -18500
rect 16347 -18548 16359 -18514
rect 16393 -18548 16405 -18514
rect 16347 -18582 16405 -18548
rect 16347 -18618 16359 -18582
rect 16393 -18618 16405 -18582
rect 16347 -18652 16405 -18618
rect 16347 -18686 16359 -18652
rect 16393 -18686 16405 -18652
rect 16347 -18700 16405 -18686
rect 16605 -18514 16663 -18500
rect 16605 -18548 16617 -18514
rect 16651 -18548 16663 -18514
rect 16605 -18582 16663 -18548
rect 16605 -18618 16617 -18582
rect 16651 -18618 16663 -18582
rect 16605 -18652 16663 -18618
rect 16605 -18686 16617 -18652
rect 16651 -18686 16663 -18652
rect 16605 -18700 16663 -18686
rect 16646 -20421 16704 -20409
rect 16646 -20481 16658 -20421
rect 16692 -20481 16704 -20421
rect 16646 -20493 16704 -20481
rect 16734 -20421 16792 -20409
rect 16734 -20481 16746 -20421
rect 16780 -20481 16792 -20421
rect 16734 -20493 16792 -20481
rect 17036 -20421 17094 -20409
rect 17036 -20481 17048 -20421
rect 17082 -20481 17094 -20421
rect 17036 -20493 17094 -20481
rect 17124 -20421 17182 -20409
rect 17124 -20481 17136 -20421
rect 17170 -20481 17182 -20421
rect 17124 -20493 17182 -20481
rect 9101 -21269 9159 -21257
rect 9101 -21305 9113 -21269
rect 9147 -21305 9159 -21269
rect 9101 -21339 9159 -21305
rect 9101 -21375 9113 -21339
rect 9147 -21375 9159 -21339
rect 9101 -21409 9159 -21375
rect 9101 -21445 9113 -21409
rect 9147 -21445 9159 -21409
rect 9101 -21457 9159 -21445
rect 9359 -21269 9417 -21257
rect 9359 -21305 9371 -21269
rect 9405 -21305 9417 -21269
rect 9359 -21339 9417 -21305
rect 9359 -21375 9371 -21339
rect 9405 -21375 9417 -21339
rect 9359 -21409 9417 -21375
rect 9359 -21445 9371 -21409
rect 9405 -21445 9417 -21409
rect 9359 -21457 9417 -21445
rect 9617 -21269 9675 -21257
rect 9617 -21305 9629 -21269
rect 9663 -21305 9675 -21269
rect 9617 -21339 9675 -21305
rect 9617 -21375 9629 -21339
rect 9663 -21375 9675 -21339
rect 9617 -21410 9675 -21375
rect 9617 -21446 9629 -21410
rect 9663 -21446 9675 -21410
rect 9617 -21457 9675 -21446
rect 9875 -21269 9933 -21257
rect 9875 -21305 9887 -21269
rect 9921 -21305 9933 -21269
rect 9875 -21339 9933 -21305
rect 9875 -21375 9887 -21339
rect 9921 -21375 9933 -21339
rect 9875 -21409 9933 -21375
rect 9875 -21445 9887 -21409
rect 9921 -21445 9933 -21409
rect 9875 -21457 9933 -21445
rect 10133 -21269 10191 -21257
rect 10133 -21305 10145 -21269
rect 10179 -21305 10191 -21269
rect 10133 -21339 10191 -21305
rect 10133 -21375 10145 -21339
rect 10179 -21375 10191 -21339
rect 10133 -21409 10191 -21375
rect 10133 -21445 10145 -21409
rect 10179 -21445 10191 -21409
rect 10133 -21457 10191 -21445
rect 10391 -21269 10449 -21257
rect 10391 -21305 10403 -21269
rect 10437 -21305 10449 -21269
rect 10391 -21339 10449 -21305
rect 10391 -21375 10403 -21339
rect 10437 -21375 10449 -21339
rect 10391 -21409 10449 -21375
rect 10391 -21445 10403 -21409
rect 10437 -21445 10449 -21409
rect 10391 -21457 10449 -21445
rect 10649 -21269 10707 -21257
rect 10649 -21305 10661 -21269
rect 10695 -21305 10707 -21269
rect 10649 -21339 10707 -21305
rect 10649 -21375 10661 -21339
rect 10695 -21375 10707 -21339
rect 10649 -21409 10707 -21375
rect 10649 -21445 10661 -21409
rect 10695 -21445 10707 -21409
rect 10649 -21457 10707 -21445
rect 10907 -21269 10965 -21257
rect 10907 -21305 10919 -21269
rect 10953 -21305 10965 -21269
rect 10907 -21339 10965 -21305
rect 10907 -21375 10919 -21339
rect 10953 -21375 10965 -21339
rect 10907 -21409 10965 -21375
rect 10907 -21445 10919 -21409
rect 10953 -21445 10965 -21409
rect 10907 -21457 10965 -21445
rect 11165 -21269 11223 -21257
rect 11165 -21305 11177 -21269
rect 11211 -21305 11223 -21269
rect 11165 -21339 11223 -21305
rect 11165 -21375 11177 -21339
rect 11211 -21375 11223 -21339
rect 11165 -21409 11223 -21375
rect 11165 -21445 11177 -21409
rect 11211 -21445 11223 -21409
rect 11165 -21457 11223 -21445
rect 11771 -21269 11829 -21257
rect 11771 -21305 11783 -21269
rect 11817 -21305 11829 -21269
rect 11771 -21339 11829 -21305
rect 11771 -21375 11783 -21339
rect 11817 -21375 11829 -21339
rect 11771 -21409 11829 -21375
rect 11771 -21445 11783 -21409
rect 11817 -21445 11829 -21409
rect 11771 -21457 11829 -21445
rect 12029 -21269 12087 -21257
rect 12029 -21305 12041 -21269
rect 12075 -21305 12087 -21269
rect 12029 -21339 12087 -21305
rect 12029 -21375 12041 -21339
rect 12075 -21375 12087 -21339
rect 12029 -21409 12087 -21375
rect 12029 -21445 12041 -21409
rect 12075 -21445 12087 -21409
rect 12029 -21457 12087 -21445
rect 12287 -21269 12345 -21257
rect 12287 -21305 12299 -21269
rect 12333 -21305 12345 -21269
rect 12287 -21339 12345 -21305
rect 12287 -21375 12299 -21339
rect 12333 -21375 12345 -21339
rect 12287 -21410 12345 -21375
rect 12287 -21446 12299 -21410
rect 12333 -21446 12345 -21410
rect 12287 -21457 12345 -21446
rect 12545 -21269 12603 -21257
rect 12545 -21305 12557 -21269
rect 12591 -21305 12603 -21269
rect 12545 -21339 12603 -21305
rect 12545 -21375 12557 -21339
rect 12591 -21375 12603 -21339
rect 12545 -21409 12603 -21375
rect 12545 -21445 12557 -21409
rect 12591 -21445 12603 -21409
rect 12545 -21457 12603 -21445
rect 12803 -21269 12861 -21257
rect 12803 -21305 12815 -21269
rect 12849 -21305 12861 -21269
rect 12803 -21339 12861 -21305
rect 12803 -21375 12815 -21339
rect 12849 -21375 12861 -21339
rect 12803 -21409 12861 -21375
rect 12803 -21445 12815 -21409
rect 12849 -21445 12861 -21409
rect 12803 -21457 12861 -21445
rect 13061 -21269 13119 -21257
rect 13061 -21305 13073 -21269
rect 13107 -21305 13119 -21269
rect 13061 -21339 13119 -21305
rect 13061 -21375 13073 -21339
rect 13107 -21375 13119 -21339
rect 13061 -21409 13119 -21375
rect 13061 -21445 13073 -21409
rect 13107 -21445 13119 -21409
rect 13061 -21457 13119 -21445
rect 13319 -21269 13377 -21257
rect 13319 -21305 13331 -21269
rect 13365 -21305 13377 -21269
rect 13319 -21339 13377 -21305
rect 13319 -21375 13331 -21339
rect 13365 -21375 13377 -21339
rect 13319 -21409 13377 -21375
rect 13319 -21445 13331 -21409
rect 13365 -21445 13377 -21409
rect 13319 -21457 13377 -21445
rect 13577 -21269 13635 -21257
rect 13577 -21305 13589 -21269
rect 13623 -21305 13635 -21269
rect 13577 -21339 13635 -21305
rect 13577 -21375 13589 -21339
rect 13623 -21375 13635 -21339
rect 13577 -21409 13635 -21375
rect 13577 -21445 13589 -21409
rect 13623 -21445 13635 -21409
rect 13577 -21457 13635 -21445
rect 13835 -21269 13893 -21257
rect 13835 -21305 13847 -21269
rect 13881 -21305 13893 -21269
rect 13835 -21339 13893 -21305
rect 13835 -21375 13847 -21339
rect 13881 -21375 13893 -21339
rect 13835 -21409 13893 -21375
rect 13835 -21445 13847 -21409
rect 13881 -21445 13893 -21409
rect 13835 -21457 13893 -21445
rect 14434 -21268 14492 -21256
rect 14434 -21304 14446 -21268
rect 14480 -21304 14492 -21268
rect 14434 -21338 14492 -21304
rect 14434 -21374 14446 -21338
rect 14480 -21374 14492 -21338
rect 14434 -21408 14492 -21374
rect 14434 -21444 14446 -21408
rect 14480 -21444 14492 -21408
rect 14434 -21456 14492 -21444
rect 14692 -21268 14750 -21256
rect 14692 -21304 14704 -21268
rect 14738 -21304 14750 -21268
rect 14692 -21338 14750 -21304
rect 14692 -21374 14704 -21338
rect 14738 -21374 14750 -21338
rect 14692 -21408 14750 -21374
rect 14692 -21444 14704 -21408
rect 14738 -21444 14750 -21408
rect 14692 -21456 14750 -21444
rect 14950 -21268 15008 -21256
rect 14950 -21304 14962 -21268
rect 14996 -21304 15008 -21268
rect 14950 -21338 15008 -21304
rect 14950 -21374 14962 -21338
rect 14996 -21374 15008 -21338
rect 14950 -21409 15008 -21374
rect 14950 -21445 14962 -21409
rect 14996 -21445 15008 -21409
rect 14950 -21456 15008 -21445
rect 15208 -21268 15266 -21256
rect 15208 -21304 15220 -21268
rect 15254 -21304 15266 -21268
rect 15208 -21338 15266 -21304
rect 15208 -21374 15220 -21338
rect 15254 -21374 15266 -21338
rect 15208 -21408 15266 -21374
rect 15208 -21444 15220 -21408
rect 15254 -21444 15266 -21408
rect 15208 -21456 15266 -21444
rect 15466 -21268 15524 -21256
rect 15466 -21304 15478 -21268
rect 15512 -21304 15524 -21268
rect 15466 -21338 15524 -21304
rect 15466 -21374 15478 -21338
rect 15512 -21374 15524 -21338
rect 15466 -21408 15524 -21374
rect 15466 -21444 15478 -21408
rect 15512 -21444 15524 -21408
rect 15466 -21456 15524 -21444
rect 15724 -21268 15782 -21256
rect 15724 -21304 15736 -21268
rect 15770 -21304 15782 -21268
rect 15724 -21338 15782 -21304
rect 15724 -21374 15736 -21338
rect 15770 -21374 15782 -21338
rect 15724 -21408 15782 -21374
rect 15724 -21444 15736 -21408
rect 15770 -21444 15782 -21408
rect 15724 -21456 15782 -21444
rect 15982 -21268 16040 -21256
rect 15982 -21304 15994 -21268
rect 16028 -21304 16040 -21268
rect 15982 -21338 16040 -21304
rect 15982 -21374 15994 -21338
rect 16028 -21374 16040 -21338
rect 15982 -21408 16040 -21374
rect 15982 -21444 15994 -21408
rect 16028 -21444 16040 -21408
rect 15982 -21456 16040 -21444
rect 16240 -21268 16298 -21256
rect 16240 -21304 16252 -21268
rect 16286 -21304 16298 -21268
rect 16240 -21338 16298 -21304
rect 16240 -21374 16252 -21338
rect 16286 -21374 16298 -21338
rect 16240 -21408 16298 -21374
rect 16240 -21444 16252 -21408
rect 16286 -21444 16298 -21408
rect 16240 -21456 16298 -21444
rect 16498 -21268 16556 -21256
rect 16498 -21304 16510 -21268
rect 16544 -21304 16556 -21268
rect 16498 -21338 16556 -21304
rect 16498 -21374 16510 -21338
rect 16544 -21374 16556 -21338
rect 16498 -21408 16556 -21374
rect 16498 -21444 16510 -21408
rect 16544 -21444 16556 -21408
rect 16498 -21456 16556 -21444
rect 9101 -21687 9159 -21675
rect 9101 -21723 9113 -21687
rect 9147 -21723 9159 -21687
rect 9101 -21757 9159 -21723
rect 9101 -21793 9113 -21757
rect 9147 -21793 9159 -21757
rect 9101 -21827 9159 -21793
rect 9101 -21863 9113 -21827
rect 9147 -21863 9159 -21827
rect 9101 -21875 9159 -21863
rect 9359 -21687 9417 -21675
rect 9359 -21723 9371 -21687
rect 9405 -21723 9417 -21687
rect 9359 -21757 9417 -21723
rect 9359 -21793 9371 -21757
rect 9405 -21793 9417 -21757
rect 9359 -21827 9417 -21793
rect 9359 -21863 9371 -21827
rect 9405 -21863 9417 -21827
rect 9359 -21875 9417 -21863
rect 9617 -21687 9675 -21675
rect 9617 -21723 9629 -21687
rect 9663 -21723 9675 -21687
rect 9617 -21757 9675 -21723
rect 9617 -21793 9629 -21757
rect 9663 -21793 9675 -21757
rect 9617 -21828 9675 -21793
rect 9617 -21864 9629 -21828
rect 9663 -21864 9675 -21828
rect 9617 -21875 9675 -21864
rect 9875 -21687 9933 -21675
rect 9875 -21723 9887 -21687
rect 9921 -21723 9933 -21687
rect 9875 -21757 9933 -21723
rect 9875 -21793 9887 -21757
rect 9921 -21793 9933 -21757
rect 9875 -21827 9933 -21793
rect 9875 -21863 9887 -21827
rect 9921 -21863 9933 -21827
rect 9875 -21875 9933 -21863
rect 10133 -21687 10191 -21675
rect 10133 -21723 10145 -21687
rect 10179 -21723 10191 -21687
rect 10133 -21757 10191 -21723
rect 10133 -21793 10145 -21757
rect 10179 -21793 10191 -21757
rect 10133 -21827 10191 -21793
rect 10133 -21863 10145 -21827
rect 10179 -21863 10191 -21827
rect 10133 -21875 10191 -21863
rect 10391 -21687 10449 -21675
rect 10391 -21723 10403 -21687
rect 10437 -21723 10449 -21687
rect 10391 -21757 10449 -21723
rect 10391 -21793 10403 -21757
rect 10437 -21793 10449 -21757
rect 10391 -21827 10449 -21793
rect 10391 -21863 10403 -21827
rect 10437 -21863 10449 -21827
rect 10391 -21875 10449 -21863
rect 10649 -21687 10707 -21675
rect 10649 -21723 10661 -21687
rect 10695 -21723 10707 -21687
rect 10649 -21757 10707 -21723
rect 10649 -21793 10661 -21757
rect 10695 -21793 10707 -21757
rect 10649 -21827 10707 -21793
rect 10649 -21863 10661 -21827
rect 10695 -21863 10707 -21827
rect 10649 -21875 10707 -21863
rect 10907 -21687 10965 -21675
rect 10907 -21723 10919 -21687
rect 10953 -21723 10965 -21687
rect 10907 -21757 10965 -21723
rect 10907 -21793 10919 -21757
rect 10953 -21793 10965 -21757
rect 10907 -21827 10965 -21793
rect 10907 -21863 10919 -21827
rect 10953 -21863 10965 -21827
rect 10907 -21875 10965 -21863
rect 11165 -21687 11223 -21675
rect 11165 -21723 11177 -21687
rect 11211 -21723 11223 -21687
rect 11165 -21757 11223 -21723
rect 11165 -21793 11177 -21757
rect 11211 -21793 11223 -21757
rect 11165 -21827 11223 -21793
rect 11165 -21863 11177 -21827
rect 11211 -21863 11223 -21827
rect 11165 -21875 11223 -21863
rect 11771 -21687 11829 -21675
rect 11771 -21723 11783 -21687
rect 11817 -21723 11829 -21687
rect 11771 -21757 11829 -21723
rect 11771 -21793 11783 -21757
rect 11817 -21793 11829 -21757
rect 11771 -21827 11829 -21793
rect 11771 -21863 11783 -21827
rect 11817 -21863 11829 -21827
rect 11771 -21875 11829 -21863
rect 12029 -21687 12087 -21675
rect 12029 -21723 12041 -21687
rect 12075 -21723 12087 -21687
rect 12029 -21757 12087 -21723
rect 12029 -21793 12041 -21757
rect 12075 -21793 12087 -21757
rect 12029 -21827 12087 -21793
rect 12029 -21863 12041 -21827
rect 12075 -21863 12087 -21827
rect 12029 -21875 12087 -21863
rect 12287 -21687 12345 -21675
rect 12287 -21723 12299 -21687
rect 12333 -21723 12345 -21687
rect 12287 -21757 12345 -21723
rect 12287 -21793 12299 -21757
rect 12333 -21793 12345 -21757
rect 12287 -21828 12345 -21793
rect 12287 -21864 12299 -21828
rect 12333 -21864 12345 -21828
rect 12287 -21875 12345 -21864
rect 12545 -21687 12603 -21675
rect 12545 -21723 12557 -21687
rect 12591 -21723 12603 -21687
rect 12545 -21757 12603 -21723
rect 12545 -21793 12557 -21757
rect 12591 -21793 12603 -21757
rect 12545 -21827 12603 -21793
rect 12545 -21863 12557 -21827
rect 12591 -21863 12603 -21827
rect 12545 -21875 12603 -21863
rect 12803 -21687 12861 -21675
rect 12803 -21723 12815 -21687
rect 12849 -21723 12861 -21687
rect 12803 -21757 12861 -21723
rect 12803 -21793 12815 -21757
rect 12849 -21793 12861 -21757
rect 12803 -21827 12861 -21793
rect 12803 -21863 12815 -21827
rect 12849 -21863 12861 -21827
rect 12803 -21875 12861 -21863
rect 13061 -21687 13119 -21675
rect 13061 -21723 13073 -21687
rect 13107 -21723 13119 -21687
rect 13061 -21757 13119 -21723
rect 13061 -21793 13073 -21757
rect 13107 -21793 13119 -21757
rect 13061 -21827 13119 -21793
rect 13061 -21863 13073 -21827
rect 13107 -21863 13119 -21827
rect 13061 -21875 13119 -21863
rect 13319 -21687 13377 -21675
rect 13319 -21723 13331 -21687
rect 13365 -21723 13377 -21687
rect 13319 -21757 13377 -21723
rect 13319 -21793 13331 -21757
rect 13365 -21793 13377 -21757
rect 13319 -21827 13377 -21793
rect 13319 -21863 13331 -21827
rect 13365 -21863 13377 -21827
rect 13319 -21875 13377 -21863
rect 13577 -21687 13635 -21675
rect 13577 -21723 13589 -21687
rect 13623 -21723 13635 -21687
rect 13577 -21757 13635 -21723
rect 13577 -21793 13589 -21757
rect 13623 -21793 13635 -21757
rect 13577 -21827 13635 -21793
rect 13577 -21863 13589 -21827
rect 13623 -21863 13635 -21827
rect 13577 -21875 13635 -21863
rect 13835 -21687 13893 -21675
rect 13835 -21723 13847 -21687
rect 13881 -21723 13893 -21687
rect 13835 -21757 13893 -21723
rect 13835 -21793 13847 -21757
rect 13881 -21793 13893 -21757
rect 13835 -21827 13893 -21793
rect 13835 -21863 13847 -21827
rect 13881 -21863 13893 -21827
rect 13835 -21875 13893 -21863
rect 14434 -21686 14492 -21674
rect 14434 -21722 14446 -21686
rect 14480 -21722 14492 -21686
rect 14434 -21756 14492 -21722
rect 14434 -21792 14446 -21756
rect 14480 -21792 14492 -21756
rect 14434 -21826 14492 -21792
rect 14434 -21862 14446 -21826
rect 14480 -21862 14492 -21826
rect 14434 -21874 14492 -21862
rect 14692 -21686 14750 -21674
rect 14692 -21722 14704 -21686
rect 14738 -21722 14750 -21686
rect 14692 -21756 14750 -21722
rect 14692 -21792 14704 -21756
rect 14738 -21792 14750 -21756
rect 14692 -21826 14750 -21792
rect 14692 -21862 14704 -21826
rect 14738 -21862 14750 -21826
rect 14692 -21874 14750 -21862
rect 14950 -21686 15008 -21674
rect 14950 -21722 14962 -21686
rect 14996 -21722 15008 -21686
rect 14950 -21756 15008 -21722
rect 14950 -21792 14962 -21756
rect 14996 -21792 15008 -21756
rect 14950 -21827 15008 -21792
rect 14950 -21863 14962 -21827
rect 14996 -21863 15008 -21827
rect 14950 -21874 15008 -21863
rect 15208 -21686 15266 -21674
rect 15208 -21722 15220 -21686
rect 15254 -21722 15266 -21686
rect 15208 -21756 15266 -21722
rect 15208 -21792 15220 -21756
rect 15254 -21792 15266 -21756
rect 15208 -21826 15266 -21792
rect 15208 -21862 15220 -21826
rect 15254 -21862 15266 -21826
rect 15208 -21874 15266 -21862
rect 15466 -21686 15524 -21674
rect 15466 -21722 15478 -21686
rect 15512 -21722 15524 -21686
rect 15466 -21756 15524 -21722
rect 15466 -21792 15478 -21756
rect 15512 -21792 15524 -21756
rect 15466 -21826 15524 -21792
rect 15466 -21862 15478 -21826
rect 15512 -21862 15524 -21826
rect 15466 -21874 15524 -21862
rect 15724 -21686 15782 -21674
rect 15724 -21722 15736 -21686
rect 15770 -21722 15782 -21686
rect 15724 -21756 15782 -21722
rect 15724 -21792 15736 -21756
rect 15770 -21792 15782 -21756
rect 15724 -21826 15782 -21792
rect 15724 -21862 15736 -21826
rect 15770 -21862 15782 -21826
rect 15724 -21874 15782 -21862
rect 15982 -21686 16040 -21674
rect 15982 -21722 15994 -21686
rect 16028 -21722 16040 -21686
rect 15982 -21756 16040 -21722
rect 15982 -21792 15994 -21756
rect 16028 -21792 16040 -21756
rect 15982 -21826 16040 -21792
rect 15982 -21862 15994 -21826
rect 16028 -21862 16040 -21826
rect 15982 -21874 16040 -21862
rect 16240 -21686 16298 -21674
rect 16240 -21722 16252 -21686
rect 16286 -21722 16298 -21686
rect 16240 -21756 16298 -21722
rect 16240 -21792 16252 -21756
rect 16286 -21792 16298 -21756
rect 16240 -21826 16298 -21792
rect 16240 -21862 16252 -21826
rect 16286 -21862 16298 -21826
rect 16240 -21874 16298 -21862
rect 16498 -21686 16556 -21674
rect 16498 -21722 16510 -21686
rect 16544 -21722 16556 -21686
rect 16498 -21756 16556 -21722
rect 16498 -21792 16510 -21756
rect 16544 -21792 16556 -21756
rect 16498 -21826 16556 -21792
rect 16498 -21862 16510 -21826
rect 16544 -21862 16556 -21826
rect 16498 -21874 16556 -21862
rect 9101 -22105 9159 -22093
rect 9101 -22141 9113 -22105
rect 9147 -22141 9159 -22105
rect 9101 -22175 9159 -22141
rect 9101 -22211 9113 -22175
rect 9147 -22211 9159 -22175
rect 9101 -22245 9159 -22211
rect 9101 -22281 9113 -22245
rect 9147 -22281 9159 -22245
rect 9101 -22293 9159 -22281
rect 9359 -22105 9417 -22093
rect 9359 -22141 9371 -22105
rect 9405 -22141 9417 -22105
rect 9359 -22175 9417 -22141
rect 9359 -22211 9371 -22175
rect 9405 -22211 9417 -22175
rect 9359 -22245 9417 -22211
rect 9359 -22281 9371 -22245
rect 9405 -22281 9417 -22245
rect 9359 -22293 9417 -22281
rect 9617 -22105 9675 -22093
rect 9617 -22141 9629 -22105
rect 9663 -22141 9675 -22105
rect 9617 -22175 9675 -22141
rect 9617 -22211 9629 -22175
rect 9663 -22211 9675 -22175
rect 9617 -22246 9675 -22211
rect 9617 -22282 9629 -22246
rect 9663 -22282 9675 -22246
rect 9617 -22293 9675 -22282
rect 9875 -22105 9933 -22093
rect 9875 -22141 9887 -22105
rect 9921 -22141 9933 -22105
rect 9875 -22175 9933 -22141
rect 9875 -22211 9887 -22175
rect 9921 -22211 9933 -22175
rect 9875 -22245 9933 -22211
rect 9875 -22281 9887 -22245
rect 9921 -22281 9933 -22245
rect 9875 -22293 9933 -22281
rect 10133 -22105 10191 -22093
rect 10133 -22141 10145 -22105
rect 10179 -22141 10191 -22105
rect 10133 -22175 10191 -22141
rect 10133 -22211 10145 -22175
rect 10179 -22211 10191 -22175
rect 10133 -22245 10191 -22211
rect 10133 -22281 10145 -22245
rect 10179 -22281 10191 -22245
rect 10133 -22293 10191 -22281
rect 10391 -22105 10449 -22093
rect 10391 -22141 10403 -22105
rect 10437 -22141 10449 -22105
rect 10391 -22175 10449 -22141
rect 10391 -22211 10403 -22175
rect 10437 -22211 10449 -22175
rect 10391 -22245 10449 -22211
rect 10391 -22281 10403 -22245
rect 10437 -22281 10449 -22245
rect 10391 -22293 10449 -22281
rect 10649 -22105 10707 -22093
rect 10649 -22141 10661 -22105
rect 10695 -22141 10707 -22105
rect 10649 -22175 10707 -22141
rect 10649 -22211 10661 -22175
rect 10695 -22211 10707 -22175
rect 10649 -22245 10707 -22211
rect 10649 -22281 10661 -22245
rect 10695 -22281 10707 -22245
rect 10649 -22293 10707 -22281
rect 10907 -22105 10965 -22093
rect 10907 -22141 10919 -22105
rect 10953 -22141 10965 -22105
rect 10907 -22175 10965 -22141
rect 10907 -22211 10919 -22175
rect 10953 -22211 10965 -22175
rect 10907 -22245 10965 -22211
rect 10907 -22281 10919 -22245
rect 10953 -22281 10965 -22245
rect 10907 -22293 10965 -22281
rect 11165 -22105 11223 -22093
rect 11165 -22141 11177 -22105
rect 11211 -22141 11223 -22105
rect 11165 -22175 11223 -22141
rect 11165 -22211 11177 -22175
rect 11211 -22211 11223 -22175
rect 11165 -22245 11223 -22211
rect 11165 -22281 11177 -22245
rect 11211 -22281 11223 -22245
rect 11165 -22293 11223 -22281
rect 11771 -22105 11829 -22093
rect 11771 -22141 11783 -22105
rect 11817 -22141 11829 -22105
rect 11771 -22175 11829 -22141
rect 11771 -22211 11783 -22175
rect 11817 -22211 11829 -22175
rect 11771 -22245 11829 -22211
rect 11771 -22281 11783 -22245
rect 11817 -22281 11829 -22245
rect 11771 -22293 11829 -22281
rect 12029 -22105 12087 -22093
rect 12029 -22141 12041 -22105
rect 12075 -22141 12087 -22105
rect 12029 -22175 12087 -22141
rect 12029 -22211 12041 -22175
rect 12075 -22211 12087 -22175
rect 12029 -22245 12087 -22211
rect 12029 -22281 12041 -22245
rect 12075 -22281 12087 -22245
rect 12029 -22293 12087 -22281
rect 12287 -22105 12345 -22093
rect 12287 -22141 12299 -22105
rect 12333 -22141 12345 -22105
rect 12287 -22175 12345 -22141
rect 12287 -22211 12299 -22175
rect 12333 -22211 12345 -22175
rect 12287 -22246 12345 -22211
rect 12287 -22282 12299 -22246
rect 12333 -22282 12345 -22246
rect 12287 -22293 12345 -22282
rect 12545 -22105 12603 -22093
rect 12545 -22141 12557 -22105
rect 12591 -22141 12603 -22105
rect 12545 -22175 12603 -22141
rect 12545 -22211 12557 -22175
rect 12591 -22211 12603 -22175
rect 12545 -22245 12603 -22211
rect 12545 -22281 12557 -22245
rect 12591 -22281 12603 -22245
rect 12545 -22293 12603 -22281
rect 12803 -22105 12861 -22093
rect 12803 -22141 12815 -22105
rect 12849 -22141 12861 -22105
rect 12803 -22175 12861 -22141
rect 12803 -22211 12815 -22175
rect 12849 -22211 12861 -22175
rect 12803 -22245 12861 -22211
rect 12803 -22281 12815 -22245
rect 12849 -22281 12861 -22245
rect 12803 -22293 12861 -22281
rect 13061 -22105 13119 -22093
rect 13061 -22141 13073 -22105
rect 13107 -22141 13119 -22105
rect 13061 -22175 13119 -22141
rect 13061 -22211 13073 -22175
rect 13107 -22211 13119 -22175
rect 13061 -22245 13119 -22211
rect 13061 -22281 13073 -22245
rect 13107 -22281 13119 -22245
rect 13061 -22293 13119 -22281
rect 13319 -22105 13377 -22093
rect 13319 -22141 13331 -22105
rect 13365 -22141 13377 -22105
rect 13319 -22175 13377 -22141
rect 13319 -22211 13331 -22175
rect 13365 -22211 13377 -22175
rect 13319 -22245 13377 -22211
rect 13319 -22281 13331 -22245
rect 13365 -22281 13377 -22245
rect 13319 -22293 13377 -22281
rect 13577 -22105 13635 -22093
rect 13577 -22141 13589 -22105
rect 13623 -22141 13635 -22105
rect 13577 -22175 13635 -22141
rect 13577 -22211 13589 -22175
rect 13623 -22211 13635 -22175
rect 13577 -22245 13635 -22211
rect 13577 -22281 13589 -22245
rect 13623 -22281 13635 -22245
rect 13577 -22293 13635 -22281
rect 13835 -22105 13893 -22093
rect 13835 -22141 13847 -22105
rect 13881 -22141 13893 -22105
rect 13835 -22175 13893 -22141
rect 13835 -22211 13847 -22175
rect 13881 -22211 13893 -22175
rect 13835 -22245 13893 -22211
rect 13835 -22281 13847 -22245
rect 13881 -22281 13893 -22245
rect 13835 -22293 13893 -22281
rect 14434 -22104 14492 -22092
rect 14434 -22140 14446 -22104
rect 14480 -22140 14492 -22104
rect 14434 -22174 14492 -22140
rect 14434 -22210 14446 -22174
rect 14480 -22210 14492 -22174
rect 14434 -22244 14492 -22210
rect 14434 -22280 14446 -22244
rect 14480 -22280 14492 -22244
rect 14434 -22292 14492 -22280
rect 14692 -22104 14750 -22092
rect 14692 -22140 14704 -22104
rect 14738 -22140 14750 -22104
rect 14692 -22174 14750 -22140
rect 14692 -22210 14704 -22174
rect 14738 -22210 14750 -22174
rect 14692 -22244 14750 -22210
rect 14692 -22280 14704 -22244
rect 14738 -22280 14750 -22244
rect 14692 -22292 14750 -22280
rect 14950 -22104 15008 -22092
rect 14950 -22140 14962 -22104
rect 14996 -22140 15008 -22104
rect 14950 -22174 15008 -22140
rect 14950 -22210 14962 -22174
rect 14996 -22210 15008 -22174
rect 14950 -22245 15008 -22210
rect 14950 -22281 14962 -22245
rect 14996 -22281 15008 -22245
rect 14950 -22292 15008 -22281
rect 15208 -22104 15266 -22092
rect 15208 -22140 15220 -22104
rect 15254 -22140 15266 -22104
rect 15208 -22174 15266 -22140
rect 15208 -22210 15220 -22174
rect 15254 -22210 15266 -22174
rect 15208 -22244 15266 -22210
rect 15208 -22280 15220 -22244
rect 15254 -22280 15266 -22244
rect 15208 -22292 15266 -22280
rect 15466 -22104 15524 -22092
rect 15466 -22140 15478 -22104
rect 15512 -22140 15524 -22104
rect 15466 -22174 15524 -22140
rect 15466 -22210 15478 -22174
rect 15512 -22210 15524 -22174
rect 15466 -22244 15524 -22210
rect 15466 -22280 15478 -22244
rect 15512 -22280 15524 -22244
rect 15466 -22292 15524 -22280
rect 15724 -22104 15782 -22092
rect 15724 -22140 15736 -22104
rect 15770 -22140 15782 -22104
rect 15724 -22174 15782 -22140
rect 15724 -22210 15736 -22174
rect 15770 -22210 15782 -22174
rect 15724 -22244 15782 -22210
rect 15724 -22280 15736 -22244
rect 15770 -22280 15782 -22244
rect 15724 -22292 15782 -22280
rect 15982 -22104 16040 -22092
rect 15982 -22140 15994 -22104
rect 16028 -22140 16040 -22104
rect 15982 -22174 16040 -22140
rect 15982 -22210 15994 -22174
rect 16028 -22210 16040 -22174
rect 15982 -22244 16040 -22210
rect 15982 -22280 15994 -22244
rect 16028 -22280 16040 -22244
rect 15982 -22292 16040 -22280
rect 16240 -22104 16298 -22092
rect 16240 -22140 16252 -22104
rect 16286 -22140 16298 -22104
rect 16240 -22174 16298 -22140
rect 16240 -22210 16252 -22174
rect 16286 -22210 16298 -22174
rect 16240 -22244 16298 -22210
rect 16240 -22280 16252 -22244
rect 16286 -22280 16298 -22244
rect 16240 -22292 16298 -22280
rect 16498 -22104 16556 -22092
rect 16498 -22140 16510 -22104
rect 16544 -22140 16556 -22104
rect 16498 -22174 16556 -22140
rect 16498 -22210 16510 -22174
rect 16544 -22210 16556 -22174
rect 16498 -22244 16556 -22210
rect 16498 -22280 16510 -22244
rect 16544 -22280 16556 -22244
rect 16498 -22292 16556 -22280
rect 9101 -22523 9159 -22511
rect 9101 -22559 9113 -22523
rect 9147 -22559 9159 -22523
rect 9101 -22593 9159 -22559
rect 9101 -22629 9113 -22593
rect 9147 -22629 9159 -22593
rect 9101 -22663 9159 -22629
rect 9101 -22699 9113 -22663
rect 9147 -22699 9159 -22663
rect 9101 -22711 9159 -22699
rect 9359 -22523 9417 -22511
rect 9359 -22559 9371 -22523
rect 9405 -22559 9417 -22523
rect 9359 -22593 9417 -22559
rect 9359 -22629 9371 -22593
rect 9405 -22629 9417 -22593
rect 9359 -22663 9417 -22629
rect 9359 -22699 9371 -22663
rect 9405 -22699 9417 -22663
rect 9359 -22711 9417 -22699
rect 9617 -22523 9675 -22511
rect 9617 -22559 9629 -22523
rect 9663 -22559 9675 -22523
rect 9617 -22593 9675 -22559
rect 9617 -22629 9629 -22593
rect 9663 -22629 9675 -22593
rect 9617 -22664 9675 -22629
rect 9617 -22700 9629 -22664
rect 9663 -22700 9675 -22664
rect 9617 -22711 9675 -22700
rect 9875 -22523 9933 -22511
rect 9875 -22559 9887 -22523
rect 9921 -22559 9933 -22523
rect 9875 -22593 9933 -22559
rect 9875 -22629 9887 -22593
rect 9921 -22629 9933 -22593
rect 9875 -22663 9933 -22629
rect 9875 -22699 9887 -22663
rect 9921 -22699 9933 -22663
rect 9875 -22711 9933 -22699
rect 10133 -22523 10191 -22511
rect 10133 -22559 10145 -22523
rect 10179 -22559 10191 -22523
rect 10133 -22593 10191 -22559
rect 10133 -22629 10145 -22593
rect 10179 -22629 10191 -22593
rect 10133 -22663 10191 -22629
rect 10133 -22699 10145 -22663
rect 10179 -22699 10191 -22663
rect 10133 -22711 10191 -22699
rect 10391 -22523 10449 -22511
rect 10391 -22559 10403 -22523
rect 10437 -22559 10449 -22523
rect 10391 -22593 10449 -22559
rect 10391 -22629 10403 -22593
rect 10437 -22629 10449 -22593
rect 10391 -22663 10449 -22629
rect 10391 -22699 10403 -22663
rect 10437 -22699 10449 -22663
rect 10391 -22711 10449 -22699
rect 10649 -22523 10707 -22511
rect 10649 -22559 10661 -22523
rect 10695 -22559 10707 -22523
rect 10649 -22593 10707 -22559
rect 10649 -22629 10661 -22593
rect 10695 -22629 10707 -22593
rect 10649 -22663 10707 -22629
rect 10649 -22699 10661 -22663
rect 10695 -22699 10707 -22663
rect 10649 -22711 10707 -22699
rect 10907 -22523 10965 -22511
rect 10907 -22559 10919 -22523
rect 10953 -22559 10965 -22523
rect 10907 -22593 10965 -22559
rect 10907 -22629 10919 -22593
rect 10953 -22629 10965 -22593
rect 10907 -22663 10965 -22629
rect 10907 -22699 10919 -22663
rect 10953 -22699 10965 -22663
rect 10907 -22711 10965 -22699
rect 11165 -22523 11223 -22511
rect 11165 -22559 11177 -22523
rect 11211 -22559 11223 -22523
rect 11165 -22593 11223 -22559
rect 11165 -22629 11177 -22593
rect 11211 -22629 11223 -22593
rect 11165 -22663 11223 -22629
rect 11165 -22699 11177 -22663
rect 11211 -22699 11223 -22663
rect 11165 -22711 11223 -22699
rect 11771 -22523 11829 -22511
rect 11771 -22559 11783 -22523
rect 11817 -22559 11829 -22523
rect 11771 -22593 11829 -22559
rect 11771 -22629 11783 -22593
rect 11817 -22629 11829 -22593
rect 11771 -22663 11829 -22629
rect 11771 -22699 11783 -22663
rect 11817 -22699 11829 -22663
rect 11771 -22711 11829 -22699
rect 12029 -22523 12087 -22511
rect 12029 -22559 12041 -22523
rect 12075 -22559 12087 -22523
rect 12029 -22593 12087 -22559
rect 12029 -22629 12041 -22593
rect 12075 -22629 12087 -22593
rect 12029 -22663 12087 -22629
rect 12029 -22699 12041 -22663
rect 12075 -22699 12087 -22663
rect 12029 -22711 12087 -22699
rect 12287 -22523 12345 -22511
rect 12287 -22559 12299 -22523
rect 12333 -22559 12345 -22523
rect 12287 -22593 12345 -22559
rect 12287 -22629 12299 -22593
rect 12333 -22629 12345 -22593
rect 12287 -22664 12345 -22629
rect 12287 -22700 12299 -22664
rect 12333 -22700 12345 -22664
rect 12287 -22711 12345 -22700
rect 12545 -22523 12603 -22511
rect 12545 -22559 12557 -22523
rect 12591 -22559 12603 -22523
rect 12545 -22593 12603 -22559
rect 12545 -22629 12557 -22593
rect 12591 -22629 12603 -22593
rect 12545 -22663 12603 -22629
rect 12545 -22699 12557 -22663
rect 12591 -22699 12603 -22663
rect 12545 -22711 12603 -22699
rect 12803 -22523 12861 -22511
rect 12803 -22559 12815 -22523
rect 12849 -22559 12861 -22523
rect 12803 -22593 12861 -22559
rect 12803 -22629 12815 -22593
rect 12849 -22629 12861 -22593
rect 12803 -22663 12861 -22629
rect 12803 -22699 12815 -22663
rect 12849 -22699 12861 -22663
rect 12803 -22711 12861 -22699
rect 13061 -22523 13119 -22511
rect 13061 -22559 13073 -22523
rect 13107 -22559 13119 -22523
rect 13061 -22593 13119 -22559
rect 13061 -22629 13073 -22593
rect 13107 -22629 13119 -22593
rect 13061 -22663 13119 -22629
rect 13061 -22699 13073 -22663
rect 13107 -22699 13119 -22663
rect 13061 -22711 13119 -22699
rect 13319 -22523 13377 -22511
rect 13319 -22559 13331 -22523
rect 13365 -22559 13377 -22523
rect 13319 -22593 13377 -22559
rect 13319 -22629 13331 -22593
rect 13365 -22629 13377 -22593
rect 13319 -22663 13377 -22629
rect 13319 -22699 13331 -22663
rect 13365 -22699 13377 -22663
rect 13319 -22711 13377 -22699
rect 13577 -22523 13635 -22511
rect 13577 -22559 13589 -22523
rect 13623 -22559 13635 -22523
rect 13577 -22593 13635 -22559
rect 13577 -22629 13589 -22593
rect 13623 -22629 13635 -22593
rect 13577 -22663 13635 -22629
rect 13577 -22699 13589 -22663
rect 13623 -22699 13635 -22663
rect 13577 -22711 13635 -22699
rect 13835 -22523 13893 -22511
rect 13835 -22559 13847 -22523
rect 13881 -22559 13893 -22523
rect 13835 -22593 13893 -22559
rect 13835 -22629 13847 -22593
rect 13881 -22629 13893 -22593
rect 13835 -22663 13893 -22629
rect 13835 -22699 13847 -22663
rect 13881 -22699 13893 -22663
rect 13835 -22711 13893 -22699
rect 14434 -22522 14492 -22510
rect 14434 -22558 14446 -22522
rect 14480 -22558 14492 -22522
rect 14434 -22592 14492 -22558
rect 14434 -22628 14446 -22592
rect 14480 -22628 14492 -22592
rect 14434 -22662 14492 -22628
rect 14434 -22698 14446 -22662
rect 14480 -22698 14492 -22662
rect 14434 -22710 14492 -22698
rect 14692 -22522 14750 -22510
rect 14692 -22558 14704 -22522
rect 14738 -22558 14750 -22522
rect 14692 -22592 14750 -22558
rect 14692 -22628 14704 -22592
rect 14738 -22628 14750 -22592
rect 14692 -22662 14750 -22628
rect 14692 -22698 14704 -22662
rect 14738 -22698 14750 -22662
rect 14692 -22710 14750 -22698
rect 14950 -22522 15008 -22510
rect 14950 -22558 14962 -22522
rect 14996 -22558 15008 -22522
rect 14950 -22592 15008 -22558
rect 14950 -22628 14962 -22592
rect 14996 -22628 15008 -22592
rect 14950 -22663 15008 -22628
rect 14950 -22699 14962 -22663
rect 14996 -22699 15008 -22663
rect 14950 -22710 15008 -22699
rect 15208 -22522 15266 -22510
rect 15208 -22558 15220 -22522
rect 15254 -22558 15266 -22522
rect 15208 -22592 15266 -22558
rect 15208 -22628 15220 -22592
rect 15254 -22628 15266 -22592
rect 15208 -22662 15266 -22628
rect 15208 -22698 15220 -22662
rect 15254 -22698 15266 -22662
rect 15208 -22710 15266 -22698
rect 15466 -22522 15524 -22510
rect 15466 -22558 15478 -22522
rect 15512 -22558 15524 -22522
rect 15466 -22592 15524 -22558
rect 15466 -22628 15478 -22592
rect 15512 -22628 15524 -22592
rect 15466 -22662 15524 -22628
rect 15466 -22698 15478 -22662
rect 15512 -22698 15524 -22662
rect 15466 -22710 15524 -22698
rect 15724 -22522 15782 -22510
rect 15724 -22558 15736 -22522
rect 15770 -22558 15782 -22522
rect 15724 -22592 15782 -22558
rect 15724 -22628 15736 -22592
rect 15770 -22628 15782 -22592
rect 15724 -22662 15782 -22628
rect 15724 -22698 15736 -22662
rect 15770 -22698 15782 -22662
rect 15724 -22710 15782 -22698
rect 15982 -22522 16040 -22510
rect 15982 -22558 15994 -22522
rect 16028 -22558 16040 -22522
rect 15982 -22592 16040 -22558
rect 15982 -22628 15994 -22592
rect 16028 -22628 16040 -22592
rect 15982 -22662 16040 -22628
rect 15982 -22698 15994 -22662
rect 16028 -22698 16040 -22662
rect 15982 -22710 16040 -22698
rect 16240 -22522 16298 -22510
rect 16240 -22558 16252 -22522
rect 16286 -22558 16298 -22522
rect 16240 -22592 16298 -22558
rect 16240 -22628 16252 -22592
rect 16286 -22628 16298 -22592
rect 16240 -22662 16298 -22628
rect 16240 -22698 16252 -22662
rect 16286 -22698 16298 -22662
rect 16240 -22710 16298 -22698
rect 16498 -22522 16556 -22510
rect 16498 -22558 16510 -22522
rect 16544 -22558 16556 -22522
rect 16498 -22592 16556 -22558
rect 16498 -22628 16510 -22592
rect 16544 -22628 16556 -22592
rect 16498 -22662 16556 -22628
rect 16498 -22698 16510 -22662
rect 16544 -22698 16556 -22662
rect 16498 -22710 16556 -22698
rect 9101 -22941 9159 -22929
rect 9101 -22977 9113 -22941
rect 9147 -22977 9159 -22941
rect 9101 -23011 9159 -22977
rect 9101 -23047 9113 -23011
rect 9147 -23047 9159 -23011
rect 9101 -23081 9159 -23047
rect 9101 -23117 9113 -23081
rect 9147 -23117 9159 -23081
rect 9101 -23129 9159 -23117
rect 9359 -22941 9417 -22929
rect 9359 -22977 9371 -22941
rect 9405 -22977 9417 -22941
rect 9359 -23011 9417 -22977
rect 9359 -23047 9371 -23011
rect 9405 -23047 9417 -23011
rect 9359 -23081 9417 -23047
rect 9359 -23117 9371 -23081
rect 9405 -23117 9417 -23081
rect 9359 -23129 9417 -23117
rect 9617 -22941 9675 -22929
rect 9617 -22977 9629 -22941
rect 9663 -22977 9675 -22941
rect 9617 -23011 9675 -22977
rect 9617 -23047 9629 -23011
rect 9663 -23047 9675 -23011
rect 9617 -23082 9675 -23047
rect 9617 -23118 9629 -23082
rect 9663 -23118 9675 -23082
rect 9617 -23129 9675 -23118
rect 9875 -22941 9933 -22929
rect 9875 -22977 9887 -22941
rect 9921 -22977 9933 -22941
rect 9875 -23011 9933 -22977
rect 9875 -23047 9887 -23011
rect 9921 -23047 9933 -23011
rect 9875 -23081 9933 -23047
rect 9875 -23117 9887 -23081
rect 9921 -23117 9933 -23081
rect 9875 -23129 9933 -23117
rect 10133 -22941 10191 -22929
rect 10133 -22977 10145 -22941
rect 10179 -22977 10191 -22941
rect 10133 -23011 10191 -22977
rect 10133 -23047 10145 -23011
rect 10179 -23047 10191 -23011
rect 10133 -23081 10191 -23047
rect 10133 -23117 10145 -23081
rect 10179 -23117 10191 -23081
rect 10133 -23129 10191 -23117
rect 10391 -22941 10449 -22929
rect 10391 -22977 10403 -22941
rect 10437 -22977 10449 -22941
rect 10391 -23011 10449 -22977
rect 10391 -23047 10403 -23011
rect 10437 -23047 10449 -23011
rect 10391 -23081 10449 -23047
rect 10391 -23117 10403 -23081
rect 10437 -23117 10449 -23081
rect 10391 -23129 10449 -23117
rect 10649 -22941 10707 -22929
rect 10649 -22977 10661 -22941
rect 10695 -22977 10707 -22941
rect 10649 -23011 10707 -22977
rect 10649 -23047 10661 -23011
rect 10695 -23047 10707 -23011
rect 10649 -23081 10707 -23047
rect 10649 -23117 10661 -23081
rect 10695 -23117 10707 -23081
rect 10649 -23129 10707 -23117
rect 10907 -22941 10965 -22929
rect 10907 -22977 10919 -22941
rect 10953 -22977 10965 -22941
rect 10907 -23011 10965 -22977
rect 10907 -23047 10919 -23011
rect 10953 -23047 10965 -23011
rect 10907 -23081 10965 -23047
rect 10907 -23117 10919 -23081
rect 10953 -23117 10965 -23081
rect 10907 -23129 10965 -23117
rect 11165 -22941 11223 -22929
rect 11165 -22977 11177 -22941
rect 11211 -22977 11223 -22941
rect 11165 -23011 11223 -22977
rect 11165 -23047 11177 -23011
rect 11211 -23047 11223 -23011
rect 11165 -23081 11223 -23047
rect 11165 -23117 11177 -23081
rect 11211 -23117 11223 -23081
rect 11165 -23129 11223 -23117
rect 11771 -22941 11829 -22929
rect 11771 -22977 11783 -22941
rect 11817 -22977 11829 -22941
rect 11771 -23011 11829 -22977
rect 11771 -23047 11783 -23011
rect 11817 -23047 11829 -23011
rect 11771 -23081 11829 -23047
rect 11771 -23117 11783 -23081
rect 11817 -23117 11829 -23081
rect 11771 -23129 11829 -23117
rect 12029 -22941 12087 -22929
rect 12029 -22977 12041 -22941
rect 12075 -22977 12087 -22941
rect 12029 -23011 12087 -22977
rect 12029 -23047 12041 -23011
rect 12075 -23047 12087 -23011
rect 12029 -23081 12087 -23047
rect 12029 -23117 12041 -23081
rect 12075 -23117 12087 -23081
rect 12029 -23129 12087 -23117
rect 12287 -22941 12345 -22929
rect 12287 -22977 12299 -22941
rect 12333 -22977 12345 -22941
rect 12287 -23011 12345 -22977
rect 12287 -23047 12299 -23011
rect 12333 -23047 12345 -23011
rect 12287 -23082 12345 -23047
rect 12287 -23118 12299 -23082
rect 12333 -23118 12345 -23082
rect 12287 -23129 12345 -23118
rect 12545 -22941 12603 -22929
rect 12545 -22977 12557 -22941
rect 12591 -22977 12603 -22941
rect 12545 -23011 12603 -22977
rect 12545 -23047 12557 -23011
rect 12591 -23047 12603 -23011
rect 12545 -23081 12603 -23047
rect 12545 -23117 12557 -23081
rect 12591 -23117 12603 -23081
rect 12545 -23129 12603 -23117
rect 12803 -22941 12861 -22929
rect 12803 -22977 12815 -22941
rect 12849 -22977 12861 -22941
rect 12803 -23011 12861 -22977
rect 12803 -23047 12815 -23011
rect 12849 -23047 12861 -23011
rect 12803 -23081 12861 -23047
rect 12803 -23117 12815 -23081
rect 12849 -23117 12861 -23081
rect 12803 -23129 12861 -23117
rect 13061 -22941 13119 -22929
rect 13061 -22977 13073 -22941
rect 13107 -22977 13119 -22941
rect 13061 -23011 13119 -22977
rect 13061 -23047 13073 -23011
rect 13107 -23047 13119 -23011
rect 13061 -23081 13119 -23047
rect 13061 -23117 13073 -23081
rect 13107 -23117 13119 -23081
rect 13061 -23129 13119 -23117
rect 13319 -22941 13377 -22929
rect 13319 -22977 13331 -22941
rect 13365 -22977 13377 -22941
rect 13319 -23011 13377 -22977
rect 13319 -23047 13331 -23011
rect 13365 -23047 13377 -23011
rect 13319 -23081 13377 -23047
rect 13319 -23117 13331 -23081
rect 13365 -23117 13377 -23081
rect 13319 -23129 13377 -23117
rect 13577 -22941 13635 -22929
rect 13577 -22977 13589 -22941
rect 13623 -22977 13635 -22941
rect 13577 -23011 13635 -22977
rect 13577 -23047 13589 -23011
rect 13623 -23047 13635 -23011
rect 13577 -23081 13635 -23047
rect 13577 -23117 13589 -23081
rect 13623 -23117 13635 -23081
rect 13577 -23129 13635 -23117
rect 13835 -22941 13893 -22929
rect 13835 -22977 13847 -22941
rect 13881 -22977 13893 -22941
rect 13835 -23011 13893 -22977
rect 13835 -23047 13847 -23011
rect 13881 -23047 13893 -23011
rect 13835 -23081 13893 -23047
rect 13835 -23117 13847 -23081
rect 13881 -23117 13893 -23081
rect 13835 -23129 13893 -23117
rect 14434 -22940 14492 -22928
rect 14434 -22976 14446 -22940
rect 14480 -22976 14492 -22940
rect 14434 -23010 14492 -22976
rect 14434 -23046 14446 -23010
rect 14480 -23046 14492 -23010
rect 14434 -23080 14492 -23046
rect 14434 -23116 14446 -23080
rect 14480 -23116 14492 -23080
rect 14434 -23128 14492 -23116
rect 14692 -22940 14750 -22928
rect 14692 -22976 14704 -22940
rect 14738 -22976 14750 -22940
rect 14692 -23010 14750 -22976
rect 14692 -23046 14704 -23010
rect 14738 -23046 14750 -23010
rect 14692 -23080 14750 -23046
rect 14692 -23116 14704 -23080
rect 14738 -23116 14750 -23080
rect 14692 -23128 14750 -23116
rect 14950 -22940 15008 -22928
rect 14950 -22976 14962 -22940
rect 14996 -22976 15008 -22940
rect 14950 -23010 15008 -22976
rect 14950 -23046 14962 -23010
rect 14996 -23046 15008 -23010
rect 14950 -23081 15008 -23046
rect 14950 -23117 14962 -23081
rect 14996 -23117 15008 -23081
rect 14950 -23128 15008 -23117
rect 15208 -22940 15266 -22928
rect 15208 -22976 15220 -22940
rect 15254 -22976 15266 -22940
rect 15208 -23010 15266 -22976
rect 15208 -23046 15220 -23010
rect 15254 -23046 15266 -23010
rect 15208 -23080 15266 -23046
rect 15208 -23116 15220 -23080
rect 15254 -23116 15266 -23080
rect 15208 -23128 15266 -23116
rect 15466 -22940 15524 -22928
rect 15466 -22976 15478 -22940
rect 15512 -22976 15524 -22940
rect 15466 -23010 15524 -22976
rect 15466 -23046 15478 -23010
rect 15512 -23046 15524 -23010
rect 15466 -23080 15524 -23046
rect 15466 -23116 15478 -23080
rect 15512 -23116 15524 -23080
rect 15466 -23128 15524 -23116
rect 15724 -22940 15782 -22928
rect 15724 -22976 15736 -22940
rect 15770 -22976 15782 -22940
rect 15724 -23010 15782 -22976
rect 15724 -23046 15736 -23010
rect 15770 -23046 15782 -23010
rect 15724 -23080 15782 -23046
rect 15724 -23116 15736 -23080
rect 15770 -23116 15782 -23080
rect 15724 -23128 15782 -23116
rect 15982 -22940 16040 -22928
rect 15982 -22976 15994 -22940
rect 16028 -22976 16040 -22940
rect 15982 -23010 16040 -22976
rect 15982 -23046 15994 -23010
rect 16028 -23046 16040 -23010
rect 15982 -23080 16040 -23046
rect 15982 -23116 15994 -23080
rect 16028 -23116 16040 -23080
rect 15982 -23128 16040 -23116
rect 16240 -22940 16298 -22928
rect 16240 -22976 16252 -22940
rect 16286 -22976 16298 -22940
rect 16240 -23010 16298 -22976
rect 16240 -23046 16252 -23010
rect 16286 -23046 16298 -23010
rect 16240 -23080 16298 -23046
rect 16240 -23116 16252 -23080
rect 16286 -23116 16298 -23080
rect 16240 -23128 16298 -23116
rect 16498 -22940 16556 -22928
rect 16498 -22976 16510 -22940
rect 16544 -22976 16556 -22940
rect 16498 -23010 16556 -22976
rect 16498 -23046 16510 -23010
rect 16544 -23046 16556 -23010
rect 16498 -23080 16556 -23046
rect 16498 -23116 16510 -23080
rect 16544 -23116 16556 -23080
rect 16498 -23128 16556 -23116
rect 9101 -23359 9159 -23347
rect 9101 -23395 9113 -23359
rect 9147 -23395 9159 -23359
rect 9101 -23429 9159 -23395
rect 9101 -23465 9113 -23429
rect 9147 -23465 9159 -23429
rect 9101 -23499 9159 -23465
rect 9101 -23535 9113 -23499
rect 9147 -23535 9159 -23499
rect 9101 -23547 9159 -23535
rect 9359 -23359 9417 -23347
rect 9359 -23395 9371 -23359
rect 9405 -23395 9417 -23359
rect 9359 -23429 9417 -23395
rect 9359 -23465 9371 -23429
rect 9405 -23465 9417 -23429
rect 9359 -23499 9417 -23465
rect 9359 -23535 9371 -23499
rect 9405 -23535 9417 -23499
rect 9359 -23547 9417 -23535
rect 9617 -23359 9675 -23347
rect 9617 -23395 9629 -23359
rect 9663 -23395 9675 -23359
rect 9617 -23429 9675 -23395
rect 9617 -23465 9629 -23429
rect 9663 -23465 9675 -23429
rect 9617 -23500 9675 -23465
rect 9617 -23536 9629 -23500
rect 9663 -23536 9675 -23500
rect 9617 -23547 9675 -23536
rect 9875 -23359 9933 -23347
rect 9875 -23395 9887 -23359
rect 9921 -23395 9933 -23359
rect 9875 -23429 9933 -23395
rect 9875 -23465 9887 -23429
rect 9921 -23465 9933 -23429
rect 9875 -23499 9933 -23465
rect 9875 -23535 9887 -23499
rect 9921 -23535 9933 -23499
rect 9875 -23547 9933 -23535
rect 10133 -23359 10191 -23347
rect 10133 -23395 10145 -23359
rect 10179 -23395 10191 -23359
rect 10133 -23429 10191 -23395
rect 10133 -23465 10145 -23429
rect 10179 -23465 10191 -23429
rect 10133 -23499 10191 -23465
rect 10133 -23535 10145 -23499
rect 10179 -23535 10191 -23499
rect 10133 -23547 10191 -23535
rect 10391 -23359 10449 -23347
rect 10391 -23395 10403 -23359
rect 10437 -23395 10449 -23359
rect 10391 -23429 10449 -23395
rect 10391 -23465 10403 -23429
rect 10437 -23465 10449 -23429
rect 10391 -23499 10449 -23465
rect 10391 -23535 10403 -23499
rect 10437 -23535 10449 -23499
rect 10391 -23547 10449 -23535
rect 10649 -23359 10707 -23347
rect 10649 -23395 10661 -23359
rect 10695 -23395 10707 -23359
rect 10649 -23429 10707 -23395
rect 10649 -23465 10661 -23429
rect 10695 -23465 10707 -23429
rect 10649 -23499 10707 -23465
rect 10649 -23535 10661 -23499
rect 10695 -23535 10707 -23499
rect 10649 -23547 10707 -23535
rect 10907 -23359 10965 -23347
rect 10907 -23395 10919 -23359
rect 10953 -23395 10965 -23359
rect 10907 -23429 10965 -23395
rect 10907 -23465 10919 -23429
rect 10953 -23465 10965 -23429
rect 10907 -23499 10965 -23465
rect 10907 -23535 10919 -23499
rect 10953 -23535 10965 -23499
rect 10907 -23547 10965 -23535
rect 11165 -23359 11223 -23347
rect 11165 -23395 11177 -23359
rect 11211 -23395 11223 -23359
rect 11165 -23429 11223 -23395
rect 11165 -23465 11177 -23429
rect 11211 -23465 11223 -23429
rect 11165 -23499 11223 -23465
rect 11165 -23535 11177 -23499
rect 11211 -23535 11223 -23499
rect 11165 -23547 11223 -23535
rect 11771 -23359 11829 -23347
rect 11771 -23395 11783 -23359
rect 11817 -23395 11829 -23359
rect 11771 -23429 11829 -23395
rect 11771 -23465 11783 -23429
rect 11817 -23465 11829 -23429
rect 11771 -23499 11829 -23465
rect 11771 -23535 11783 -23499
rect 11817 -23535 11829 -23499
rect 11771 -23547 11829 -23535
rect 12029 -23359 12087 -23347
rect 12029 -23395 12041 -23359
rect 12075 -23395 12087 -23359
rect 12029 -23429 12087 -23395
rect 12029 -23465 12041 -23429
rect 12075 -23465 12087 -23429
rect 12029 -23499 12087 -23465
rect 12029 -23535 12041 -23499
rect 12075 -23535 12087 -23499
rect 12029 -23547 12087 -23535
rect 12287 -23359 12345 -23347
rect 12287 -23395 12299 -23359
rect 12333 -23395 12345 -23359
rect 12287 -23429 12345 -23395
rect 12287 -23465 12299 -23429
rect 12333 -23465 12345 -23429
rect 12287 -23500 12345 -23465
rect 12287 -23536 12299 -23500
rect 12333 -23536 12345 -23500
rect 12287 -23547 12345 -23536
rect 12545 -23359 12603 -23347
rect 12545 -23395 12557 -23359
rect 12591 -23395 12603 -23359
rect 12545 -23429 12603 -23395
rect 12545 -23465 12557 -23429
rect 12591 -23465 12603 -23429
rect 12545 -23499 12603 -23465
rect 12545 -23535 12557 -23499
rect 12591 -23535 12603 -23499
rect 12545 -23547 12603 -23535
rect 12803 -23359 12861 -23347
rect 12803 -23395 12815 -23359
rect 12849 -23395 12861 -23359
rect 12803 -23429 12861 -23395
rect 12803 -23465 12815 -23429
rect 12849 -23465 12861 -23429
rect 12803 -23499 12861 -23465
rect 12803 -23535 12815 -23499
rect 12849 -23535 12861 -23499
rect 12803 -23547 12861 -23535
rect 13061 -23359 13119 -23347
rect 13061 -23395 13073 -23359
rect 13107 -23395 13119 -23359
rect 13061 -23429 13119 -23395
rect 13061 -23465 13073 -23429
rect 13107 -23465 13119 -23429
rect 13061 -23499 13119 -23465
rect 13061 -23535 13073 -23499
rect 13107 -23535 13119 -23499
rect 13061 -23547 13119 -23535
rect 13319 -23359 13377 -23347
rect 13319 -23395 13331 -23359
rect 13365 -23395 13377 -23359
rect 13319 -23429 13377 -23395
rect 13319 -23465 13331 -23429
rect 13365 -23465 13377 -23429
rect 13319 -23499 13377 -23465
rect 13319 -23535 13331 -23499
rect 13365 -23535 13377 -23499
rect 13319 -23547 13377 -23535
rect 13577 -23359 13635 -23347
rect 13577 -23395 13589 -23359
rect 13623 -23395 13635 -23359
rect 13577 -23429 13635 -23395
rect 13577 -23465 13589 -23429
rect 13623 -23465 13635 -23429
rect 13577 -23499 13635 -23465
rect 13577 -23535 13589 -23499
rect 13623 -23535 13635 -23499
rect 13577 -23547 13635 -23535
rect 13835 -23359 13893 -23347
rect 13835 -23395 13847 -23359
rect 13881 -23395 13893 -23359
rect 13835 -23429 13893 -23395
rect 13835 -23465 13847 -23429
rect 13881 -23465 13893 -23429
rect 13835 -23499 13893 -23465
rect 13835 -23535 13847 -23499
rect 13881 -23535 13893 -23499
rect 13835 -23547 13893 -23535
rect 14434 -23358 14492 -23346
rect 14434 -23394 14446 -23358
rect 14480 -23394 14492 -23358
rect 14434 -23428 14492 -23394
rect 14434 -23464 14446 -23428
rect 14480 -23464 14492 -23428
rect 14434 -23498 14492 -23464
rect 14434 -23534 14446 -23498
rect 14480 -23534 14492 -23498
rect 14434 -23546 14492 -23534
rect 14692 -23358 14750 -23346
rect 14692 -23394 14704 -23358
rect 14738 -23394 14750 -23358
rect 14692 -23428 14750 -23394
rect 14692 -23464 14704 -23428
rect 14738 -23464 14750 -23428
rect 14692 -23498 14750 -23464
rect 14692 -23534 14704 -23498
rect 14738 -23534 14750 -23498
rect 14692 -23546 14750 -23534
rect 14950 -23358 15008 -23346
rect 14950 -23394 14962 -23358
rect 14996 -23394 15008 -23358
rect 14950 -23428 15008 -23394
rect 14950 -23464 14962 -23428
rect 14996 -23464 15008 -23428
rect 14950 -23499 15008 -23464
rect 14950 -23535 14962 -23499
rect 14996 -23535 15008 -23499
rect 14950 -23546 15008 -23535
rect 15208 -23358 15266 -23346
rect 15208 -23394 15220 -23358
rect 15254 -23394 15266 -23358
rect 15208 -23428 15266 -23394
rect 15208 -23464 15220 -23428
rect 15254 -23464 15266 -23428
rect 15208 -23498 15266 -23464
rect 15208 -23534 15220 -23498
rect 15254 -23534 15266 -23498
rect 15208 -23546 15266 -23534
rect 15466 -23358 15524 -23346
rect 15466 -23394 15478 -23358
rect 15512 -23394 15524 -23358
rect 15466 -23428 15524 -23394
rect 15466 -23464 15478 -23428
rect 15512 -23464 15524 -23428
rect 15466 -23498 15524 -23464
rect 15466 -23534 15478 -23498
rect 15512 -23534 15524 -23498
rect 15466 -23546 15524 -23534
rect 15724 -23358 15782 -23346
rect 15724 -23394 15736 -23358
rect 15770 -23394 15782 -23358
rect 15724 -23428 15782 -23394
rect 15724 -23464 15736 -23428
rect 15770 -23464 15782 -23428
rect 15724 -23498 15782 -23464
rect 15724 -23534 15736 -23498
rect 15770 -23534 15782 -23498
rect 15724 -23546 15782 -23534
rect 15982 -23358 16040 -23346
rect 15982 -23394 15994 -23358
rect 16028 -23394 16040 -23358
rect 15982 -23428 16040 -23394
rect 15982 -23464 15994 -23428
rect 16028 -23464 16040 -23428
rect 15982 -23498 16040 -23464
rect 15982 -23534 15994 -23498
rect 16028 -23534 16040 -23498
rect 15982 -23546 16040 -23534
rect 16240 -23358 16298 -23346
rect 16240 -23394 16252 -23358
rect 16286 -23394 16298 -23358
rect 16240 -23428 16298 -23394
rect 16240 -23464 16252 -23428
rect 16286 -23464 16298 -23428
rect 16240 -23498 16298 -23464
rect 16240 -23534 16252 -23498
rect 16286 -23534 16298 -23498
rect 16240 -23546 16298 -23534
rect 16498 -23358 16556 -23346
rect 16498 -23394 16510 -23358
rect 16544 -23394 16556 -23358
rect 16498 -23428 16556 -23394
rect 16498 -23464 16510 -23428
rect 16544 -23464 16556 -23428
rect 16498 -23498 16556 -23464
rect 16498 -23534 16510 -23498
rect 16544 -23534 16556 -23498
rect 16498 -23546 16556 -23534
rect 9101 -23777 9159 -23765
rect 9101 -23813 9113 -23777
rect 9147 -23813 9159 -23777
rect 9101 -23847 9159 -23813
rect 9101 -23883 9113 -23847
rect 9147 -23883 9159 -23847
rect 9101 -23917 9159 -23883
rect 9101 -23953 9113 -23917
rect 9147 -23953 9159 -23917
rect 9101 -23965 9159 -23953
rect 9359 -23777 9417 -23765
rect 9359 -23813 9371 -23777
rect 9405 -23813 9417 -23777
rect 9359 -23847 9417 -23813
rect 9359 -23883 9371 -23847
rect 9405 -23883 9417 -23847
rect 9359 -23917 9417 -23883
rect 9359 -23953 9371 -23917
rect 9405 -23953 9417 -23917
rect 9359 -23965 9417 -23953
rect 9617 -23777 9675 -23765
rect 9617 -23813 9629 -23777
rect 9663 -23813 9675 -23777
rect 9617 -23847 9675 -23813
rect 9617 -23883 9629 -23847
rect 9663 -23883 9675 -23847
rect 9617 -23918 9675 -23883
rect 9617 -23954 9629 -23918
rect 9663 -23954 9675 -23918
rect 9617 -23965 9675 -23954
rect 9875 -23777 9933 -23765
rect 9875 -23813 9887 -23777
rect 9921 -23813 9933 -23777
rect 9875 -23847 9933 -23813
rect 9875 -23883 9887 -23847
rect 9921 -23883 9933 -23847
rect 9875 -23917 9933 -23883
rect 9875 -23953 9887 -23917
rect 9921 -23953 9933 -23917
rect 9875 -23965 9933 -23953
rect 10133 -23777 10191 -23765
rect 10133 -23813 10145 -23777
rect 10179 -23813 10191 -23777
rect 10133 -23847 10191 -23813
rect 10133 -23883 10145 -23847
rect 10179 -23883 10191 -23847
rect 10133 -23917 10191 -23883
rect 10133 -23953 10145 -23917
rect 10179 -23953 10191 -23917
rect 10133 -23965 10191 -23953
rect 10391 -23777 10449 -23765
rect 10391 -23813 10403 -23777
rect 10437 -23813 10449 -23777
rect 10391 -23847 10449 -23813
rect 10391 -23883 10403 -23847
rect 10437 -23883 10449 -23847
rect 10391 -23917 10449 -23883
rect 10391 -23953 10403 -23917
rect 10437 -23953 10449 -23917
rect 10391 -23965 10449 -23953
rect 10649 -23777 10707 -23765
rect 10649 -23813 10661 -23777
rect 10695 -23813 10707 -23777
rect 10649 -23847 10707 -23813
rect 10649 -23883 10661 -23847
rect 10695 -23883 10707 -23847
rect 10649 -23917 10707 -23883
rect 10649 -23953 10661 -23917
rect 10695 -23953 10707 -23917
rect 10649 -23965 10707 -23953
rect 10907 -23777 10965 -23765
rect 10907 -23813 10919 -23777
rect 10953 -23813 10965 -23777
rect 10907 -23847 10965 -23813
rect 10907 -23883 10919 -23847
rect 10953 -23883 10965 -23847
rect 10907 -23917 10965 -23883
rect 10907 -23953 10919 -23917
rect 10953 -23953 10965 -23917
rect 10907 -23965 10965 -23953
rect 11165 -23777 11223 -23765
rect 11165 -23813 11177 -23777
rect 11211 -23813 11223 -23777
rect 11165 -23847 11223 -23813
rect 11165 -23883 11177 -23847
rect 11211 -23883 11223 -23847
rect 11165 -23917 11223 -23883
rect 11165 -23953 11177 -23917
rect 11211 -23953 11223 -23917
rect 11165 -23965 11223 -23953
rect 11771 -23777 11829 -23765
rect 11771 -23813 11783 -23777
rect 11817 -23813 11829 -23777
rect 11771 -23847 11829 -23813
rect 11771 -23883 11783 -23847
rect 11817 -23883 11829 -23847
rect 11771 -23917 11829 -23883
rect 11771 -23953 11783 -23917
rect 11817 -23953 11829 -23917
rect 11771 -23965 11829 -23953
rect 12029 -23777 12087 -23765
rect 12029 -23813 12041 -23777
rect 12075 -23813 12087 -23777
rect 12029 -23847 12087 -23813
rect 12029 -23883 12041 -23847
rect 12075 -23883 12087 -23847
rect 12029 -23917 12087 -23883
rect 12029 -23953 12041 -23917
rect 12075 -23953 12087 -23917
rect 12029 -23965 12087 -23953
rect 12287 -23777 12345 -23765
rect 12287 -23813 12299 -23777
rect 12333 -23813 12345 -23777
rect 12287 -23847 12345 -23813
rect 12287 -23883 12299 -23847
rect 12333 -23883 12345 -23847
rect 12287 -23918 12345 -23883
rect 12287 -23954 12299 -23918
rect 12333 -23954 12345 -23918
rect 12287 -23965 12345 -23954
rect 12545 -23777 12603 -23765
rect 12545 -23813 12557 -23777
rect 12591 -23813 12603 -23777
rect 12545 -23847 12603 -23813
rect 12545 -23883 12557 -23847
rect 12591 -23883 12603 -23847
rect 12545 -23917 12603 -23883
rect 12545 -23953 12557 -23917
rect 12591 -23953 12603 -23917
rect 12545 -23965 12603 -23953
rect 12803 -23777 12861 -23765
rect 12803 -23813 12815 -23777
rect 12849 -23813 12861 -23777
rect 12803 -23847 12861 -23813
rect 12803 -23883 12815 -23847
rect 12849 -23883 12861 -23847
rect 12803 -23917 12861 -23883
rect 12803 -23953 12815 -23917
rect 12849 -23953 12861 -23917
rect 12803 -23965 12861 -23953
rect 13061 -23777 13119 -23765
rect 13061 -23813 13073 -23777
rect 13107 -23813 13119 -23777
rect 13061 -23847 13119 -23813
rect 13061 -23883 13073 -23847
rect 13107 -23883 13119 -23847
rect 13061 -23917 13119 -23883
rect 13061 -23953 13073 -23917
rect 13107 -23953 13119 -23917
rect 13061 -23965 13119 -23953
rect 13319 -23777 13377 -23765
rect 13319 -23813 13331 -23777
rect 13365 -23813 13377 -23777
rect 13319 -23847 13377 -23813
rect 13319 -23883 13331 -23847
rect 13365 -23883 13377 -23847
rect 13319 -23917 13377 -23883
rect 13319 -23953 13331 -23917
rect 13365 -23953 13377 -23917
rect 13319 -23965 13377 -23953
rect 13577 -23777 13635 -23765
rect 13577 -23813 13589 -23777
rect 13623 -23813 13635 -23777
rect 13577 -23847 13635 -23813
rect 13577 -23883 13589 -23847
rect 13623 -23883 13635 -23847
rect 13577 -23917 13635 -23883
rect 13577 -23953 13589 -23917
rect 13623 -23953 13635 -23917
rect 13577 -23965 13635 -23953
rect 13835 -23777 13893 -23765
rect 13835 -23813 13847 -23777
rect 13881 -23813 13893 -23777
rect 13835 -23847 13893 -23813
rect 13835 -23883 13847 -23847
rect 13881 -23883 13893 -23847
rect 13835 -23917 13893 -23883
rect 13835 -23953 13847 -23917
rect 13881 -23953 13893 -23917
rect 13835 -23965 13893 -23953
rect 14434 -23776 14492 -23764
rect 14434 -23812 14446 -23776
rect 14480 -23812 14492 -23776
rect 14434 -23846 14492 -23812
rect 14434 -23882 14446 -23846
rect 14480 -23882 14492 -23846
rect 14434 -23916 14492 -23882
rect 14434 -23952 14446 -23916
rect 14480 -23952 14492 -23916
rect 14434 -23964 14492 -23952
rect 14692 -23776 14750 -23764
rect 14692 -23812 14704 -23776
rect 14738 -23812 14750 -23776
rect 14692 -23846 14750 -23812
rect 14692 -23882 14704 -23846
rect 14738 -23882 14750 -23846
rect 14692 -23916 14750 -23882
rect 14692 -23952 14704 -23916
rect 14738 -23952 14750 -23916
rect 14692 -23964 14750 -23952
rect 14950 -23776 15008 -23764
rect 14950 -23812 14962 -23776
rect 14996 -23812 15008 -23776
rect 14950 -23846 15008 -23812
rect 14950 -23882 14962 -23846
rect 14996 -23882 15008 -23846
rect 14950 -23917 15008 -23882
rect 14950 -23953 14962 -23917
rect 14996 -23953 15008 -23917
rect 14950 -23964 15008 -23953
rect 15208 -23776 15266 -23764
rect 15208 -23812 15220 -23776
rect 15254 -23812 15266 -23776
rect 15208 -23846 15266 -23812
rect 15208 -23882 15220 -23846
rect 15254 -23882 15266 -23846
rect 15208 -23916 15266 -23882
rect 15208 -23952 15220 -23916
rect 15254 -23952 15266 -23916
rect 15208 -23964 15266 -23952
rect 15466 -23776 15524 -23764
rect 15466 -23812 15478 -23776
rect 15512 -23812 15524 -23776
rect 15466 -23846 15524 -23812
rect 15466 -23882 15478 -23846
rect 15512 -23882 15524 -23846
rect 15466 -23916 15524 -23882
rect 15466 -23952 15478 -23916
rect 15512 -23952 15524 -23916
rect 15466 -23964 15524 -23952
rect 15724 -23776 15782 -23764
rect 15724 -23812 15736 -23776
rect 15770 -23812 15782 -23776
rect 15724 -23846 15782 -23812
rect 15724 -23882 15736 -23846
rect 15770 -23882 15782 -23846
rect 15724 -23916 15782 -23882
rect 15724 -23952 15736 -23916
rect 15770 -23952 15782 -23916
rect 15724 -23964 15782 -23952
rect 15982 -23776 16040 -23764
rect 15982 -23812 15994 -23776
rect 16028 -23812 16040 -23776
rect 15982 -23846 16040 -23812
rect 15982 -23882 15994 -23846
rect 16028 -23882 16040 -23846
rect 15982 -23916 16040 -23882
rect 15982 -23952 15994 -23916
rect 16028 -23952 16040 -23916
rect 15982 -23964 16040 -23952
rect 16240 -23776 16298 -23764
rect 16240 -23812 16252 -23776
rect 16286 -23812 16298 -23776
rect 16240 -23846 16298 -23812
rect 16240 -23882 16252 -23846
rect 16286 -23882 16298 -23846
rect 16240 -23916 16298 -23882
rect 16240 -23952 16252 -23916
rect 16286 -23952 16298 -23916
rect 16240 -23964 16298 -23952
rect 16498 -23776 16556 -23764
rect 16498 -23812 16510 -23776
rect 16544 -23812 16556 -23776
rect 16498 -23846 16556 -23812
rect 16498 -23882 16510 -23846
rect 16544 -23882 16556 -23846
rect 16498 -23916 16556 -23882
rect 16498 -23952 16510 -23916
rect 16544 -23952 16556 -23916
rect 16498 -23964 16556 -23952
rect 8981 -24431 9039 -24417
rect 8981 -24465 8993 -24431
rect 9027 -24465 9039 -24431
rect 8981 -24499 9039 -24465
rect 8981 -24535 8993 -24499
rect 9027 -24535 9039 -24499
rect 8981 -24569 9039 -24535
rect 8981 -24603 8993 -24569
rect 9027 -24603 9039 -24569
rect 8981 -24617 9039 -24603
rect 9239 -24431 9297 -24417
rect 9239 -24465 9251 -24431
rect 9285 -24465 9297 -24431
rect 9239 -24499 9297 -24465
rect 9239 -24535 9251 -24499
rect 9285 -24535 9297 -24499
rect 9239 -24569 9297 -24535
rect 9239 -24603 9251 -24569
rect 9285 -24603 9297 -24569
rect 9239 -24617 9297 -24603
rect 9521 -24431 9579 -24417
rect 9521 -24465 9533 -24431
rect 9567 -24465 9579 -24431
rect 9521 -24499 9579 -24465
rect 9521 -24535 9533 -24499
rect 9567 -24535 9579 -24499
rect 9521 -24569 9579 -24535
rect 9521 -24603 9533 -24569
rect 9567 -24603 9579 -24569
rect 9521 -24617 9579 -24603
rect 9779 -24431 9837 -24417
rect 9779 -24465 9791 -24431
rect 9825 -24465 9837 -24431
rect 9779 -24499 9837 -24465
rect 9779 -24535 9791 -24499
rect 9825 -24535 9837 -24499
rect 9779 -24569 9837 -24535
rect 9779 -24603 9791 -24569
rect 9825 -24603 9837 -24569
rect 9779 -24617 9837 -24603
rect 10001 -24431 10059 -24417
rect 10001 -24465 10013 -24431
rect 10047 -24465 10059 -24431
rect 10001 -24499 10059 -24465
rect 10001 -24535 10013 -24499
rect 10047 -24535 10059 -24499
rect 10001 -24569 10059 -24535
rect 10001 -24603 10013 -24569
rect 10047 -24603 10059 -24569
rect 10001 -24617 10059 -24603
rect 10259 -24431 10317 -24417
rect 10259 -24465 10271 -24431
rect 10305 -24465 10317 -24431
rect 10259 -24499 10317 -24465
rect 10259 -24535 10271 -24499
rect 10305 -24535 10317 -24499
rect 10259 -24569 10317 -24535
rect 10259 -24603 10271 -24569
rect 10305 -24603 10317 -24569
rect 10259 -24617 10317 -24603
rect 10504 -24429 10562 -24415
rect 10504 -24463 10516 -24429
rect 10550 -24463 10562 -24429
rect 10504 -24497 10562 -24463
rect 10504 -24533 10516 -24497
rect 10550 -24533 10562 -24497
rect 10504 -24567 10562 -24533
rect 10504 -24601 10516 -24567
rect 10550 -24601 10562 -24567
rect 10504 -24615 10562 -24601
rect 10762 -24429 10820 -24415
rect 10762 -24463 10774 -24429
rect 10808 -24463 10820 -24429
rect 10762 -24497 10820 -24463
rect 10762 -24533 10774 -24497
rect 10808 -24533 10820 -24497
rect 10762 -24567 10820 -24533
rect 10762 -24601 10774 -24567
rect 10808 -24601 10820 -24567
rect 10762 -24615 10820 -24601
rect 11014 -24419 11072 -24405
rect 11014 -24453 11026 -24419
rect 11060 -24453 11072 -24419
rect 11014 -24487 11072 -24453
rect 11014 -24523 11026 -24487
rect 11060 -24523 11072 -24487
rect 11014 -24557 11072 -24523
rect 11014 -24591 11026 -24557
rect 11060 -24591 11072 -24557
rect 11014 -24605 11072 -24591
rect 11272 -24419 11330 -24405
rect 11272 -24453 11284 -24419
rect 11318 -24453 11330 -24419
rect 11272 -24487 11330 -24453
rect 11272 -24523 11284 -24487
rect 11318 -24523 11330 -24487
rect 11272 -24557 11330 -24523
rect 11272 -24591 11284 -24557
rect 11318 -24591 11330 -24557
rect 11272 -24605 11330 -24591
rect 11651 -24431 11709 -24417
rect 11651 -24465 11663 -24431
rect 11697 -24465 11709 -24431
rect 11651 -24499 11709 -24465
rect 11651 -24535 11663 -24499
rect 11697 -24535 11709 -24499
rect 11651 -24569 11709 -24535
rect 11651 -24603 11663 -24569
rect 11697 -24603 11709 -24569
rect 11651 -24617 11709 -24603
rect 11909 -24431 11967 -24417
rect 11909 -24465 11921 -24431
rect 11955 -24465 11967 -24431
rect 11909 -24499 11967 -24465
rect 11909 -24535 11921 -24499
rect 11955 -24535 11967 -24499
rect 11909 -24569 11967 -24535
rect 11909 -24603 11921 -24569
rect 11955 -24603 11967 -24569
rect 11909 -24617 11967 -24603
rect 12191 -24431 12249 -24417
rect 12191 -24465 12203 -24431
rect 12237 -24465 12249 -24431
rect 12191 -24499 12249 -24465
rect 12191 -24535 12203 -24499
rect 12237 -24535 12249 -24499
rect 12191 -24569 12249 -24535
rect 12191 -24603 12203 -24569
rect 12237 -24603 12249 -24569
rect 12191 -24617 12249 -24603
rect 12449 -24431 12507 -24417
rect 12449 -24465 12461 -24431
rect 12495 -24465 12507 -24431
rect 12449 -24499 12507 -24465
rect 12449 -24535 12461 -24499
rect 12495 -24535 12507 -24499
rect 12449 -24569 12507 -24535
rect 12449 -24603 12461 -24569
rect 12495 -24603 12507 -24569
rect 12449 -24617 12507 -24603
rect 12671 -24431 12729 -24417
rect 12671 -24465 12683 -24431
rect 12717 -24465 12729 -24431
rect 12671 -24499 12729 -24465
rect 12671 -24535 12683 -24499
rect 12717 -24535 12729 -24499
rect 12671 -24569 12729 -24535
rect 12671 -24603 12683 -24569
rect 12717 -24603 12729 -24569
rect 12671 -24617 12729 -24603
rect 12929 -24431 12987 -24417
rect 12929 -24465 12941 -24431
rect 12975 -24465 12987 -24431
rect 12929 -24499 12987 -24465
rect 12929 -24535 12941 -24499
rect 12975 -24535 12987 -24499
rect 12929 -24569 12987 -24535
rect 12929 -24603 12941 -24569
rect 12975 -24603 12987 -24569
rect 12929 -24617 12987 -24603
rect 13174 -24429 13232 -24415
rect 13174 -24463 13186 -24429
rect 13220 -24463 13232 -24429
rect 13174 -24497 13232 -24463
rect 13174 -24533 13186 -24497
rect 13220 -24533 13232 -24497
rect 13174 -24567 13232 -24533
rect 13174 -24601 13186 -24567
rect 13220 -24601 13232 -24567
rect 13174 -24615 13232 -24601
rect 13432 -24429 13490 -24415
rect 13432 -24463 13444 -24429
rect 13478 -24463 13490 -24429
rect 13432 -24497 13490 -24463
rect 13432 -24533 13444 -24497
rect 13478 -24533 13490 -24497
rect 13432 -24567 13490 -24533
rect 13432 -24601 13444 -24567
rect 13478 -24601 13490 -24567
rect 13432 -24615 13490 -24601
rect 13684 -24419 13742 -24405
rect 13684 -24453 13696 -24419
rect 13730 -24453 13742 -24419
rect 13684 -24487 13742 -24453
rect 13684 -24523 13696 -24487
rect 13730 -24523 13742 -24487
rect 13684 -24557 13742 -24523
rect 13684 -24591 13696 -24557
rect 13730 -24591 13742 -24557
rect 13684 -24605 13742 -24591
rect 13942 -24419 14000 -24405
rect 13942 -24453 13954 -24419
rect 13988 -24453 14000 -24419
rect 13942 -24487 14000 -24453
rect 13942 -24523 13954 -24487
rect 13988 -24523 14000 -24487
rect 13942 -24557 14000 -24523
rect 13942 -24591 13954 -24557
rect 13988 -24591 14000 -24557
rect 13942 -24605 14000 -24591
rect 14314 -24430 14372 -24416
rect 14314 -24464 14326 -24430
rect 14360 -24464 14372 -24430
rect 14314 -24498 14372 -24464
rect 14314 -24534 14326 -24498
rect 14360 -24534 14372 -24498
rect 14314 -24568 14372 -24534
rect 14314 -24602 14326 -24568
rect 14360 -24602 14372 -24568
rect 14314 -24616 14372 -24602
rect 14572 -24430 14630 -24416
rect 14572 -24464 14584 -24430
rect 14618 -24464 14630 -24430
rect 14572 -24498 14630 -24464
rect 14572 -24534 14584 -24498
rect 14618 -24534 14630 -24498
rect 14572 -24568 14630 -24534
rect 14572 -24602 14584 -24568
rect 14618 -24602 14630 -24568
rect 14572 -24616 14630 -24602
rect 14854 -24430 14912 -24416
rect 14854 -24464 14866 -24430
rect 14900 -24464 14912 -24430
rect 14854 -24498 14912 -24464
rect 14854 -24534 14866 -24498
rect 14900 -24534 14912 -24498
rect 14854 -24568 14912 -24534
rect 14854 -24602 14866 -24568
rect 14900 -24602 14912 -24568
rect 14854 -24616 14912 -24602
rect 15112 -24430 15170 -24416
rect 15112 -24464 15124 -24430
rect 15158 -24464 15170 -24430
rect 15112 -24498 15170 -24464
rect 15112 -24534 15124 -24498
rect 15158 -24534 15170 -24498
rect 15112 -24568 15170 -24534
rect 15112 -24602 15124 -24568
rect 15158 -24602 15170 -24568
rect 15112 -24616 15170 -24602
rect 15334 -24430 15392 -24416
rect 15334 -24464 15346 -24430
rect 15380 -24464 15392 -24430
rect 15334 -24498 15392 -24464
rect 15334 -24534 15346 -24498
rect 15380 -24534 15392 -24498
rect 15334 -24568 15392 -24534
rect 15334 -24602 15346 -24568
rect 15380 -24602 15392 -24568
rect 15334 -24616 15392 -24602
rect 15592 -24430 15650 -24416
rect 15592 -24464 15604 -24430
rect 15638 -24464 15650 -24430
rect 15592 -24498 15650 -24464
rect 15592 -24534 15604 -24498
rect 15638 -24534 15650 -24498
rect 15592 -24568 15650 -24534
rect 15592 -24602 15604 -24568
rect 15638 -24602 15650 -24568
rect 15592 -24616 15650 -24602
rect 15837 -24428 15895 -24414
rect 15837 -24462 15849 -24428
rect 15883 -24462 15895 -24428
rect 15837 -24496 15895 -24462
rect 15837 -24532 15849 -24496
rect 15883 -24532 15895 -24496
rect 15837 -24566 15895 -24532
rect 15837 -24600 15849 -24566
rect 15883 -24600 15895 -24566
rect 15837 -24614 15895 -24600
rect 16095 -24428 16153 -24414
rect 16095 -24462 16107 -24428
rect 16141 -24462 16153 -24428
rect 16095 -24496 16153 -24462
rect 16095 -24532 16107 -24496
rect 16141 -24532 16153 -24496
rect 16095 -24566 16153 -24532
rect 16095 -24600 16107 -24566
rect 16141 -24600 16153 -24566
rect 16095 -24614 16153 -24600
rect 16347 -24418 16405 -24404
rect 16347 -24452 16359 -24418
rect 16393 -24452 16405 -24418
rect 16347 -24486 16405 -24452
rect 16347 -24522 16359 -24486
rect 16393 -24522 16405 -24486
rect 16347 -24556 16405 -24522
rect 16347 -24590 16359 -24556
rect 16393 -24590 16405 -24556
rect 16347 -24604 16405 -24590
rect 16605 -24418 16663 -24404
rect 16605 -24452 16617 -24418
rect 16651 -24452 16663 -24418
rect 16605 -24486 16663 -24452
rect 16605 -24522 16617 -24486
rect 16651 -24522 16663 -24486
rect 16605 -24556 16663 -24522
rect 16605 -24590 16617 -24556
rect 16651 -24590 16663 -24556
rect 16605 -24604 16663 -24590
rect 17978 -7634 18036 -7622
rect 17978 -9010 17990 -7634
rect 18024 -9010 18036 -7634
rect 17978 -9022 18036 -9010
rect 19636 -7634 19694 -7622
rect 19636 -9010 19648 -7634
rect 19682 -9010 19694 -7634
rect 19636 -9022 19694 -9010
rect 21294 -7634 21352 -7622
rect 21294 -9010 21306 -7634
rect 21340 -9010 21352 -7634
rect 21294 -9022 21352 -9010
rect 17978 -9144 18036 -9132
rect 17978 -10520 17990 -9144
rect 18024 -10520 18036 -9144
rect 17978 -10532 18036 -10520
rect 19636 -9144 19694 -9132
rect 19636 -10520 19648 -9144
rect 19682 -10520 19694 -9144
rect 19636 -10532 19694 -10520
rect 21294 -9144 21352 -9132
rect 21294 -10520 21306 -9144
rect 21340 -10520 21352 -9144
rect 21294 -10532 21352 -10520
rect 17978 -10654 18036 -10642
rect 17978 -12030 17990 -10654
rect 18024 -12030 18036 -10654
rect 17978 -12042 18036 -12030
rect 19636 -10654 19694 -10642
rect 19636 -12030 19648 -10654
rect 19682 -12030 19694 -10654
rect 19636 -12042 19694 -12030
rect 21294 -10654 21352 -10642
rect 21294 -12030 21306 -10654
rect 21340 -12030 21352 -10654
rect 21294 -12042 21352 -12030
rect 17978 -12164 18036 -12152
rect 17978 -13540 17990 -12164
rect 18024 -13540 18036 -12164
rect 17978 -13552 18036 -13540
rect 19636 -12164 19694 -12152
rect 19636 -13540 19648 -12164
rect 19682 -13540 19694 -12164
rect 19636 -13552 19694 -13540
rect 21294 -12164 21352 -12152
rect 21294 -13540 21306 -12164
rect 21340 -13540 21352 -12164
rect 21294 -13552 21352 -13540
rect 17978 -13674 18036 -13662
rect 17978 -15050 17990 -13674
rect 18024 -15050 18036 -13674
rect 17978 -15062 18036 -15050
rect 19636 -13674 19694 -13662
rect 19636 -15050 19648 -13674
rect 19682 -15050 19694 -13674
rect 19636 -15062 19694 -15050
rect 21294 -13674 21352 -13662
rect 21294 -15050 21306 -13674
rect 21340 -15050 21352 -13674
rect 21294 -15062 21352 -15050
rect 17978 -15184 18036 -15172
rect 17978 -16560 17990 -15184
rect 18024 -16560 18036 -15184
rect 17978 -16572 18036 -16560
rect 19636 -15184 19694 -15172
rect 19636 -16560 19648 -15184
rect 19682 -16560 19694 -15184
rect 19636 -16572 19694 -16560
rect 21294 -15184 21352 -15172
rect 21294 -16560 21306 -15184
rect 21340 -16560 21352 -15184
rect 21294 -16572 21352 -16560
rect 17978 -16694 18036 -16682
rect 17978 -18070 17990 -16694
rect 18024 -18070 18036 -16694
rect 17978 -18082 18036 -18070
rect 19636 -16694 19694 -16682
rect 19636 -18070 19648 -16694
rect 19682 -18070 19694 -16694
rect 19636 -18082 19694 -18070
rect 21294 -16694 21352 -16682
rect 21294 -18070 21306 -16694
rect 21340 -18070 21352 -16694
rect 21294 -18082 21352 -18070
rect 17978 -18204 18036 -18192
rect 17978 -19580 17990 -18204
rect 18024 -19580 18036 -18204
rect 17978 -19592 18036 -19580
rect 19636 -18204 19694 -18192
rect 19636 -19580 19648 -18204
rect 19682 -19580 19694 -18204
rect 19636 -19592 19694 -19580
rect 21294 -18204 21352 -18192
rect 21294 -19580 21306 -18204
rect 21340 -19580 21352 -18204
rect 21294 -19592 21352 -19580
rect 17978 -19714 18036 -19702
rect 17978 -21090 17990 -19714
rect 18024 -21090 18036 -19714
rect 17978 -21102 18036 -21090
rect 19636 -19714 19694 -19702
rect 19636 -21090 19648 -19714
rect 19682 -21090 19694 -19714
rect 19636 -21102 19694 -21090
rect 21294 -19714 21352 -19702
rect 21294 -21090 21306 -19714
rect 21340 -21090 21352 -19714
rect 21294 -21102 21352 -21090
rect 17978 -21224 18036 -21212
rect 17978 -22600 17990 -21224
rect 18024 -22600 18036 -21224
rect 17978 -22612 18036 -22600
rect 19636 -21224 19694 -21212
rect 19636 -22600 19648 -21224
rect 19682 -22600 19694 -21224
rect 19636 -22612 19694 -22600
rect 21294 -21224 21352 -21212
rect 21294 -22600 21306 -21224
rect 21340 -22600 21352 -21224
rect 21294 -22612 21352 -22600
rect 17978 -22734 18036 -22722
rect 17978 -24110 17990 -22734
rect 18024 -24110 18036 -22734
rect 17978 -24122 18036 -24110
rect 19636 -22734 19694 -22722
rect 19636 -24110 19648 -22734
rect 19682 -24110 19694 -22734
rect 19636 -24122 19694 -24110
rect 21294 -22734 21352 -22722
rect 21294 -24110 21306 -22734
rect 21340 -24110 21352 -22734
rect 21294 -24122 21352 -24110
rect 17978 -24244 18036 -24232
rect 17978 -25620 17990 -24244
rect 18024 -25620 18036 -24244
rect 17978 -25632 18036 -25620
rect 19636 -24244 19694 -24232
rect 19636 -25620 19648 -24244
rect 19682 -25620 19694 -24244
rect 19636 -25632 19694 -25620
rect 21294 -24244 21352 -24232
rect 21294 -25620 21306 -24244
rect 21340 -25620 21352 -24244
rect 21294 -25632 21352 -25620
<< pdiff >>
rect -94622 20212 -94564 20568
rect -94622 19524 -94610 20212
rect -94576 19524 -94564 20212
rect -94622 19168 -94564 19524
rect -92964 20212 -92906 20568
rect -92964 19524 -92952 20212
rect -92918 19524 -92906 20212
rect -92964 19168 -92906 19524
rect -91306 20212 -91248 20568
rect -91306 19524 -91294 20212
rect -91260 19524 -91248 20212
rect -91306 19168 -91248 19524
rect -89648 20212 -89590 20568
rect -89648 19524 -89636 20212
rect -89602 19524 -89590 20212
rect -89648 19168 -89590 19524
rect -87990 20212 -87932 20568
rect -87990 19524 -87978 20212
rect -87944 19524 -87932 20212
rect -87990 19168 -87932 19524
rect -86332 20212 -86274 20568
rect -86332 19524 -86320 20212
rect -86286 19524 -86274 20212
rect -86332 19168 -86274 19524
rect -84674 20212 -84616 20568
rect -84674 19524 -84662 20212
rect -84628 19524 -84616 20212
rect -84674 19168 -84616 19524
rect -83016 20212 -82958 20568
rect -83016 19524 -83004 20212
rect -82970 19524 -82958 20212
rect -83016 19168 -82958 19524
rect -81358 20212 -81300 20568
rect -81358 19524 -81346 20212
rect -81312 19524 -81300 20212
rect -81358 19168 -81300 19524
rect -79700 20212 -79642 20568
rect -79700 19524 -79688 20212
rect -79654 19524 -79642 20212
rect -79700 19168 -79642 19524
rect -78042 20212 -77984 20568
rect -78042 19524 -78030 20212
rect -77996 19524 -77984 20212
rect -78042 19168 -77984 19524
rect -76384 20212 -76326 20568
rect -76384 19524 -76372 20212
rect -76338 19524 -76326 20212
rect -76384 19168 -76326 19524
rect -74726 20212 -74668 20568
rect -74726 19524 -74714 20212
rect -74680 19524 -74668 20212
rect -74726 19168 -74668 19524
rect -73068 20212 -73010 20568
rect -73068 19524 -73056 20212
rect -73022 19524 -73010 20212
rect -73068 19168 -73010 19524
rect -71410 20212 -71352 20568
rect -71410 19524 -71398 20212
rect -71364 19524 -71352 20212
rect -71410 19168 -71352 19524
rect -69752 20212 -69694 20568
rect -69752 19524 -69740 20212
rect -69706 19524 -69694 20212
rect -69752 19168 -69694 19524
rect -68094 20212 -68036 20568
rect -68094 19524 -68082 20212
rect -68048 19524 -68036 20212
rect -68094 19168 -68036 19524
rect -66436 20212 -66378 20568
rect -66436 19524 -66424 20212
rect -66390 19524 -66378 20212
rect -66436 19168 -66378 19524
rect -64778 20212 -64720 20568
rect -64778 19524 -64766 20212
rect -64732 19524 -64720 20212
rect -64778 19168 -64720 19524
rect -63120 20212 -63062 20568
rect -63120 19524 -63108 20212
rect -63074 19524 -63062 20212
rect -63120 19168 -63062 19524
rect -61462 20212 -61404 20568
rect -61462 19524 -61450 20212
rect -61416 19524 -61404 20212
rect -61462 19168 -61404 19524
rect -59804 20212 -59746 20568
rect -59804 19524 -59792 20212
rect -59758 19524 -59746 20212
rect -59804 19168 -59746 19524
rect -58146 20212 -58088 20568
rect -58146 19524 -58134 20212
rect -58100 19524 -58088 20212
rect -58146 19168 -58088 19524
rect -56488 20212 -56430 20568
rect -56488 19524 -56476 20212
rect -56442 19524 -56430 20212
rect -56488 19168 -56430 19524
rect -54830 20212 -54772 20568
rect -54830 19524 -54818 20212
rect -54784 19524 -54772 20212
rect -54830 19168 -54772 19524
rect -53172 20212 -53114 20568
rect -53172 19524 -53160 20212
rect -53126 19524 -53114 20212
rect -53172 19168 -53114 19524
rect -51514 20212 -51456 20568
rect -51514 19524 -51502 20212
rect -51468 19524 -51456 20212
rect -51514 19168 -51456 19524
rect -49856 20212 -49798 20568
rect -49856 19524 -49844 20212
rect -49810 19524 -49798 20212
rect -49856 19168 -49798 19524
rect -48198 20212 -48140 20568
rect -48198 19524 -48186 20212
rect -48152 19524 -48140 20212
rect -48198 19168 -48140 19524
rect -46540 20212 -46482 20568
rect -46540 19524 -46528 20212
rect -46494 19524 -46482 20212
rect -46540 19168 -46482 19524
rect -44882 20212 -44824 20568
rect -44882 19524 -44870 20212
rect -44836 19524 -44824 20212
rect -44882 19168 -44824 19524
rect -43224 20212 -43166 20568
rect -43224 19524 -43212 20212
rect -43178 19524 -43166 20212
rect -43224 19168 -43166 19524
rect -41566 20212 -41508 20568
rect -41566 19524 -41554 20212
rect -41520 19524 -41508 20212
rect -41566 19168 -41508 19524
rect -39908 20212 -39850 20568
rect -39908 19524 -39896 20212
rect -39862 19524 -39850 20212
rect -39908 19168 -39850 19524
rect -38250 20212 -38192 20568
rect -38250 19524 -38238 20212
rect -38204 19524 -38192 20212
rect -38250 19168 -38192 19524
rect -36592 20212 -36534 20568
rect -36592 19524 -36580 20212
rect -36546 19524 -36534 20212
rect -36592 19168 -36534 19524
rect -34934 20212 -34876 20568
rect -34934 19524 -34922 20212
rect -34888 19524 -34876 20212
rect -34934 19168 -34876 19524
rect -33276 20212 -33218 20568
rect -33276 19524 -33264 20212
rect -33230 19524 -33218 20212
rect -33276 19168 -33218 19524
rect -31618 20212 -31560 20568
rect -31618 19524 -31606 20212
rect -31572 19524 -31560 20212
rect -31618 19168 -31560 19524
rect -29960 20212 -29902 20568
rect -29960 19524 -29948 20212
rect -29914 19524 -29902 20212
rect -29960 19168 -29902 19524
rect -28302 20212 -28244 20568
rect -28302 19524 -28290 20212
rect -28256 19524 -28244 20212
rect -28302 19168 -28244 19524
rect -94622 18576 -94564 18932
rect -94622 17888 -94610 18576
rect -94576 17888 -94564 18576
rect -94622 17532 -94564 17888
rect -92964 18576 -92906 18932
rect -92964 17888 -92952 18576
rect -92918 17888 -92906 18576
rect -92964 17532 -92906 17888
rect -91306 18576 -91248 18932
rect -91306 17888 -91294 18576
rect -91260 17888 -91248 18576
rect -91306 17532 -91248 17888
rect -89648 18576 -89590 18932
rect -89648 17888 -89636 18576
rect -89602 17888 -89590 18576
rect -89648 17532 -89590 17888
rect -87990 18576 -87932 18932
rect -87990 17888 -87978 18576
rect -87944 17888 -87932 18576
rect -87990 17532 -87932 17888
rect -86332 18576 -86274 18932
rect -86332 17888 -86320 18576
rect -86286 17888 -86274 18576
rect -86332 17532 -86274 17888
rect -84674 18576 -84616 18932
rect -84674 17888 -84662 18576
rect -84628 17888 -84616 18576
rect -84674 17532 -84616 17888
rect -83016 18576 -82958 18932
rect -83016 17888 -83004 18576
rect -82970 17888 -82958 18576
rect -83016 17532 -82958 17888
rect -81358 18576 -81300 18932
rect -81358 17888 -81346 18576
rect -81312 17888 -81300 18576
rect -81358 17532 -81300 17888
rect -79700 18576 -79642 18932
rect -79700 17888 -79688 18576
rect -79654 17888 -79642 18576
rect -79700 17532 -79642 17888
rect -78042 18576 -77984 18932
rect -78042 17888 -78030 18576
rect -77996 17888 -77984 18576
rect -78042 17532 -77984 17888
rect -76384 18576 -76326 18932
rect -76384 17888 -76372 18576
rect -76338 17888 -76326 18576
rect -76384 17532 -76326 17888
rect -74726 18576 -74668 18932
rect -74726 17888 -74714 18576
rect -74680 17888 -74668 18576
rect -74726 17532 -74668 17888
rect -73068 18576 -73010 18932
rect -73068 17888 -73056 18576
rect -73022 17888 -73010 18576
rect -73068 17532 -73010 17888
rect -71410 18576 -71352 18932
rect -71410 17888 -71398 18576
rect -71364 17888 -71352 18576
rect -71410 17532 -71352 17888
rect -69752 18576 -69694 18932
rect -69752 17888 -69740 18576
rect -69706 17888 -69694 18576
rect -69752 17532 -69694 17888
rect -68094 18576 -68036 18932
rect -68094 17888 -68082 18576
rect -68048 17888 -68036 18576
rect -68094 17532 -68036 17888
rect -66436 18576 -66378 18932
rect -66436 17888 -66424 18576
rect -66390 17888 -66378 18576
rect -66436 17532 -66378 17888
rect -64778 18576 -64720 18932
rect -64778 17888 -64766 18576
rect -64732 17888 -64720 18576
rect -64778 17532 -64720 17888
rect -63120 18576 -63062 18932
rect -63120 17888 -63108 18576
rect -63074 17888 -63062 18576
rect -63120 17532 -63062 17888
rect -61462 18576 -61404 18932
rect -61462 17888 -61450 18576
rect -61416 17888 -61404 18576
rect -61462 17532 -61404 17888
rect -59804 18576 -59746 18932
rect -59804 17888 -59792 18576
rect -59758 17888 -59746 18576
rect -59804 17532 -59746 17888
rect -58146 18576 -58088 18932
rect -58146 17888 -58134 18576
rect -58100 17888 -58088 18576
rect -58146 17532 -58088 17888
rect -56488 18576 -56430 18932
rect -56488 17888 -56476 18576
rect -56442 17888 -56430 18576
rect -56488 17532 -56430 17888
rect -54830 18576 -54772 18932
rect -54830 17888 -54818 18576
rect -54784 17888 -54772 18576
rect -54830 17532 -54772 17888
rect -53172 18576 -53114 18932
rect -53172 17888 -53160 18576
rect -53126 17888 -53114 18576
rect -53172 17532 -53114 17888
rect -51514 18576 -51456 18932
rect -51514 17888 -51502 18576
rect -51468 17888 -51456 18576
rect -51514 17532 -51456 17888
rect -49856 18576 -49798 18932
rect -49856 17888 -49844 18576
rect -49810 17888 -49798 18576
rect -49856 17532 -49798 17888
rect -48198 18576 -48140 18932
rect -48198 17888 -48186 18576
rect -48152 17888 -48140 18576
rect -48198 17532 -48140 17888
rect -46540 18576 -46482 18932
rect -46540 17888 -46528 18576
rect -46494 17888 -46482 18576
rect -46540 17532 -46482 17888
rect -44882 18576 -44824 18932
rect -44882 17888 -44870 18576
rect -44836 17888 -44824 18576
rect -44882 17532 -44824 17888
rect -43224 18576 -43166 18932
rect -43224 17888 -43212 18576
rect -43178 17888 -43166 18576
rect -43224 17532 -43166 17888
rect -41566 18576 -41508 18932
rect -41566 17888 -41554 18576
rect -41520 17888 -41508 18576
rect -41566 17532 -41508 17888
rect -39908 18576 -39850 18932
rect -39908 17888 -39896 18576
rect -39862 17888 -39850 18576
rect -39908 17532 -39850 17888
rect -38250 18576 -38192 18932
rect -38250 17888 -38238 18576
rect -38204 17888 -38192 18576
rect -38250 17532 -38192 17888
rect -36592 18576 -36534 18932
rect -36592 17888 -36580 18576
rect -36546 17888 -36534 18576
rect -36592 17532 -36534 17888
rect -34934 18576 -34876 18932
rect -34934 17888 -34922 18576
rect -34888 17888 -34876 18576
rect -34934 17532 -34876 17888
rect -33276 18576 -33218 18932
rect -33276 17888 -33264 18576
rect -33230 17888 -33218 18576
rect -33276 17532 -33218 17888
rect -31618 18576 -31560 18932
rect -31618 17888 -31606 18576
rect -31572 17888 -31560 18576
rect -31618 17532 -31560 17888
rect -29960 18576 -29902 18932
rect -29960 17888 -29948 18576
rect -29914 17888 -29902 18576
rect -29960 17532 -29902 17888
rect -28302 18576 -28244 18932
rect -28302 17888 -28290 18576
rect -28256 17888 -28244 18576
rect -28302 17532 -28244 17888
rect -94620 16830 -94562 17186
rect -94620 16142 -94608 16830
rect -94574 16142 -94562 16830
rect -94620 15786 -94562 16142
rect -92962 16830 -92904 17186
rect -92962 16142 -92950 16830
rect -92916 16142 -92904 16830
rect -92962 15786 -92904 16142
rect -91304 16830 -91246 17186
rect -91304 16142 -91292 16830
rect -91258 16142 -91246 16830
rect -91304 15786 -91246 16142
rect -89646 16830 -89588 17186
rect -89646 16142 -89634 16830
rect -89600 16142 -89588 16830
rect -89646 15786 -89588 16142
rect -87988 16830 -87930 17186
rect -87988 16142 -87976 16830
rect -87942 16142 -87930 16830
rect -87988 15786 -87930 16142
rect -86330 16830 -86272 17186
rect -86330 16142 -86318 16830
rect -86284 16142 -86272 16830
rect -86330 15786 -86272 16142
rect -84672 16830 -84614 17186
rect -84672 16142 -84660 16830
rect -84626 16142 -84614 16830
rect -84672 15786 -84614 16142
rect -83014 16830 -82956 17186
rect -83014 16142 -83002 16830
rect -82968 16142 -82956 16830
rect -83014 15786 -82956 16142
rect -81356 16830 -81298 17186
rect -81356 16142 -81344 16830
rect -81310 16142 -81298 16830
rect -81356 15786 -81298 16142
rect -79698 16830 -79640 17186
rect -79698 16142 -79686 16830
rect -79652 16142 -79640 16830
rect -79698 15786 -79640 16142
rect -78040 16830 -77982 17186
rect -78040 16142 -78028 16830
rect -77994 16142 -77982 16830
rect -78040 15786 -77982 16142
rect -76382 16830 -76324 17186
rect -76382 16142 -76370 16830
rect -76336 16142 -76324 16830
rect -76382 15786 -76324 16142
rect -74724 16830 -74666 17186
rect -74724 16142 -74712 16830
rect -74678 16142 -74666 16830
rect -74724 15786 -74666 16142
rect -73066 16830 -73008 17186
rect -73066 16142 -73054 16830
rect -73020 16142 -73008 16830
rect -73066 15786 -73008 16142
rect -71408 16830 -71350 17186
rect -71408 16142 -71396 16830
rect -71362 16142 -71350 16830
rect -71408 15786 -71350 16142
rect -69750 16830 -69692 17186
rect -69750 16142 -69738 16830
rect -69704 16142 -69692 16830
rect -69750 15786 -69692 16142
rect -68092 16830 -68034 17186
rect -68092 16142 -68080 16830
rect -68046 16142 -68034 16830
rect -68092 15786 -68034 16142
rect -66434 16830 -66376 17186
rect -66434 16142 -66422 16830
rect -66388 16142 -66376 16830
rect -66434 15786 -66376 16142
rect -64776 16830 -64718 17186
rect -64776 16142 -64764 16830
rect -64730 16142 -64718 16830
rect -64776 15786 -64718 16142
rect -63118 16830 -63060 17186
rect -63118 16142 -63106 16830
rect -63072 16142 -63060 16830
rect -63118 15786 -63060 16142
rect -61460 16830 -61402 17186
rect -61460 16142 -61448 16830
rect -61414 16142 -61402 16830
rect -61460 15786 -61402 16142
rect -59802 16830 -59744 17186
rect -59802 16142 -59790 16830
rect -59756 16142 -59744 16830
rect -59802 15786 -59744 16142
rect -58144 16830 -58086 17186
rect -58144 16142 -58132 16830
rect -58098 16142 -58086 16830
rect -58144 15786 -58086 16142
rect -56486 16830 -56428 17186
rect -56486 16142 -56474 16830
rect -56440 16142 -56428 16830
rect -56486 15786 -56428 16142
rect -54828 16830 -54770 17186
rect -54828 16142 -54816 16830
rect -54782 16142 -54770 16830
rect -54828 15786 -54770 16142
rect -53170 16830 -53112 17186
rect -53170 16142 -53158 16830
rect -53124 16142 -53112 16830
rect -53170 15786 -53112 16142
rect -51512 16830 -51454 17186
rect -51512 16142 -51500 16830
rect -51466 16142 -51454 16830
rect -51512 15786 -51454 16142
rect -49854 16830 -49796 17186
rect -49854 16142 -49842 16830
rect -49808 16142 -49796 16830
rect -49854 15786 -49796 16142
rect -48196 16830 -48138 17186
rect -48196 16142 -48184 16830
rect -48150 16142 -48138 16830
rect -48196 15786 -48138 16142
rect -46538 16830 -46480 17186
rect -46538 16142 -46526 16830
rect -46492 16142 -46480 16830
rect -46538 15786 -46480 16142
rect -44880 16830 -44822 17186
rect -44880 16142 -44868 16830
rect -44834 16142 -44822 16830
rect -44880 15786 -44822 16142
rect -43222 16830 -43164 17186
rect -43222 16142 -43210 16830
rect -43176 16142 -43164 16830
rect -43222 15786 -43164 16142
rect -41564 16830 -41506 17186
rect -41564 16142 -41552 16830
rect -41518 16142 -41506 16830
rect -41564 15786 -41506 16142
rect -39906 16830 -39848 17186
rect -39906 16142 -39894 16830
rect -39860 16142 -39848 16830
rect -39906 15786 -39848 16142
rect -38248 16830 -38190 17186
rect -38248 16142 -38236 16830
rect -38202 16142 -38190 16830
rect -38248 15786 -38190 16142
rect -36590 16830 -36532 17186
rect -36590 16142 -36578 16830
rect -36544 16142 -36532 16830
rect -36590 15786 -36532 16142
rect -34932 16830 -34874 17186
rect -34932 16142 -34920 16830
rect -34886 16142 -34874 16830
rect -34932 15786 -34874 16142
rect -33274 16830 -33216 17186
rect -33274 16142 -33262 16830
rect -33228 16142 -33216 16830
rect -33274 15786 -33216 16142
rect -31616 16830 -31558 17186
rect -31616 16142 -31604 16830
rect -31570 16142 -31558 16830
rect -31616 15786 -31558 16142
rect -29958 16830 -29900 17186
rect -29958 16142 -29946 16830
rect -29912 16142 -29900 16830
rect -29958 15786 -29900 16142
rect -28300 16830 -28242 17186
rect -28300 16142 -28288 16830
rect -28254 16142 -28242 16830
rect -28300 15786 -28242 16142
rect -94620 15194 -94562 15550
rect -94620 14506 -94608 15194
rect -94574 14506 -94562 15194
rect -94620 14150 -94562 14506
rect -92962 15194 -92904 15550
rect -92962 14506 -92950 15194
rect -92916 14506 -92904 15194
rect -92962 14150 -92904 14506
rect -91304 15194 -91246 15550
rect -91304 14506 -91292 15194
rect -91258 14506 -91246 15194
rect -91304 14150 -91246 14506
rect -89646 15194 -89588 15550
rect -89646 14506 -89634 15194
rect -89600 14506 -89588 15194
rect -89646 14150 -89588 14506
rect -87988 15194 -87930 15550
rect -87988 14506 -87976 15194
rect -87942 14506 -87930 15194
rect -87988 14150 -87930 14506
rect -86330 15194 -86272 15550
rect -86330 14506 -86318 15194
rect -86284 14506 -86272 15194
rect -86330 14150 -86272 14506
rect -84672 15194 -84614 15550
rect -84672 14506 -84660 15194
rect -84626 14506 -84614 15194
rect -84672 14150 -84614 14506
rect -83014 15194 -82956 15550
rect -83014 14506 -83002 15194
rect -82968 14506 -82956 15194
rect -83014 14150 -82956 14506
rect -81356 15194 -81298 15550
rect -81356 14506 -81344 15194
rect -81310 14506 -81298 15194
rect -81356 14150 -81298 14506
rect -79698 15194 -79640 15550
rect -79698 14506 -79686 15194
rect -79652 14506 -79640 15194
rect -79698 14150 -79640 14506
rect -78040 15194 -77982 15550
rect -78040 14506 -78028 15194
rect -77994 14506 -77982 15194
rect -78040 14150 -77982 14506
rect -76382 15194 -76324 15550
rect -76382 14506 -76370 15194
rect -76336 14506 -76324 15194
rect -76382 14150 -76324 14506
rect -74724 15194 -74666 15550
rect -74724 14506 -74712 15194
rect -74678 14506 -74666 15194
rect -74724 14150 -74666 14506
rect -73066 15194 -73008 15550
rect -73066 14506 -73054 15194
rect -73020 14506 -73008 15194
rect -73066 14150 -73008 14506
rect -71408 15194 -71350 15550
rect -71408 14506 -71396 15194
rect -71362 14506 -71350 15194
rect -71408 14150 -71350 14506
rect -69750 15194 -69692 15550
rect -69750 14506 -69738 15194
rect -69704 14506 -69692 15194
rect -69750 14150 -69692 14506
rect -68092 15194 -68034 15550
rect -68092 14506 -68080 15194
rect -68046 14506 -68034 15194
rect -68092 14150 -68034 14506
rect -66434 15194 -66376 15550
rect -66434 14506 -66422 15194
rect -66388 14506 -66376 15194
rect -66434 14150 -66376 14506
rect -64776 15194 -64718 15550
rect -64776 14506 -64764 15194
rect -64730 14506 -64718 15194
rect -64776 14150 -64718 14506
rect -63118 15194 -63060 15550
rect -63118 14506 -63106 15194
rect -63072 14506 -63060 15194
rect -63118 14150 -63060 14506
rect -61460 15194 -61402 15550
rect -61460 14506 -61448 15194
rect -61414 14506 -61402 15194
rect -61460 14150 -61402 14506
rect -59802 15194 -59744 15550
rect -59802 14506 -59790 15194
rect -59756 14506 -59744 15194
rect -59802 14150 -59744 14506
rect -58144 15194 -58086 15550
rect -58144 14506 -58132 15194
rect -58098 14506 -58086 15194
rect -58144 14150 -58086 14506
rect -56486 15194 -56428 15550
rect -56486 14506 -56474 15194
rect -56440 14506 -56428 15194
rect -56486 14150 -56428 14506
rect -54828 15194 -54770 15550
rect -54828 14506 -54816 15194
rect -54782 14506 -54770 15194
rect -54828 14150 -54770 14506
rect -53170 15194 -53112 15550
rect -53170 14506 -53158 15194
rect -53124 14506 -53112 15194
rect -53170 14150 -53112 14506
rect -51512 15194 -51454 15550
rect -51512 14506 -51500 15194
rect -51466 14506 -51454 15194
rect -51512 14150 -51454 14506
rect -49854 15194 -49796 15550
rect -49854 14506 -49842 15194
rect -49808 14506 -49796 15194
rect -49854 14150 -49796 14506
rect -48196 15194 -48138 15550
rect -48196 14506 -48184 15194
rect -48150 14506 -48138 15194
rect -48196 14150 -48138 14506
rect -46538 15194 -46480 15550
rect -46538 14506 -46526 15194
rect -46492 14506 -46480 15194
rect -46538 14150 -46480 14506
rect -44880 15194 -44822 15550
rect -44880 14506 -44868 15194
rect -44834 14506 -44822 15194
rect -44880 14150 -44822 14506
rect -43222 15194 -43164 15550
rect -43222 14506 -43210 15194
rect -43176 14506 -43164 15194
rect -43222 14150 -43164 14506
rect -41564 15194 -41506 15550
rect -41564 14506 -41552 15194
rect -41518 14506 -41506 15194
rect -41564 14150 -41506 14506
rect -39906 15194 -39848 15550
rect -39906 14506 -39894 15194
rect -39860 14506 -39848 15194
rect -39906 14150 -39848 14506
rect -38248 15194 -38190 15550
rect -38248 14506 -38236 15194
rect -38202 14506 -38190 15194
rect -38248 14150 -38190 14506
rect -36590 15194 -36532 15550
rect -36590 14506 -36578 15194
rect -36544 14506 -36532 15194
rect -36590 14150 -36532 14506
rect -34932 15194 -34874 15550
rect -34932 14506 -34920 15194
rect -34886 14506 -34874 15194
rect -34932 14150 -34874 14506
rect -33274 15194 -33216 15550
rect -33274 14506 -33262 15194
rect -33228 14506 -33216 15194
rect -33274 14150 -33216 14506
rect -31616 15194 -31558 15550
rect -31616 14506 -31604 15194
rect -31570 14506 -31558 15194
rect -31616 14150 -31558 14506
rect -29958 15194 -29900 15550
rect -29958 14506 -29946 15194
rect -29912 14506 -29900 15194
rect -29958 14150 -29900 14506
rect -28300 15194 -28242 15550
rect -28300 14506 -28288 15194
rect -28254 14506 -28242 15194
rect -28300 14150 -28242 14506
rect -94620 13558 -94562 13914
rect -94620 12870 -94608 13558
rect -94574 12870 -94562 13558
rect -94620 12514 -94562 12870
rect -92962 13558 -92904 13914
rect -92962 12870 -92950 13558
rect -92916 12870 -92904 13558
rect -92962 12514 -92904 12870
rect -91304 13558 -91246 13914
rect -91304 12870 -91292 13558
rect -91258 12870 -91246 13558
rect -91304 12514 -91246 12870
rect -89646 13558 -89588 13914
rect -89646 12870 -89634 13558
rect -89600 12870 -89588 13558
rect -89646 12514 -89588 12870
rect -87988 13558 -87930 13914
rect -87988 12870 -87976 13558
rect -87942 12870 -87930 13558
rect -87988 12514 -87930 12870
rect -86330 13558 -86272 13914
rect -86330 12870 -86318 13558
rect -86284 12870 -86272 13558
rect -86330 12514 -86272 12870
rect -84672 13558 -84614 13914
rect -84672 12870 -84660 13558
rect -84626 12870 -84614 13558
rect -84672 12514 -84614 12870
rect -83014 13558 -82956 13914
rect -83014 12870 -83002 13558
rect -82968 12870 -82956 13558
rect -83014 12514 -82956 12870
rect -81356 13558 -81298 13914
rect -81356 12870 -81344 13558
rect -81310 12870 -81298 13558
rect -81356 12514 -81298 12870
rect -79698 13558 -79640 13914
rect -79698 12870 -79686 13558
rect -79652 12870 -79640 13558
rect -79698 12514 -79640 12870
rect -78040 13558 -77982 13914
rect -78040 12870 -78028 13558
rect -77994 12870 -77982 13558
rect -78040 12514 -77982 12870
rect -76382 13558 -76324 13914
rect -76382 12870 -76370 13558
rect -76336 12870 -76324 13558
rect -76382 12514 -76324 12870
rect -74724 13558 -74666 13914
rect -74724 12870 -74712 13558
rect -74678 12870 -74666 13558
rect -74724 12514 -74666 12870
rect -73066 13558 -73008 13914
rect -73066 12870 -73054 13558
rect -73020 12870 -73008 13558
rect -73066 12514 -73008 12870
rect -71408 13558 -71350 13914
rect -71408 12870 -71396 13558
rect -71362 12870 -71350 13558
rect -71408 12514 -71350 12870
rect -69750 13558 -69692 13914
rect -69750 12870 -69738 13558
rect -69704 12870 -69692 13558
rect -69750 12514 -69692 12870
rect -68092 13558 -68034 13914
rect -68092 12870 -68080 13558
rect -68046 12870 -68034 13558
rect -68092 12514 -68034 12870
rect -66434 13558 -66376 13914
rect -66434 12870 -66422 13558
rect -66388 12870 -66376 13558
rect -66434 12514 -66376 12870
rect -64776 13558 -64718 13914
rect -64776 12870 -64764 13558
rect -64730 12870 -64718 13558
rect -64776 12514 -64718 12870
rect -63118 13558 -63060 13914
rect -63118 12870 -63106 13558
rect -63072 12870 -63060 13558
rect -63118 12514 -63060 12870
rect -61460 13558 -61402 13914
rect -61460 12870 -61448 13558
rect -61414 12870 -61402 13558
rect -61460 12514 -61402 12870
rect -59802 13558 -59744 13914
rect -59802 12870 -59790 13558
rect -59756 12870 -59744 13558
rect -59802 12514 -59744 12870
rect -58144 13558 -58086 13914
rect -58144 12870 -58132 13558
rect -58098 12870 -58086 13558
rect -58144 12514 -58086 12870
rect -56486 13558 -56428 13914
rect -56486 12870 -56474 13558
rect -56440 12870 -56428 13558
rect -56486 12514 -56428 12870
rect -54828 13558 -54770 13914
rect -54828 12870 -54816 13558
rect -54782 12870 -54770 13558
rect -54828 12514 -54770 12870
rect -53170 13558 -53112 13914
rect -53170 12870 -53158 13558
rect -53124 12870 -53112 13558
rect -53170 12514 -53112 12870
rect -51512 13558 -51454 13914
rect -51512 12870 -51500 13558
rect -51466 12870 -51454 13558
rect -51512 12514 -51454 12870
rect -49854 13558 -49796 13914
rect -49854 12870 -49842 13558
rect -49808 12870 -49796 13558
rect -49854 12514 -49796 12870
rect -48196 13558 -48138 13914
rect -48196 12870 -48184 13558
rect -48150 12870 -48138 13558
rect -48196 12514 -48138 12870
rect -46538 13558 -46480 13914
rect -46538 12870 -46526 13558
rect -46492 12870 -46480 13558
rect -46538 12514 -46480 12870
rect -44880 13558 -44822 13914
rect -44880 12870 -44868 13558
rect -44834 12870 -44822 13558
rect -44880 12514 -44822 12870
rect -43222 13558 -43164 13914
rect -43222 12870 -43210 13558
rect -43176 12870 -43164 13558
rect -43222 12514 -43164 12870
rect -41564 13558 -41506 13914
rect -41564 12870 -41552 13558
rect -41518 12870 -41506 13558
rect -41564 12514 -41506 12870
rect -39906 13558 -39848 13914
rect -39906 12870 -39894 13558
rect -39860 12870 -39848 13558
rect -39906 12514 -39848 12870
rect -38248 13558 -38190 13914
rect -38248 12870 -38236 13558
rect -38202 12870 -38190 13558
rect -38248 12514 -38190 12870
rect -36590 13558 -36532 13914
rect -36590 12870 -36578 13558
rect -36544 12870 -36532 13558
rect -36590 12514 -36532 12870
rect -34932 13558 -34874 13914
rect -34932 12870 -34920 13558
rect -34886 12870 -34874 13558
rect -34932 12514 -34874 12870
rect -33274 13558 -33216 13914
rect -33274 12870 -33262 13558
rect -33228 12870 -33216 13558
rect -33274 12514 -33216 12870
rect -31616 13558 -31558 13914
rect -31616 12870 -31604 13558
rect -31570 12870 -31558 13558
rect -31616 12514 -31558 12870
rect -29958 13558 -29900 13914
rect -29958 12870 -29946 13558
rect -29912 12870 -29900 13558
rect -29958 12514 -29900 12870
rect -28300 13558 -28242 13914
rect -28300 12870 -28288 13558
rect -28254 12870 -28242 13558
rect -28300 12514 -28242 12870
rect -94620 11922 -94562 12278
rect -94620 11234 -94608 11922
rect -94574 11234 -94562 11922
rect -94620 10878 -94562 11234
rect -92962 11922 -92904 12278
rect -92962 11234 -92950 11922
rect -92916 11234 -92904 11922
rect -92962 10878 -92904 11234
rect -91304 11922 -91246 12278
rect -91304 11234 -91292 11922
rect -91258 11234 -91246 11922
rect -91304 10878 -91246 11234
rect -89646 11922 -89588 12278
rect -89646 11234 -89634 11922
rect -89600 11234 -89588 11922
rect -89646 10878 -89588 11234
rect -87988 11922 -87930 12278
rect -87988 11234 -87976 11922
rect -87942 11234 -87930 11922
rect -87988 10878 -87930 11234
rect -86330 11922 -86272 12278
rect -86330 11234 -86318 11922
rect -86284 11234 -86272 11922
rect -86330 10878 -86272 11234
rect -84672 11922 -84614 12278
rect -84672 11234 -84660 11922
rect -84626 11234 -84614 11922
rect -84672 10878 -84614 11234
rect -83014 11922 -82956 12278
rect -83014 11234 -83002 11922
rect -82968 11234 -82956 11922
rect -83014 10878 -82956 11234
rect -81356 11922 -81298 12278
rect -81356 11234 -81344 11922
rect -81310 11234 -81298 11922
rect -81356 10878 -81298 11234
rect -79698 11922 -79640 12278
rect -79698 11234 -79686 11922
rect -79652 11234 -79640 11922
rect -79698 10878 -79640 11234
rect -78040 11922 -77982 12278
rect -78040 11234 -78028 11922
rect -77994 11234 -77982 11922
rect -78040 10878 -77982 11234
rect -76382 11922 -76324 12278
rect -76382 11234 -76370 11922
rect -76336 11234 -76324 11922
rect -76382 10878 -76324 11234
rect -74724 11922 -74666 12278
rect -74724 11234 -74712 11922
rect -74678 11234 -74666 11922
rect -74724 10878 -74666 11234
rect -73066 11922 -73008 12278
rect -73066 11234 -73054 11922
rect -73020 11234 -73008 11922
rect -73066 10878 -73008 11234
rect -71408 11922 -71350 12278
rect -71408 11234 -71396 11922
rect -71362 11234 -71350 11922
rect -71408 10878 -71350 11234
rect -69750 11922 -69692 12278
rect -69750 11234 -69738 11922
rect -69704 11234 -69692 11922
rect -69750 10878 -69692 11234
rect -68092 11922 -68034 12278
rect -68092 11234 -68080 11922
rect -68046 11234 -68034 11922
rect -68092 10878 -68034 11234
rect -66434 11922 -66376 12278
rect -66434 11234 -66422 11922
rect -66388 11234 -66376 11922
rect -66434 10878 -66376 11234
rect -64776 11922 -64718 12278
rect -64776 11234 -64764 11922
rect -64730 11234 -64718 11922
rect -64776 10878 -64718 11234
rect -63118 11922 -63060 12278
rect -63118 11234 -63106 11922
rect -63072 11234 -63060 11922
rect -63118 10878 -63060 11234
rect -61460 11922 -61402 12278
rect -61460 11234 -61448 11922
rect -61414 11234 -61402 11922
rect -61460 10878 -61402 11234
rect -59802 11922 -59744 12278
rect -59802 11234 -59790 11922
rect -59756 11234 -59744 11922
rect -59802 10878 -59744 11234
rect -58144 11922 -58086 12278
rect -58144 11234 -58132 11922
rect -58098 11234 -58086 11922
rect -58144 10878 -58086 11234
rect -56486 11922 -56428 12278
rect -56486 11234 -56474 11922
rect -56440 11234 -56428 11922
rect -56486 10878 -56428 11234
rect -54828 11922 -54770 12278
rect -54828 11234 -54816 11922
rect -54782 11234 -54770 11922
rect -54828 10878 -54770 11234
rect -53170 11922 -53112 12278
rect -53170 11234 -53158 11922
rect -53124 11234 -53112 11922
rect -53170 10878 -53112 11234
rect -51512 11922 -51454 12278
rect -51512 11234 -51500 11922
rect -51466 11234 -51454 11922
rect -51512 10878 -51454 11234
rect -49854 11922 -49796 12278
rect -49854 11234 -49842 11922
rect -49808 11234 -49796 11922
rect -49854 10878 -49796 11234
rect -48196 11922 -48138 12278
rect -48196 11234 -48184 11922
rect -48150 11234 -48138 11922
rect -48196 10878 -48138 11234
rect -46538 11922 -46480 12278
rect -46538 11234 -46526 11922
rect -46492 11234 -46480 11922
rect -46538 10878 -46480 11234
rect -44880 11922 -44822 12278
rect -44880 11234 -44868 11922
rect -44834 11234 -44822 11922
rect -44880 10878 -44822 11234
rect -43222 11922 -43164 12278
rect -43222 11234 -43210 11922
rect -43176 11234 -43164 11922
rect -43222 10878 -43164 11234
rect -41564 11922 -41506 12278
rect -41564 11234 -41552 11922
rect -41518 11234 -41506 11922
rect -41564 10878 -41506 11234
rect -39906 11922 -39848 12278
rect -39906 11234 -39894 11922
rect -39860 11234 -39848 11922
rect -39906 10878 -39848 11234
rect -38248 11922 -38190 12278
rect -38248 11234 -38236 11922
rect -38202 11234 -38190 11922
rect -38248 10878 -38190 11234
rect -36590 11922 -36532 12278
rect -36590 11234 -36578 11922
rect -36544 11234 -36532 11922
rect -36590 10878 -36532 11234
rect -34932 11922 -34874 12278
rect -34932 11234 -34920 11922
rect -34886 11234 -34874 11922
rect -34932 10878 -34874 11234
rect -33274 11922 -33216 12278
rect -33274 11234 -33262 11922
rect -33228 11234 -33216 11922
rect -33274 10878 -33216 11234
rect -31616 11922 -31558 12278
rect -31616 11234 -31604 11922
rect -31570 11234 -31558 11922
rect -31616 10878 -31558 11234
rect -29958 11922 -29900 12278
rect -29958 11234 -29946 11922
rect -29912 11234 -29900 11922
rect -29958 10878 -29900 11234
rect -28300 11922 -28242 12278
rect -28300 11234 -28288 11922
rect -28254 11234 -28242 11922
rect -28300 10878 -28242 11234
rect -94620 10284 -94562 10640
rect -94620 9596 -94608 10284
rect -94574 9596 -94562 10284
rect -94620 9240 -94562 9596
rect -92962 10284 -92904 10640
rect -92962 9596 -92950 10284
rect -92916 9596 -92904 10284
rect -92962 9240 -92904 9596
rect -91304 10284 -91246 10640
rect -91304 9596 -91292 10284
rect -91258 9596 -91246 10284
rect -91304 9240 -91246 9596
rect -89646 10284 -89588 10640
rect -89646 9596 -89634 10284
rect -89600 9596 -89588 10284
rect -89646 9240 -89588 9596
rect -87988 10284 -87930 10640
rect -87988 9596 -87976 10284
rect -87942 9596 -87930 10284
rect -87988 9240 -87930 9596
rect -86330 10284 -86272 10640
rect -86330 9596 -86318 10284
rect -86284 9596 -86272 10284
rect -86330 9240 -86272 9596
rect -84672 10284 -84614 10640
rect -84672 9596 -84660 10284
rect -84626 9596 -84614 10284
rect -84672 9240 -84614 9596
rect -83014 10284 -82956 10640
rect -83014 9596 -83002 10284
rect -82968 9596 -82956 10284
rect -83014 9240 -82956 9596
rect -81356 10284 -81298 10640
rect -81356 9596 -81344 10284
rect -81310 9596 -81298 10284
rect -81356 9240 -81298 9596
rect -79698 10284 -79640 10640
rect -79698 9596 -79686 10284
rect -79652 9596 -79640 10284
rect -79698 9240 -79640 9596
rect -78040 10284 -77982 10640
rect -78040 9596 -78028 10284
rect -77994 9596 -77982 10284
rect -78040 9240 -77982 9596
rect -76382 10284 -76324 10640
rect -76382 9596 -76370 10284
rect -76336 9596 -76324 10284
rect -76382 9240 -76324 9596
rect -74724 10284 -74666 10640
rect -74724 9596 -74712 10284
rect -74678 9596 -74666 10284
rect -74724 9240 -74666 9596
rect -73066 10284 -73008 10640
rect -73066 9596 -73054 10284
rect -73020 9596 -73008 10284
rect -73066 9240 -73008 9596
rect -71408 10284 -71350 10640
rect -71408 9596 -71396 10284
rect -71362 9596 -71350 10284
rect -71408 9240 -71350 9596
rect -69750 10284 -69692 10640
rect -69750 9596 -69738 10284
rect -69704 9596 -69692 10284
rect -69750 9240 -69692 9596
rect -68092 10284 -68034 10640
rect -68092 9596 -68080 10284
rect -68046 9596 -68034 10284
rect -68092 9240 -68034 9596
rect -66434 10284 -66376 10640
rect -66434 9596 -66422 10284
rect -66388 9596 -66376 10284
rect -66434 9240 -66376 9596
rect -64776 10284 -64718 10640
rect -64776 9596 -64764 10284
rect -64730 9596 -64718 10284
rect -64776 9240 -64718 9596
rect -63118 10284 -63060 10640
rect -63118 9596 -63106 10284
rect -63072 9596 -63060 10284
rect -63118 9240 -63060 9596
rect -61460 10284 -61402 10640
rect -61460 9596 -61448 10284
rect -61414 9596 -61402 10284
rect -61460 9240 -61402 9596
rect -59802 10284 -59744 10640
rect -59802 9596 -59790 10284
rect -59756 9596 -59744 10284
rect -59802 9240 -59744 9596
rect -58144 10284 -58086 10640
rect -58144 9596 -58132 10284
rect -58098 9596 -58086 10284
rect -58144 9240 -58086 9596
rect -56486 10284 -56428 10640
rect -56486 9596 -56474 10284
rect -56440 9596 -56428 10284
rect -56486 9240 -56428 9596
rect -54828 10284 -54770 10640
rect -54828 9596 -54816 10284
rect -54782 9596 -54770 10284
rect -54828 9240 -54770 9596
rect -53170 10284 -53112 10640
rect -53170 9596 -53158 10284
rect -53124 9596 -53112 10284
rect -53170 9240 -53112 9596
rect -51512 10284 -51454 10640
rect -51512 9596 -51500 10284
rect -51466 9596 -51454 10284
rect -51512 9240 -51454 9596
rect -49854 10284 -49796 10640
rect -49854 9596 -49842 10284
rect -49808 9596 -49796 10284
rect -49854 9240 -49796 9596
rect -48196 10284 -48138 10640
rect -48196 9596 -48184 10284
rect -48150 9596 -48138 10284
rect -48196 9240 -48138 9596
rect -46538 10284 -46480 10640
rect -46538 9596 -46526 10284
rect -46492 9596 -46480 10284
rect -46538 9240 -46480 9596
rect -44880 10284 -44822 10640
rect -44880 9596 -44868 10284
rect -44834 9596 -44822 10284
rect -44880 9240 -44822 9596
rect -43222 10284 -43164 10640
rect -43222 9596 -43210 10284
rect -43176 9596 -43164 10284
rect -43222 9240 -43164 9596
rect -41564 10284 -41506 10640
rect -41564 9596 -41552 10284
rect -41518 9596 -41506 10284
rect -41564 9240 -41506 9596
rect -39906 10284 -39848 10640
rect -39906 9596 -39894 10284
rect -39860 9596 -39848 10284
rect -39906 9240 -39848 9596
rect -38248 10284 -38190 10640
rect -38248 9596 -38236 10284
rect -38202 9596 -38190 10284
rect -38248 9240 -38190 9596
rect -36590 10284 -36532 10640
rect -36590 9596 -36578 10284
rect -36544 9596 -36532 10284
rect -36590 9240 -36532 9596
rect -34932 10284 -34874 10640
rect -34932 9596 -34920 10284
rect -34886 9596 -34874 10284
rect -34932 9240 -34874 9596
rect -33274 10284 -33216 10640
rect -33274 9596 -33262 10284
rect -33228 9596 -33216 10284
rect -33274 9240 -33216 9596
rect -31616 10284 -31558 10640
rect -31616 9596 -31604 10284
rect -31570 9596 -31558 10284
rect -31616 9240 -31558 9596
rect -29958 10284 -29900 10640
rect -29958 9596 -29946 10284
rect -29912 9596 -29900 10284
rect -29958 9240 -29900 9596
rect -28300 10284 -28242 10640
rect -28300 9596 -28288 10284
rect -28254 9596 -28242 10284
rect -28300 9240 -28242 9596
rect -94620 8648 -94562 9004
rect -94620 7960 -94608 8648
rect -94574 7960 -94562 8648
rect -94620 7604 -94562 7960
rect -92962 8648 -92904 9004
rect -92962 7960 -92950 8648
rect -92916 7960 -92904 8648
rect -92962 7604 -92904 7960
rect -91304 8648 -91246 9004
rect -91304 7960 -91292 8648
rect -91258 7960 -91246 8648
rect -91304 7604 -91246 7960
rect -89646 8648 -89588 9004
rect -89646 7960 -89634 8648
rect -89600 7960 -89588 8648
rect -89646 7604 -89588 7960
rect -87988 8648 -87930 9004
rect -87988 7960 -87976 8648
rect -87942 7960 -87930 8648
rect -87988 7604 -87930 7960
rect -86330 8648 -86272 9004
rect -86330 7960 -86318 8648
rect -86284 7960 -86272 8648
rect -86330 7604 -86272 7960
rect -84672 8648 -84614 9004
rect -84672 7960 -84660 8648
rect -84626 7960 -84614 8648
rect -84672 7604 -84614 7960
rect -83014 8648 -82956 9004
rect -83014 7960 -83002 8648
rect -82968 7960 -82956 8648
rect -83014 7604 -82956 7960
rect -81356 8648 -81298 9004
rect -81356 7960 -81344 8648
rect -81310 7960 -81298 8648
rect -81356 7604 -81298 7960
rect -79698 8648 -79640 9004
rect -79698 7960 -79686 8648
rect -79652 7960 -79640 8648
rect -79698 7604 -79640 7960
rect -78040 8648 -77982 9004
rect -78040 7960 -78028 8648
rect -77994 7960 -77982 8648
rect -78040 7604 -77982 7960
rect -76382 8648 -76324 9004
rect -76382 7960 -76370 8648
rect -76336 7960 -76324 8648
rect -76382 7604 -76324 7960
rect -74724 8648 -74666 9004
rect -74724 7960 -74712 8648
rect -74678 7960 -74666 8648
rect -74724 7604 -74666 7960
rect -73066 8648 -73008 9004
rect -73066 7960 -73054 8648
rect -73020 7960 -73008 8648
rect -73066 7604 -73008 7960
rect -71408 8648 -71350 9004
rect -71408 7960 -71396 8648
rect -71362 7960 -71350 8648
rect -71408 7604 -71350 7960
rect -69750 8648 -69692 9004
rect -69750 7960 -69738 8648
rect -69704 7960 -69692 8648
rect -69750 7604 -69692 7960
rect -68092 8648 -68034 9004
rect -68092 7960 -68080 8648
rect -68046 7960 -68034 8648
rect -68092 7604 -68034 7960
rect -66434 8648 -66376 9004
rect -66434 7960 -66422 8648
rect -66388 7960 -66376 8648
rect -66434 7604 -66376 7960
rect -64776 8648 -64718 9004
rect -64776 7960 -64764 8648
rect -64730 7960 -64718 8648
rect -64776 7604 -64718 7960
rect -63118 8648 -63060 9004
rect -63118 7960 -63106 8648
rect -63072 7960 -63060 8648
rect -63118 7604 -63060 7960
rect -61460 8648 -61402 9004
rect -61460 7960 -61448 8648
rect -61414 7960 -61402 8648
rect -61460 7604 -61402 7960
rect -59802 8648 -59744 9004
rect -59802 7960 -59790 8648
rect -59756 7960 -59744 8648
rect -59802 7604 -59744 7960
rect -58144 8648 -58086 9004
rect -58144 7960 -58132 8648
rect -58098 7960 -58086 8648
rect -58144 7604 -58086 7960
rect -56486 8648 -56428 9004
rect -56486 7960 -56474 8648
rect -56440 7960 -56428 8648
rect -56486 7604 -56428 7960
rect -54828 8648 -54770 9004
rect -54828 7960 -54816 8648
rect -54782 7960 -54770 8648
rect -54828 7604 -54770 7960
rect -53170 8648 -53112 9004
rect -53170 7960 -53158 8648
rect -53124 7960 -53112 8648
rect -53170 7604 -53112 7960
rect -51512 8648 -51454 9004
rect -51512 7960 -51500 8648
rect -51466 7960 -51454 8648
rect -51512 7604 -51454 7960
rect -49854 8648 -49796 9004
rect -49854 7960 -49842 8648
rect -49808 7960 -49796 8648
rect -49854 7604 -49796 7960
rect -48196 8648 -48138 9004
rect -48196 7960 -48184 8648
rect -48150 7960 -48138 8648
rect -48196 7604 -48138 7960
rect -46538 8648 -46480 9004
rect -46538 7960 -46526 8648
rect -46492 7960 -46480 8648
rect -46538 7604 -46480 7960
rect -44880 8648 -44822 9004
rect -44880 7960 -44868 8648
rect -44834 7960 -44822 8648
rect -44880 7604 -44822 7960
rect -43222 8648 -43164 9004
rect -43222 7960 -43210 8648
rect -43176 7960 -43164 8648
rect -43222 7604 -43164 7960
rect -41564 8648 -41506 9004
rect -41564 7960 -41552 8648
rect -41518 7960 -41506 8648
rect -41564 7604 -41506 7960
rect -39906 8648 -39848 9004
rect -39906 7960 -39894 8648
rect -39860 7960 -39848 8648
rect -39906 7604 -39848 7960
rect -38248 8648 -38190 9004
rect -38248 7960 -38236 8648
rect -38202 7960 -38190 8648
rect -38248 7604 -38190 7960
rect -36590 8648 -36532 9004
rect -36590 7960 -36578 8648
rect -36544 7960 -36532 8648
rect -36590 7604 -36532 7960
rect -34932 8648 -34874 9004
rect -34932 7960 -34920 8648
rect -34886 7960 -34874 8648
rect -34932 7604 -34874 7960
rect -33274 8648 -33216 9004
rect -33274 7960 -33262 8648
rect -33228 7960 -33216 8648
rect -33274 7604 -33216 7960
rect -31616 8648 -31558 9004
rect -31616 7960 -31604 8648
rect -31570 7960 -31558 8648
rect -31616 7604 -31558 7960
rect -29958 8648 -29900 9004
rect -29958 7960 -29946 8648
rect -29912 7960 -29900 8648
rect -29958 7604 -29900 7960
rect -28300 8648 -28242 9004
rect -28300 7960 -28288 8648
rect -28254 7960 -28242 8648
rect -28300 7604 -28242 7960
rect -94620 7012 -94562 7368
rect -94620 6324 -94608 7012
rect -94574 6324 -94562 7012
rect -94620 5968 -94562 6324
rect -92962 7012 -92904 7368
rect -92962 6324 -92950 7012
rect -92916 6324 -92904 7012
rect -92962 5968 -92904 6324
rect -91304 7012 -91246 7368
rect -91304 6324 -91292 7012
rect -91258 6324 -91246 7012
rect -91304 5968 -91246 6324
rect -89646 7012 -89588 7368
rect -89646 6324 -89634 7012
rect -89600 6324 -89588 7012
rect -89646 5968 -89588 6324
rect -87988 7012 -87930 7368
rect -87988 6324 -87976 7012
rect -87942 6324 -87930 7012
rect -87988 5968 -87930 6324
rect -86330 7012 -86272 7368
rect -86330 6324 -86318 7012
rect -86284 6324 -86272 7012
rect -86330 5968 -86272 6324
rect -84672 7012 -84614 7368
rect -84672 6324 -84660 7012
rect -84626 6324 -84614 7012
rect -84672 5968 -84614 6324
rect -83014 7012 -82956 7368
rect -83014 6324 -83002 7012
rect -82968 6324 -82956 7012
rect -83014 5968 -82956 6324
rect -81356 7012 -81298 7368
rect -81356 6324 -81344 7012
rect -81310 6324 -81298 7012
rect -81356 5968 -81298 6324
rect -79698 7012 -79640 7368
rect -79698 6324 -79686 7012
rect -79652 6324 -79640 7012
rect -79698 5968 -79640 6324
rect -78040 7012 -77982 7368
rect -78040 6324 -78028 7012
rect -77994 6324 -77982 7012
rect -78040 5968 -77982 6324
rect -76382 7012 -76324 7368
rect -76382 6324 -76370 7012
rect -76336 6324 -76324 7012
rect -76382 5968 -76324 6324
rect -74724 7012 -74666 7368
rect -74724 6324 -74712 7012
rect -74678 6324 -74666 7012
rect -74724 5968 -74666 6324
rect -73066 7012 -73008 7368
rect -73066 6324 -73054 7012
rect -73020 6324 -73008 7012
rect -73066 5968 -73008 6324
rect -71408 7012 -71350 7368
rect -71408 6324 -71396 7012
rect -71362 6324 -71350 7012
rect -71408 5968 -71350 6324
rect -69750 7012 -69692 7368
rect -69750 6324 -69738 7012
rect -69704 6324 -69692 7012
rect -69750 5968 -69692 6324
rect -68092 7012 -68034 7368
rect -68092 6324 -68080 7012
rect -68046 6324 -68034 7012
rect -68092 5968 -68034 6324
rect -66434 7012 -66376 7368
rect -66434 6324 -66422 7012
rect -66388 6324 -66376 7012
rect -66434 5968 -66376 6324
rect -64776 7012 -64718 7368
rect -64776 6324 -64764 7012
rect -64730 6324 -64718 7012
rect -64776 5968 -64718 6324
rect -63118 7012 -63060 7368
rect -63118 6324 -63106 7012
rect -63072 6324 -63060 7012
rect -63118 5968 -63060 6324
rect -61460 7012 -61402 7368
rect -61460 6324 -61448 7012
rect -61414 6324 -61402 7012
rect -61460 5968 -61402 6324
rect -59802 7012 -59744 7368
rect -59802 6324 -59790 7012
rect -59756 6324 -59744 7012
rect -59802 5968 -59744 6324
rect -58144 7012 -58086 7368
rect -58144 6324 -58132 7012
rect -58098 6324 -58086 7012
rect -58144 5968 -58086 6324
rect -56486 7012 -56428 7368
rect -56486 6324 -56474 7012
rect -56440 6324 -56428 7012
rect -56486 5968 -56428 6324
rect -54828 7012 -54770 7368
rect -54828 6324 -54816 7012
rect -54782 6324 -54770 7012
rect -54828 5968 -54770 6324
rect -53170 7012 -53112 7368
rect -53170 6324 -53158 7012
rect -53124 6324 -53112 7012
rect -53170 5968 -53112 6324
rect -51512 7012 -51454 7368
rect -51512 6324 -51500 7012
rect -51466 6324 -51454 7012
rect -51512 5968 -51454 6324
rect -49854 7012 -49796 7368
rect -49854 6324 -49842 7012
rect -49808 6324 -49796 7012
rect -49854 5968 -49796 6324
rect -48196 7012 -48138 7368
rect -48196 6324 -48184 7012
rect -48150 6324 -48138 7012
rect -48196 5968 -48138 6324
rect -46538 7012 -46480 7368
rect -46538 6324 -46526 7012
rect -46492 6324 -46480 7012
rect -46538 5968 -46480 6324
rect -44880 7012 -44822 7368
rect -44880 6324 -44868 7012
rect -44834 6324 -44822 7012
rect -44880 5968 -44822 6324
rect -43222 7012 -43164 7368
rect -43222 6324 -43210 7012
rect -43176 6324 -43164 7012
rect -43222 5968 -43164 6324
rect -41564 7012 -41506 7368
rect -41564 6324 -41552 7012
rect -41518 6324 -41506 7012
rect -41564 5968 -41506 6324
rect -39906 7012 -39848 7368
rect -39906 6324 -39894 7012
rect -39860 6324 -39848 7012
rect -39906 5968 -39848 6324
rect -38248 7012 -38190 7368
rect -38248 6324 -38236 7012
rect -38202 6324 -38190 7012
rect -38248 5968 -38190 6324
rect -36590 7012 -36532 7368
rect -36590 6324 -36578 7012
rect -36544 6324 -36532 7012
rect -36590 5968 -36532 6324
rect -34932 7012 -34874 7368
rect -34932 6324 -34920 7012
rect -34886 6324 -34874 7012
rect -34932 5968 -34874 6324
rect -33274 7012 -33216 7368
rect -33274 6324 -33262 7012
rect -33228 6324 -33216 7012
rect -33274 5968 -33216 6324
rect -31616 7012 -31558 7368
rect -31616 6324 -31604 7012
rect -31570 6324 -31558 7012
rect -31616 5968 -31558 6324
rect -29958 7012 -29900 7368
rect -29958 6324 -29946 7012
rect -29912 6324 -29900 7012
rect -29958 5968 -29900 6324
rect -28300 7012 -28242 7368
rect -28300 6324 -28288 7012
rect -28254 6324 -28242 7012
rect -28300 5968 -28242 6324
rect -94620 5376 -94562 5732
rect -94620 4688 -94608 5376
rect -94574 4688 -94562 5376
rect -94620 4332 -94562 4688
rect -92962 5376 -92904 5732
rect -92962 4688 -92950 5376
rect -92916 4688 -92904 5376
rect -92962 4332 -92904 4688
rect -91304 5376 -91246 5732
rect -91304 4688 -91292 5376
rect -91258 4688 -91246 5376
rect -91304 4332 -91246 4688
rect -89646 5376 -89588 5732
rect -89646 4688 -89634 5376
rect -89600 4688 -89588 5376
rect -89646 4332 -89588 4688
rect -87988 5376 -87930 5732
rect -87988 4688 -87976 5376
rect -87942 4688 -87930 5376
rect -87988 4332 -87930 4688
rect -86330 5376 -86272 5732
rect -86330 4688 -86318 5376
rect -86284 4688 -86272 5376
rect -86330 4332 -86272 4688
rect -84672 5376 -84614 5732
rect -84672 4688 -84660 5376
rect -84626 4688 -84614 5376
rect -84672 4332 -84614 4688
rect -83014 5376 -82956 5732
rect -83014 4688 -83002 5376
rect -82968 4688 -82956 5376
rect -83014 4332 -82956 4688
rect -81356 5376 -81298 5732
rect -81356 4688 -81344 5376
rect -81310 4688 -81298 5376
rect -81356 4332 -81298 4688
rect -79698 5376 -79640 5732
rect -79698 4688 -79686 5376
rect -79652 4688 -79640 5376
rect -79698 4332 -79640 4688
rect -78040 5376 -77982 5732
rect -78040 4688 -78028 5376
rect -77994 4688 -77982 5376
rect -78040 4332 -77982 4688
rect -76382 5376 -76324 5732
rect -76382 4688 -76370 5376
rect -76336 4688 -76324 5376
rect -76382 4332 -76324 4688
rect -74724 5376 -74666 5732
rect -74724 4688 -74712 5376
rect -74678 4688 -74666 5376
rect -74724 4332 -74666 4688
rect -73066 5376 -73008 5732
rect -73066 4688 -73054 5376
rect -73020 4688 -73008 5376
rect -73066 4332 -73008 4688
rect -71408 5376 -71350 5732
rect -71408 4688 -71396 5376
rect -71362 4688 -71350 5376
rect -71408 4332 -71350 4688
rect -69750 5376 -69692 5732
rect -69750 4688 -69738 5376
rect -69704 4688 -69692 5376
rect -69750 4332 -69692 4688
rect -68092 5376 -68034 5732
rect -68092 4688 -68080 5376
rect -68046 4688 -68034 5376
rect -68092 4332 -68034 4688
rect -66434 5376 -66376 5732
rect -66434 4688 -66422 5376
rect -66388 4688 -66376 5376
rect -66434 4332 -66376 4688
rect -64776 5376 -64718 5732
rect -64776 4688 -64764 5376
rect -64730 4688 -64718 5376
rect -64776 4332 -64718 4688
rect -63118 5376 -63060 5732
rect -63118 4688 -63106 5376
rect -63072 4688 -63060 5376
rect -63118 4332 -63060 4688
rect -61460 5376 -61402 5732
rect -61460 4688 -61448 5376
rect -61414 4688 -61402 5376
rect -61460 4332 -61402 4688
rect -59802 5376 -59744 5732
rect -59802 4688 -59790 5376
rect -59756 4688 -59744 5376
rect -59802 4332 -59744 4688
rect -58144 5376 -58086 5732
rect -58144 4688 -58132 5376
rect -58098 4688 -58086 5376
rect -58144 4332 -58086 4688
rect -56486 5376 -56428 5732
rect -56486 4688 -56474 5376
rect -56440 4688 -56428 5376
rect -56486 4332 -56428 4688
rect -54828 5376 -54770 5732
rect -54828 4688 -54816 5376
rect -54782 4688 -54770 5376
rect -54828 4332 -54770 4688
rect -53170 5376 -53112 5732
rect -53170 4688 -53158 5376
rect -53124 4688 -53112 5376
rect -53170 4332 -53112 4688
rect -51512 5376 -51454 5732
rect -51512 4688 -51500 5376
rect -51466 4688 -51454 5376
rect -51512 4332 -51454 4688
rect -49854 5376 -49796 5732
rect -49854 4688 -49842 5376
rect -49808 4688 -49796 5376
rect -49854 4332 -49796 4688
rect -48196 5376 -48138 5732
rect -48196 4688 -48184 5376
rect -48150 4688 -48138 5376
rect -48196 4332 -48138 4688
rect -46538 5376 -46480 5732
rect -46538 4688 -46526 5376
rect -46492 4688 -46480 5376
rect -46538 4332 -46480 4688
rect -44880 5376 -44822 5732
rect -44880 4688 -44868 5376
rect -44834 4688 -44822 5376
rect -44880 4332 -44822 4688
rect -43222 5376 -43164 5732
rect -43222 4688 -43210 5376
rect -43176 4688 -43164 5376
rect -43222 4332 -43164 4688
rect -41564 5376 -41506 5732
rect -41564 4688 -41552 5376
rect -41518 4688 -41506 5376
rect -41564 4332 -41506 4688
rect -39906 5376 -39848 5732
rect -39906 4688 -39894 5376
rect -39860 4688 -39848 5376
rect -39906 4332 -39848 4688
rect -38248 5376 -38190 5732
rect -38248 4688 -38236 5376
rect -38202 4688 -38190 5376
rect -38248 4332 -38190 4688
rect -36590 5376 -36532 5732
rect -36590 4688 -36578 5376
rect -36544 4688 -36532 5376
rect -36590 4332 -36532 4688
rect -34932 5376 -34874 5732
rect -34932 4688 -34920 5376
rect -34886 4688 -34874 5376
rect -34932 4332 -34874 4688
rect -33274 5376 -33216 5732
rect -33274 4688 -33262 5376
rect -33228 4688 -33216 5376
rect -33274 4332 -33216 4688
rect -31616 5376 -31558 5732
rect -31616 4688 -31604 5376
rect -31570 4688 -31558 5376
rect -31616 4332 -31558 4688
rect -29958 5376 -29900 5732
rect -29958 4688 -29946 5376
rect -29912 4688 -29900 5376
rect -29958 4332 -29900 4688
rect -28300 5376 -28242 5732
rect -28300 4688 -28288 5376
rect -28254 4688 -28242 5376
rect -28300 4332 -28242 4688
rect -61778 3796 -61720 3890
rect -61782 3784 -61720 3796
rect -61782 3596 -61770 3784
rect -61736 3596 -61720 3784
rect -61782 3584 -61720 3596
rect -61778 3490 -61720 3584
rect -61690 3784 -61624 3890
rect -61690 3596 -61674 3784
rect -61640 3596 -61624 3784
rect -61690 3490 -61624 3596
rect -61594 3784 -61528 3890
rect -61594 3596 -61578 3784
rect -61544 3596 -61528 3784
rect -61594 3490 -61528 3596
rect -61498 3784 -61432 3890
rect -61498 3596 -61482 3784
rect -61448 3596 -61432 3784
rect -61498 3490 -61432 3596
rect -61402 3796 -61344 3890
rect 2608 5660 2666 5916
rect 2608 5172 2620 5660
rect 2654 5172 2666 5660
rect 1062 4932 1120 5038
rect 1062 4744 1074 4932
rect 1108 4744 1120 4932
rect 1062 4638 1120 4744
rect 1150 4932 1208 5038
rect 1150 4744 1162 4932
rect 1196 4744 1208 4932
rect 1150 4638 1208 4744
rect 1294 4930 1352 5036
rect 1294 4742 1306 4930
rect 1340 4742 1352 4930
rect 1294 4636 1352 4742
rect 1382 4930 1440 5036
rect 1382 4742 1394 4930
rect 1428 4742 1440 4930
rect 1382 4636 1440 4742
rect 1522 4928 1580 5034
rect 1522 4740 1534 4928
rect 1568 4740 1580 4928
rect 1522 4634 1580 4740
rect 1610 4928 1668 5034
rect 1610 4740 1622 4928
rect 1656 4740 1668 4928
rect 1610 4634 1668 4740
rect 1740 4930 1798 5036
rect 1740 4742 1752 4930
rect 1786 4742 1798 4930
rect 1740 4636 1798 4742
rect 1828 4930 1886 5036
rect 1828 4742 1840 4930
rect 1874 4742 1886 4930
rect 2608 4916 2666 5172
rect 2866 5660 2924 5916
rect 2866 5172 2878 5660
rect 2912 5172 2924 5660
rect 2866 4916 2924 5172
rect 3264 5668 3322 5924
rect 3264 5180 3276 5668
rect 3310 5180 3322 5668
rect 3264 4924 3322 5180
rect 3522 5668 3580 5924
rect 3522 5180 3534 5668
rect 3568 5180 3580 5668
rect 3522 4924 3580 5180
rect 3780 5668 3838 5924
rect 3780 5180 3792 5668
rect 3826 5180 3838 5668
rect 3780 4924 3838 5180
rect 4264 5668 4322 5924
rect 4264 5180 4276 5668
rect 4310 5180 4322 5668
rect 4264 4924 4322 5180
rect 4522 5668 4580 5924
rect 4522 5180 4534 5668
rect 4568 5180 4580 5668
rect 4522 4924 4580 5180
rect 4780 5668 4838 5924
rect 4780 5180 4792 5668
rect 4826 5180 4838 5668
rect 4780 4924 4838 5180
rect 5170 5672 5228 5928
rect 5170 5184 5182 5672
rect 5216 5184 5228 5672
rect 5170 4928 5228 5184
rect 5428 5672 5486 5928
rect 5428 5184 5440 5672
rect 5474 5184 5486 5672
rect 5428 4928 5486 5184
rect 8544 5400 8602 5656
rect 6248 4950 6306 5056
rect 1828 4636 1886 4742
rect 6248 4762 6260 4950
rect 6294 4762 6306 4950
rect 6248 4656 6306 4762
rect 6336 4950 6394 5056
rect 6336 4762 6348 4950
rect 6382 4762 6394 4950
rect 6336 4656 6394 4762
rect 6480 4948 6538 5054
rect 6480 4760 6492 4948
rect 6526 4760 6538 4948
rect 6480 4654 6538 4760
rect 6568 4948 6626 5054
rect 6568 4760 6580 4948
rect 6614 4760 6626 4948
rect 6568 4654 6626 4760
rect 6708 4946 6766 5052
rect 6708 4758 6720 4946
rect 6754 4758 6766 4946
rect 6708 4652 6766 4758
rect 6796 4946 6854 5052
rect 6796 4758 6808 4946
rect 6842 4758 6854 4946
rect 6796 4652 6854 4758
rect 6926 4948 6984 5054
rect 6926 4760 6938 4948
rect 6972 4760 6984 4948
rect 6926 4654 6984 4760
rect 7014 4948 7072 5054
rect 7014 4760 7026 4948
rect 7060 4760 7072 4948
rect 7014 4654 7072 4760
rect 8544 4912 8556 5400
rect 8590 4912 8602 5400
rect 8544 4656 8602 4912
rect 8802 5400 8860 5656
rect 8802 4912 8814 5400
rect 8848 4912 8860 5400
rect 8802 4656 8860 4912
rect 9023 5392 9081 5648
rect 9023 4904 9035 5392
rect 9069 4904 9081 5392
rect 9023 4648 9081 4904
rect 9281 5392 9339 5648
rect 9281 4904 9293 5392
rect 9327 4904 9339 5392
rect 9281 4648 9339 4904
rect 9539 5392 9597 5648
rect 9539 4904 9551 5392
rect 9585 4904 9597 5392
rect 9539 4648 9597 4904
rect 9681 5394 9739 5650
rect 9681 4906 9693 5394
rect 9727 4906 9739 5394
rect 9681 4650 9739 4906
rect 9939 5394 9997 5650
rect 9939 5040 9951 5394
rect 9985 5040 9997 5394
rect 9939 4650 9997 5040
rect 10197 5394 10255 5650
rect 10197 4906 10209 5394
rect 10243 4906 10255 5394
rect 10197 4650 10255 4906
rect 10338 5374 10396 5630
rect 10338 4886 10350 5374
rect 10384 4886 10396 5374
rect 10338 4630 10396 4886
rect 10596 5374 10654 5630
rect 10596 4886 10608 5374
rect 10642 4886 10654 5374
rect 13818 5272 13876 5528
rect 10596 4630 10654 4886
rect 11424 4962 11482 5068
rect 11424 4774 11436 4962
rect 11470 4774 11482 4962
rect 11424 4668 11482 4774
rect 11512 4962 11570 5068
rect 11512 4774 11524 4962
rect 11558 4774 11570 4962
rect 11512 4668 11570 4774
rect 11656 4960 11714 5066
rect 11656 4772 11668 4960
rect 11702 4772 11714 4960
rect 11656 4666 11714 4772
rect 11744 4960 11802 5066
rect 11744 4772 11756 4960
rect 11790 4772 11802 4960
rect 11744 4666 11802 4772
rect 11884 4958 11942 5064
rect 11884 4770 11896 4958
rect 11930 4770 11942 4958
rect 11884 4664 11942 4770
rect 11972 4958 12030 5064
rect 11972 4770 11984 4958
rect 12018 4770 12030 4958
rect 11972 4664 12030 4770
rect 12102 4960 12160 5066
rect 12102 4772 12114 4960
rect 12148 4772 12160 4960
rect 12102 4666 12160 4772
rect 12190 4960 12248 5066
rect 12190 4772 12202 4960
rect 12236 4772 12248 4960
rect 12190 4666 12248 4772
rect 13818 4784 13830 5272
rect 13864 4784 13876 5272
rect 13818 4528 13876 4784
rect 14076 5272 14134 5528
rect 14076 4784 14088 5272
rect 14122 4784 14134 5272
rect 14076 4528 14134 4784
rect 14212 5254 14270 5510
rect 14212 4766 14224 5254
rect 14258 4766 14270 5254
rect 14212 4510 14270 4766
rect 14670 5254 14728 5510
rect 14670 4766 14682 5254
rect 14716 4766 14728 5254
rect 14670 4510 14728 4766
rect 14784 5254 14842 5510
rect 14784 4766 14796 5254
rect 14830 4766 14842 5254
rect 14784 4510 14842 4766
rect 15242 5254 15300 5510
rect 15242 4766 15254 5254
rect 15288 4766 15300 5254
rect 15242 4510 15300 4766
rect 15406 5284 15464 5540
rect 15406 4796 15418 5284
rect 15452 4796 15464 5284
rect 15406 4540 15464 4796
rect 15664 5284 15722 5540
rect 15664 4796 15676 5284
rect 15710 4796 15722 5284
rect 15664 4540 15722 4796
rect 17080 4754 17138 4860
rect 17080 4566 17092 4754
rect 17126 4566 17138 4754
rect 17080 4460 17138 4566
rect 17168 4754 17226 4860
rect 17168 4566 17180 4754
rect 17214 4566 17226 4754
rect 17168 4460 17226 4566
rect 17312 4752 17370 4858
rect 17312 4564 17324 4752
rect 17358 4564 17370 4752
rect 17312 4458 17370 4564
rect 17400 4752 17458 4858
rect 17400 4564 17412 4752
rect 17446 4564 17458 4752
rect 17400 4458 17458 4564
rect 17540 4750 17598 4856
rect 17540 4562 17552 4750
rect 17586 4562 17598 4750
rect 17540 4456 17598 4562
rect 17628 4750 17686 4856
rect 17628 4562 17640 4750
rect 17674 4562 17686 4750
rect 17628 4456 17686 4562
rect 17758 4752 17816 4858
rect 17758 4564 17770 4752
rect 17804 4564 17816 4752
rect 17758 4458 17816 4564
rect 17846 4752 17904 4858
rect 17846 4564 17858 4752
rect 17892 4564 17904 4752
rect 17846 4458 17904 4564
rect -61402 3784 -61340 3796
rect -61402 3596 -61386 3784
rect -61352 3596 -61340 3784
rect -61402 3584 -61340 3596
rect -61402 3490 -61344 3584
rect 27078 2832 27136 2844
rect 26874 2794 26932 2806
rect 26874 2482 26886 2794
rect 26920 2482 26932 2794
rect 26874 2470 26932 2482
rect 26962 2794 27020 2806
rect 26962 2482 26974 2794
rect 27008 2482 27020 2794
rect 27078 2520 27090 2832
rect 27124 2520 27136 2832
rect 27078 2508 27136 2520
rect 27166 2832 27224 2844
rect 27166 2520 27178 2832
rect 27212 2520 27224 2832
rect 27690 2840 27748 2852
rect 27166 2508 27224 2520
rect 27486 2802 27544 2814
rect 26962 2470 27020 2482
rect 27486 2490 27498 2802
rect 27532 2490 27544 2802
rect 27486 2478 27544 2490
rect 27574 2802 27632 2814
rect 27574 2490 27586 2802
rect 27620 2490 27632 2802
rect 27690 2528 27702 2840
rect 27736 2528 27748 2840
rect 27690 2516 27748 2528
rect 27778 2840 27836 2852
rect 27778 2528 27790 2840
rect 27824 2528 27836 2840
rect 28268 2836 28326 2848
rect 27778 2516 27836 2528
rect 28064 2798 28122 2810
rect 27574 2478 27632 2490
rect 28064 2486 28076 2798
rect 28110 2486 28122 2798
rect 28064 2474 28122 2486
rect 28152 2798 28210 2810
rect 28152 2486 28164 2798
rect 28198 2486 28210 2798
rect 28268 2524 28280 2836
rect 28314 2524 28326 2836
rect 28268 2512 28326 2524
rect 28356 2836 28414 2848
rect 28356 2524 28368 2836
rect 28402 2524 28414 2836
rect 28842 2844 28900 2856
rect 28356 2512 28414 2524
rect 28638 2806 28696 2818
rect 28152 2474 28210 2486
rect 28638 2494 28650 2806
rect 28684 2494 28696 2806
rect 28638 2482 28696 2494
rect 28726 2806 28784 2818
rect 28726 2494 28738 2806
rect 28772 2494 28784 2806
rect 28842 2532 28854 2844
rect 28888 2532 28900 2844
rect 28842 2520 28900 2532
rect 28930 2844 28988 2856
rect 28930 2532 28942 2844
rect 28976 2532 28988 2844
rect 29420 2844 29478 2856
rect 28930 2520 28988 2532
rect 29216 2806 29274 2818
rect 28726 2482 28784 2494
rect 29216 2494 29228 2806
rect 29262 2494 29274 2806
rect 29216 2482 29274 2494
rect 29304 2806 29362 2818
rect 29304 2494 29316 2806
rect 29350 2494 29362 2806
rect 29420 2532 29432 2844
rect 29466 2532 29478 2844
rect 29420 2520 29478 2532
rect 29508 2844 29566 2856
rect 29508 2532 29520 2844
rect 29554 2532 29566 2844
rect 29998 2844 30056 2856
rect 29508 2520 29566 2532
rect 29794 2806 29852 2818
rect 29304 2482 29362 2494
rect 29794 2494 29806 2806
rect 29840 2494 29852 2806
rect 29794 2482 29852 2494
rect 29882 2806 29940 2818
rect 29882 2494 29894 2806
rect 29928 2494 29940 2806
rect 29998 2532 30010 2844
rect 30044 2532 30056 2844
rect 29998 2520 30056 2532
rect 30086 2844 30144 2856
rect 30086 2532 30098 2844
rect 30132 2532 30144 2844
rect 30580 2848 30638 2860
rect 30086 2520 30144 2532
rect 30376 2810 30434 2822
rect 29882 2482 29940 2494
rect 30376 2498 30388 2810
rect 30422 2498 30434 2810
rect 30376 2486 30434 2498
rect 30464 2810 30522 2822
rect 30464 2498 30476 2810
rect 30510 2498 30522 2810
rect 30580 2536 30592 2848
rect 30626 2536 30638 2848
rect 30580 2524 30638 2536
rect 30668 2848 30726 2860
rect 30668 2536 30680 2848
rect 30714 2536 30726 2848
rect 31156 2844 31214 2856
rect 30668 2524 30726 2536
rect 30952 2806 31010 2818
rect 30464 2486 30522 2498
rect 30952 2494 30964 2806
rect 30998 2494 31010 2806
rect 30952 2482 31010 2494
rect 31040 2806 31098 2818
rect 31040 2494 31052 2806
rect 31086 2494 31098 2806
rect 31156 2532 31168 2844
rect 31202 2532 31214 2844
rect 31156 2520 31214 2532
rect 31244 2844 31302 2856
rect 31244 2532 31256 2844
rect 31290 2532 31302 2844
rect 31726 2840 31784 2852
rect 31244 2520 31302 2532
rect 31522 2802 31580 2814
rect 31040 2482 31098 2494
rect 31522 2490 31534 2802
rect 31568 2490 31580 2802
rect 31522 2478 31580 2490
rect 31610 2802 31668 2814
rect 31610 2490 31622 2802
rect 31656 2490 31668 2802
rect 31726 2528 31738 2840
rect 31772 2528 31784 2840
rect 31726 2516 31784 2528
rect 31814 2840 31872 2852
rect 31814 2528 31826 2840
rect 31860 2528 31872 2840
rect 31814 2516 31872 2528
rect 31610 2478 31668 2490
rect 28468 778 28526 790
rect 28268 740 28326 752
rect 28268 428 28280 740
rect 28314 428 28326 740
rect 28268 416 28326 428
rect 28356 740 28414 752
rect 28356 428 28368 740
rect 28402 428 28414 740
rect 28468 466 28480 778
rect 28514 466 28526 778
rect 28468 454 28526 466
rect 28556 778 28614 790
rect 28556 466 28568 778
rect 28602 466 28614 778
rect 28556 454 28614 466
rect 28670 738 28728 750
rect 28356 416 28414 428
rect 28670 426 28682 738
rect 28716 426 28728 738
rect 28670 414 28728 426
rect 28758 738 28816 750
rect 28758 426 28770 738
rect 28804 426 28816 738
rect 28758 414 28816 426
rect 28468 272 28526 284
rect 28268 234 28326 246
rect 28268 -78 28280 234
rect 28314 -78 28326 234
rect 28268 -90 28326 -78
rect 28356 234 28414 246
rect 28356 -78 28368 234
rect 28402 -78 28414 234
rect 28468 -40 28480 272
rect 28514 -40 28526 272
rect 28468 -52 28526 -40
rect 28556 272 28614 284
rect 28556 -40 28568 272
rect 28602 -40 28614 272
rect 28556 -52 28614 -40
rect 28668 234 28726 246
rect 28356 -90 28414 -78
rect 28668 -78 28680 234
rect 28714 -78 28726 234
rect 28668 -90 28726 -78
rect 28756 234 28814 246
rect 28756 -78 28768 234
rect 28802 -78 28814 234
rect 28756 -90 28814 -78
rect 28468 -236 28526 -224
rect 28268 -274 28326 -262
rect 28268 -586 28280 -274
rect 28314 -586 28326 -274
rect 28268 -598 28326 -586
rect 28356 -274 28414 -262
rect 28356 -586 28368 -274
rect 28402 -586 28414 -274
rect 28468 -548 28480 -236
rect 28514 -548 28526 -236
rect 28468 -560 28526 -548
rect 28556 -236 28614 -224
rect 28556 -548 28568 -236
rect 28602 -548 28614 -236
rect 28556 -560 28614 -548
rect 28668 -274 28726 -262
rect 28356 -598 28414 -586
rect 28668 -586 28680 -274
rect 28714 -586 28726 -274
rect 28668 -598 28726 -586
rect 28756 -274 28814 -262
rect 28756 -586 28768 -274
rect 28802 -586 28814 -274
rect 28756 -598 28814 -586
rect 8761 -1042 8813 -1028
rect 8761 -1076 8769 -1042
rect 8803 -1076 8813 -1042
rect 8761 -1110 8813 -1076
rect 8761 -1144 8769 -1110
rect 8803 -1144 8813 -1110
rect 8761 -1156 8813 -1144
rect 8843 -1058 8897 -1028
rect 8843 -1092 8853 -1058
rect 8887 -1092 8897 -1058
rect 8843 -1156 8897 -1092
rect 8927 -1042 8979 -1028
rect 8927 -1076 8937 -1042
rect 8971 -1076 8979 -1042
rect 8927 -1110 8979 -1076
rect 9112 -1034 9164 -1022
rect 9112 -1068 9120 -1034
rect 9154 -1068 9164 -1034
rect 9112 -1106 9164 -1068
rect 9194 -1042 9256 -1022
rect 9194 -1076 9204 -1042
rect 9238 -1076 9256 -1042
rect 9194 -1106 9256 -1076
rect 9286 -1036 9355 -1022
rect 9286 -1070 9297 -1036
rect 9331 -1070 9355 -1036
rect 9286 -1106 9355 -1070
rect 9385 -1060 9495 -1022
rect 9385 -1094 9451 -1060
rect 9485 -1094 9495 -1060
rect 9385 -1106 9495 -1094
rect 9525 -1044 9592 -1022
rect 9525 -1078 9548 -1044
rect 9582 -1078 9592 -1044
rect 9525 -1106 9592 -1078
rect 9622 -1060 9674 -1022
rect 9622 -1094 9632 -1060
rect 9666 -1094 9674 -1060
rect 9622 -1106 9674 -1094
rect 9737 -1034 9789 -1022
rect 9737 -1068 9745 -1034
rect 9779 -1068 9789 -1034
rect 8927 -1144 8937 -1110
rect 8971 -1144 8979 -1110
rect 8927 -1156 8979 -1144
rect 9737 -1190 9789 -1068
rect 9819 -1042 9888 -1022
rect 9819 -1076 9833 -1042
rect 9867 -1076 9888 -1042
rect 9819 -1106 9888 -1076
rect 9918 -1035 9974 -1022
rect 9918 -1069 9930 -1035
rect 9964 -1069 9974 -1035
rect 9918 -1106 9974 -1069
rect 10004 -1106 10058 -1022
rect 10088 -1034 10166 -1022
rect 10088 -1068 10122 -1034
rect 10156 -1068 10166 -1034
rect 10088 -1106 10166 -1068
rect 10196 -1060 10250 -1022
rect 10196 -1094 10206 -1060
rect 10240 -1094 10250 -1060
rect 10196 -1106 10250 -1094
rect 10280 -1034 10414 -1022
rect 10280 -1068 10292 -1034
rect 10326 -1068 10370 -1034
rect 10404 -1068 10414 -1034
rect 10280 -1106 10414 -1068
rect 9819 -1190 9873 -1106
rect 10364 -1222 10414 -1106
rect 10444 -1042 10500 -1022
rect 10444 -1076 10454 -1042
rect 10488 -1076 10500 -1042
rect 10444 -1110 10500 -1076
rect 10444 -1144 10454 -1110
rect 10488 -1144 10500 -1110
rect 10444 -1178 10500 -1144
rect 10581 -1034 10633 -1022
rect 10581 -1068 10589 -1034
rect 10623 -1068 10633 -1034
rect 10581 -1102 10633 -1068
rect 10581 -1136 10589 -1102
rect 10623 -1136 10633 -1102
rect 10581 -1150 10633 -1136
rect 10663 -1034 10730 -1022
rect 10663 -1068 10686 -1034
rect 10720 -1068 10730 -1034
rect 10663 -1102 10730 -1068
rect 10663 -1136 10686 -1102
rect 10720 -1136 10730 -1102
rect 10663 -1150 10730 -1136
rect 10444 -1212 10454 -1178
rect 10488 -1212 10500 -1178
rect 10444 -1222 10500 -1212
rect 10678 -1170 10730 -1150
rect 10678 -1204 10686 -1170
rect 10720 -1204 10730 -1170
rect 10678 -1222 10730 -1204
rect 10760 -1070 10812 -1022
rect 10760 -1104 10770 -1070
rect 10804 -1104 10812 -1070
rect 10760 -1138 10812 -1104
rect 10760 -1172 10770 -1138
rect 10804 -1172 10812 -1138
rect 11227 -1042 11279 -1028
rect 11227 -1076 11235 -1042
rect 11269 -1076 11279 -1042
rect 11227 -1110 11279 -1076
rect 11227 -1144 11235 -1110
rect 11269 -1144 11279 -1110
rect 11227 -1156 11279 -1144
rect 11309 -1058 11363 -1028
rect 11309 -1092 11319 -1058
rect 11353 -1092 11363 -1058
rect 11309 -1156 11363 -1092
rect 11393 -1042 11445 -1028
rect 11393 -1076 11403 -1042
rect 11437 -1076 11445 -1042
rect 11393 -1110 11445 -1076
rect 11578 -1034 11630 -1022
rect 11578 -1068 11586 -1034
rect 11620 -1068 11630 -1034
rect 11578 -1106 11630 -1068
rect 11660 -1042 11722 -1022
rect 11660 -1076 11670 -1042
rect 11704 -1076 11722 -1042
rect 11660 -1106 11722 -1076
rect 11752 -1036 11821 -1022
rect 11752 -1070 11763 -1036
rect 11797 -1070 11821 -1036
rect 11752 -1106 11821 -1070
rect 11851 -1060 11961 -1022
rect 11851 -1094 11917 -1060
rect 11951 -1094 11961 -1060
rect 11851 -1106 11961 -1094
rect 11991 -1044 12058 -1022
rect 11991 -1078 12014 -1044
rect 12048 -1078 12058 -1044
rect 11991 -1106 12058 -1078
rect 12088 -1060 12140 -1022
rect 12088 -1094 12098 -1060
rect 12132 -1094 12140 -1060
rect 12088 -1106 12140 -1094
rect 12203 -1034 12255 -1022
rect 12203 -1068 12211 -1034
rect 12245 -1068 12255 -1034
rect 11393 -1144 11403 -1110
rect 11437 -1144 11445 -1110
rect 11393 -1156 11445 -1144
rect 10760 -1222 10812 -1172
rect 12203 -1190 12255 -1068
rect 12285 -1042 12354 -1022
rect 12285 -1076 12299 -1042
rect 12333 -1076 12354 -1042
rect 12285 -1106 12354 -1076
rect 12384 -1035 12440 -1022
rect 12384 -1069 12396 -1035
rect 12430 -1069 12440 -1035
rect 12384 -1106 12440 -1069
rect 12470 -1106 12524 -1022
rect 12554 -1034 12632 -1022
rect 12554 -1068 12588 -1034
rect 12622 -1068 12632 -1034
rect 12554 -1106 12632 -1068
rect 12662 -1060 12716 -1022
rect 12662 -1094 12672 -1060
rect 12706 -1094 12716 -1060
rect 12662 -1106 12716 -1094
rect 12746 -1034 12880 -1022
rect 12746 -1068 12758 -1034
rect 12792 -1068 12836 -1034
rect 12870 -1068 12880 -1034
rect 12746 -1106 12880 -1068
rect 12285 -1190 12339 -1106
rect 12830 -1222 12880 -1106
rect 12910 -1042 12966 -1022
rect 12910 -1076 12920 -1042
rect 12954 -1076 12966 -1042
rect 12910 -1110 12966 -1076
rect 12910 -1144 12920 -1110
rect 12954 -1144 12966 -1110
rect 12910 -1178 12966 -1144
rect 13047 -1034 13099 -1022
rect 13047 -1068 13055 -1034
rect 13089 -1068 13099 -1034
rect 13047 -1102 13099 -1068
rect 13047 -1136 13055 -1102
rect 13089 -1136 13099 -1102
rect 13047 -1150 13099 -1136
rect 13129 -1034 13196 -1022
rect 13129 -1068 13152 -1034
rect 13186 -1068 13196 -1034
rect 13129 -1102 13196 -1068
rect 13129 -1136 13152 -1102
rect 13186 -1136 13196 -1102
rect 13129 -1150 13196 -1136
rect 12910 -1212 12920 -1178
rect 12954 -1212 12966 -1178
rect 12910 -1222 12966 -1212
rect 13144 -1170 13196 -1150
rect 13144 -1204 13152 -1170
rect 13186 -1204 13196 -1170
rect 13144 -1222 13196 -1204
rect 13226 -1070 13278 -1022
rect 13226 -1104 13236 -1070
rect 13270 -1104 13278 -1070
rect 13226 -1138 13278 -1104
rect 13226 -1172 13236 -1138
rect 13270 -1172 13278 -1138
rect 13226 -1222 13278 -1172
rect 10181 -1836 10233 -1824
rect 10181 -1870 10189 -1836
rect 10223 -1870 10233 -1836
rect 10181 -1904 10233 -1870
rect 10181 -1938 10189 -1904
rect 10223 -1938 10233 -1904
rect 10181 -1972 10233 -1938
rect 10181 -2006 10189 -1972
rect 10223 -2006 10233 -1972
rect 10181 -2024 10233 -2006
rect 10263 -1836 10317 -1824
rect 10263 -1870 10273 -1836
rect 10307 -1870 10317 -1836
rect 10263 -1904 10317 -1870
rect 10263 -1938 10273 -1904
rect 10307 -1938 10317 -1904
rect 10263 -1972 10317 -1938
rect 10263 -2006 10273 -1972
rect 10307 -2006 10317 -1972
rect 10263 -2024 10317 -2006
rect 10347 -1836 10399 -1824
rect 10347 -1870 10357 -1836
rect 10391 -1870 10399 -1836
rect 10347 -1904 10399 -1870
rect 10347 -1938 10357 -1904
rect 10391 -1938 10399 -1904
rect 10347 -1972 10399 -1938
rect 11227 -1844 11279 -1830
rect 11227 -1878 11235 -1844
rect 11269 -1878 11279 -1844
rect 11227 -1912 11279 -1878
rect 11227 -1946 11235 -1912
rect 11269 -1946 11279 -1912
rect 11227 -1958 11279 -1946
rect 11309 -1860 11363 -1830
rect 11309 -1894 11319 -1860
rect 11353 -1894 11363 -1860
rect 11309 -1958 11363 -1894
rect 11393 -1844 11445 -1830
rect 11393 -1878 11403 -1844
rect 11437 -1878 11445 -1844
rect 11393 -1912 11445 -1878
rect 11578 -1836 11630 -1824
rect 11578 -1870 11586 -1836
rect 11620 -1870 11630 -1836
rect 11578 -1908 11630 -1870
rect 11660 -1844 11722 -1824
rect 11660 -1878 11670 -1844
rect 11704 -1878 11722 -1844
rect 11660 -1908 11722 -1878
rect 11752 -1838 11821 -1824
rect 11752 -1872 11763 -1838
rect 11797 -1872 11821 -1838
rect 11752 -1908 11821 -1872
rect 11851 -1862 11961 -1824
rect 11851 -1896 11917 -1862
rect 11951 -1896 11961 -1862
rect 11851 -1908 11961 -1896
rect 11991 -1846 12058 -1824
rect 11991 -1880 12014 -1846
rect 12048 -1880 12058 -1846
rect 11991 -1908 12058 -1880
rect 12088 -1862 12140 -1824
rect 12088 -1896 12098 -1862
rect 12132 -1896 12140 -1862
rect 12088 -1908 12140 -1896
rect 12203 -1836 12255 -1824
rect 12203 -1870 12211 -1836
rect 12245 -1870 12255 -1836
rect 11393 -1946 11403 -1912
rect 11437 -1946 11445 -1912
rect 11393 -1958 11445 -1946
rect 10347 -2006 10357 -1972
rect 10391 -2006 10399 -1972
rect 10347 -2024 10399 -2006
rect 12203 -1992 12255 -1870
rect 12285 -1844 12354 -1824
rect 12285 -1878 12299 -1844
rect 12333 -1878 12354 -1844
rect 12285 -1908 12354 -1878
rect 12384 -1837 12440 -1824
rect 12384 -1871 12396 -1837
rect 12430 -1871 12440 -1837
rect 12384 -1908 12440 -1871
rect 12470 -1908 12524 -1824
rect 12554 -1836 12632 -1824
rect 12554 -1870 12588 -1836
rect 12622 -1870 12632 -1836
rect 12554 -1908 12632 -1870
rect 12662 -1862 12716 -1824
rect 12662 -1896 12672 -1862
rect 12706 -1896 12716 -1862
rect 12662 -1908 12716 -1896
rect 12746 -1836 12880 -1824
rect 12746 -1870 12758 -1836
rect 12792 -1870 12836 -1836
rect 12870 -1870 12880 -1836
rect 12746 -1908 12880 -1870
rect 12285 -1992 12339 -1908
rect 12830 -2024 12880 -1908
rect 12910 -1844 12966 -1824
rect 12910 -1878 12920 -1844
rect 12954 -1878 12966 -1844
rect 12910 -1912 12966 -1878
rect 12910 -1946 12920 -1912
rect 12954 -1946 12966 -1912
rect 12910 -1980 12966 -1946
rect 13047 -1836 13099 -1824
rect 13047 -1870 13055 -1836
rect 13089 -1870 13099 -1836
rect 13047 -1904 13099 -1870
rect 13047 -1938 13055 -1904
rect 13089 -1938 13099 -1904
rect 13047 -1952 13099 -1938
rect 13129 -1836 13196 -1824
rect 13129 -1870 13152 -1836
rect 13186 -1870 13196 -1836
rect 13129 -1904 13196 -1870
rect 13129 -1938 13152 -1904
rect 13186 -1938 13196 -1904
rect 13129 -1952 13196 -1938
rect 12910 -2014 12920 -1980
rect 12954 -2014 12966 -1980
rect 12910 -2024 12966 -2014
rect 13144 -1972 13196 -1952
rect 13144 -2006 13152 -1972
rect 13186 -2006 13196 -1972
rect 13144 -2024 13196 -2006
rect 13226 -1872 13278 -1824
rect 13226 -1906 13236 -1872
rect 13270 -1906 13278 -1872
rect 13226 -1940 13278 -1906
rect 13226 -1974 13236 -1940
rect 13270 -1974 13278 -1940
rect 13226 -2024 13278 -1974
rect -9131 -4312 -9079 -4298
rect -9131 -4346 -9123 -4312
rect -9089 -4346 -9079 -4312
rect -9131 -4380 -9079 -4346
rect -9131 -4414 -9123 -4380
rect -9089 -4414 -9079 -4380
rect -9131 -4426 -9079 -4414
rect -9049 -4328 -8995 -4298
rect -9049 -4362 -9039 -4328
rect -9005 -4362 -8995 -4328
rect -9049 -4426 -8995 -4362
rect -8965 -4312 -8913 -4298
rect -8965 -4346 -8955 -4312
rect -8921 -4346 -8913 -4312
rect -8965 -4380 -8913 -4346
rect -8780 -4304 -8728 -4292
rect -8780 -4338 -8772 -4304
rect -8738 -4338 -8728 -4304
rect -8780 -4376 -8728 -4338
rect -8698 -4312 -8636 -4292
rect -8698 -4346 -8688 -4312
rect -8654 -4346 -8636 -4312
rect -8698 -4376 -8636 -4346
rect -8606 -4306 -8537 -4292
rect -8606 -4340 -8595 -4306
rect -8561 -4340 -8537 -4306
rect -8606 -4376 -8537 -4340
rect -8507 -4330 -8397 -4292
rect -8507 -4364 -8441 -4330
rect -8407 -4364 -8397 -4330
rect -8507 -4376 -8397 -4364
rect -8367 -4314 -8300 -4292
rect -8367 -4348 -8344 -4314
rect -8310 -4348 -8300 -4314
rect -8367 -4376 -8300 -4348
rect -8270 -4330 -8218 -4292
rect -8270 -4364 -8260 -4330
rect -8226 -4364 -8218 -4330
rect -8270 -4376 -8218 -4364
rect -8155 -4304 -8103 -4292
rect -8155 -4338 -8147 -4304
rect -8113 -4338 -8103 -4304
rect -8965 -4414 -8955 -4380
rect -8921 -4414 -8913 -4380
rect -8965 -4426 -8913 -4414
rect -8155 -4460 -8103 -4338
rect -8073 -4312 -8004 -4292
rect -8073 -4346 -8059 -4312
rect -8025 -4346 -8004 -4312
rect -8073 -4376 -8004 -4346
rect -7974 -4305 -7918 -4292
rect -7974 -4339 -7962 -4305
rect -7928 -4339 -7918 -4305
rect -7974 -4376 -7918 -4339
rect -7888 -4376 -7834 -4292
rect -7804 -4304 -7726 -4292
rect -7804 -4338 -7770 -4304
rect -7736 -4338 -7726 -4304
rect -7804 -4376 -7726 -4338
rect -7696 -4330 -7642 -4292
rect -7696 -4364 -7686 -4330
rect -7652 -4364 -7642 -4330
rect -7696 -4376 -7642 -4364
rect -7612 -4304 -7478 -4292
rect -7612 -4338 -7600 -4304
rect -7566 -4338 -7522 -4304
rect -7488 -4338 -7478 -4304
rect -7612 -4376 -7478 -4338
rect -8073 -4460 -8019 -4376
rect -7528 -4492 -7478 -4376
rect -7448 -4312 -7392 -4292
rect -7448 -4346 -7438 -4312
rect -7404 -4346 -7392 -4312
rect -7448 -4380 -7392 -4346
rect -7448 -4414 -7438 -4380
rect -7404 -4414 -7392 -4380
rect -7448 -4448 -7392 -4414
rect -7311 -4304 -7259 -4292
rect -7311 -4338 -7303 -4304
rect -7269 -4338 -7259 -4304
rect -7311 -4372 -7259 -4338
rect -7311 -4406 -7303 -4372
rect -7269 -4406 -7259 -4372
rect -7311 -4420 -7259 -4406
rect -7229 -4304 -7162 -4292
rect -7229 -4338 -7206 -4304
rect -7172 -4338 -7162 -4304
rect -7229 -4372 -7162 -4338
rect -7229 -4406 -7206 -4372
rect -7172 -4406 -7162 -4372
rect -7229 -4420 -7162 -4406
rect -7448 -4482 -7438 -4448
rect -7404 -4482 -7392 -4448
rect -7448 -4492 -7392 -4482
rect -7214 -4440 -7162 -4420
rect -7214 -4474 -7206 -4440
rect -7172 -4474 -7162 -4440
rect -7214 -4492 -7162 -4474
rect -7132 -4340 -7080 -4292
rect -7132 -4374 -7122 -4340
rect -7088 -4374 -7080 -4340
rect -7132 -4408 -7080 -4374
rect -7132 -4442 -7122 -4408
rect -7088 -4442 -7080 -4408
rect -7015 -4312 -6963 -4298
rect -7015 -4346 -7007 -4312
rect -6973 -4346 -6963 -4312
rect -7015 -4380 -6963 -4346
rect -7015 -4414 -7007 -4380
rect -6973 -4414 -6963 -4380
rect -7015 -4426 -6963 -4414
rect -6933 -4328 -6879 -4298
rect -6933 -4362 -6923 -4328
rect -6889 -4362 -6879 -4328
rect -6933 -4426 -6879 -4362
rect -6849 -4312 -6797 -4298
rect -6849 -4346 -6839 -4312
rect -6805 -4346 -6797 -4312
rect -6849 -4380 -6797 -4346
rect -6664 -4304 -6612 -4292
rect -6664 -4338 -6656 -4304
rect -6622 -4338 -6612 -4304
rect -6664 -4376 -6612 -4338
rect -6582 -4312 -6520 -4292
rect -6582 -4346 -6572 -4312
rect -6538 -4346 -6520 -4312
rect -6582 -4376 -6520 -4346
rect -6490 -4306 -6421 -4292
rect -6490 -4340 -6479 -4306
rect -6445 -4340 -6421 -4306
rect -6490 -4376 -6421 -4340
rect -6391 -4330 -6281 -4292
rect -6391 -4364 -6325 -4330
rect -6291 -4364 -6281 -4330
rect -6391 -4376 -6281 -4364
rect -6251 -4314 -6184 -4292
rect -6251 -4348 -6228 -4314
rect -6194 -4348 -6184 -4314
rect -6251 -4376 -6184 -4348
rect -6154 -4330 -6102 -4292
rect -6154 -4364 -6144 -4330
rect -6110 -4364 -6102 -4330
rect -6154 -4376 -6102 -4364
rect -6039 -4304 -5987 -4292
rect -6039 -4338 -6031 -4304
rect -5997 -4338 -5987 -4304
rect -6849 -4414 -6839 -4380
rect -6805 -4414 -6797 -4380
rect -6849 -4426 -6797 -4414
rect -7132 -4492 -7080 -4442
rect -6039 -4460 -5987 -4338
rect -5957 -4312 -5888 -4292
rect -5957 -4346 -5943 -4312
rect -5909 -4346 -5888 -4312
rect -5957 -4376 -5888 -4346
rect -5858 -4305 -5802 -4292
rect -5858 -4339 -5846 -4305
rect -5812 -4339 -5802 -4305
rect -5858 -4376 -5802 -4339
rect -5772 -4376 -5718 -4292
rect -5688 -4304 -5610 -4292
rect -5688 -4338 -5654 -4304
rect -5620 -4338 -5610 -4304
rect -5688 -4376 -5610 -4338
rect -5580 -4330 -5526 -4292
rect -5580 -4364 -5570 -4330
rect -5536 -4364 -5526 -4330
rect -5580 -4376 -5526 -4364
rect -5496 -4304 -5362 -4292
rect -5496 -4338 -5484 -4304
rect -5450 -4338 -5406 -4304
rect -5372 -4338 -5362 -4304
rect -5496 -4376 -5362 -4338
rect -5957 -4460 -5903 -4376
rect -5412 -4492 -5362 -4376
rect -5332 -4312 -5276 -4292
rect -5332 -4346 -5322 -4312
rect -5288 -4346 -5276 -4312
rect -5332 -4380 -5276 -4346
rect -5332 -4414 -5322 -4380
rect -5288 -4414 -5276 -4380
rect -5332 -4448 -5276 -4414
rect -5195 -4304 -5143 -4292
rect -5195 -4338 -5187 -4304
rect -5153 -4338 -5143 -4304
rect -5195 -4372 -5143 -4338
rect -5195 -4406 -5187 -4372
rect -5153 -4406 -5143 -4372
rect -5195 -4420 -5143 -4406
rect -5113 -4304 -5046 -4292
rect -5113 -4338 -5090 -4304
rect -5056 -4338 -5046 -4304
rect -5113 -4372 -5046 -4338
rect -5113 -4406 -5090 -4372
rect -5056 -4406 -5046 -4372
rect -5113 -4420 -5046 -4406
rect -5332 -4482 -5322 -4448
rect -5288 -4482 -5276 -4448
rect -5332 -4492 -5276 -4482
rect -5098 -4440 -5046 -4420
rect -5098 -4474 -5090 -4440
rect -5056 -4474 -5046 -4440
rect -5098 -4492 -5046 -4474
rect -5016 -4340 -4964 -4292
rect -5016 -4374 -5006 -4340
rect -4972 -4374 -4964 -4340
rect -5016 -4408 -4964 -4374
rect -5016 -4442 -5006 -4408
rect -4972 -4442 -4964 -4408
rect -4899 -4312 -4847 -4298
rect -4899 -4346 -4891 -4312
rect -4857 -4346 -4847 -4312
rect -4899 -4380 -4847 -4346
rect -4899 -4414 -4891 -4380
rect -4857 -4414 -4847 -4380
rect -4899 -4426 -4847 -4414
rect -4817 -4328 -4763 -4298
rect -4817 -4362 -4807 -4328
rect -4773 -4362 -4763 -4328
rect -4817 -4426 -4763 -4362
rect -4733 -4312 -4681 -4298
rect -4733 -4346 -4723 -4312
rect -4689 -4346 -4681 -4312
rect -4733 -4380 -4681 -4346
rect -4548 -4304 -4496 -4292
rect -4548 -4338 -4540 -4304
rect -4506 -4338 -4496 -4304
rect -4548 -4376 -4496 -4338
rect -4466 -4312 -4404 -4292
rect -4466 -4346 -4456 -4312
rect -4422 -4346 -4404 -4312
rect -4466 -4376 -4404 -4346
rect -4374 -4306 -4305 -4292
rect -4374 -4340 -4363 -4306
rect -4329 -4340 -4305 -4306
rect -4374 -4376 -4305 -4340
rect -4275 -4330 -4165 -4292
rect -4275 -4364 -4209 -4330
rect -4175 -4364 -4165 -4330
rect -4275 -4376 -4165 -4364
rect -4135 -4314 -4068 -4292
rect -4135 -4348 -4112 -4314
rect -4078 -4348 -4068 -4314
rect -4135 -4376 -4068 -4348
rect -4038 -4330 -3986 -4292
rect -4038 -4364 -4028 -4330
rect -3994 -4364 -3986 -4330
rect -4038 -4376 -3986 -4364
rect -3923 -4304 -3871 -4292
rect -3923 -4338 -3915 -4304
rect -3881 -4338 -3871 -4304
rect -4733 -4414 -4723 -4380
rect -4689 -4414 -4681 -4380
rect -4733 -4426 -4681 -4414
rect -5016 -4492 -4964 -4442
rect -3923 -4460 -3871 -4338
rect -3841 -4312 -3772 -4292
rect -3841 -4346 -3827 -4312
rect -3793 -4346 -3772 -4312
rect -3841 -4376 -3772 -4346
rect -3742 -4305 -3686 -4292
rect -3742 -4339 -3730 -4305
rect -3696 -4339 -3686 -4305
rect -3742 -4376 -3686 -4339
rect -3656 -4376 -3602 -4292
rect -3572 -4304 -3494 -4292
rect -3572 -4338 -3538 -4304
rect -3504 -4338 -3494 -4304
rect -3572 -4376 -3494 -4338
rect -3464 -4330 -3410 -4292
rect -3464 -4364 -3454 -4330
rect -3420 -4364 -3410 -4330
rect -3464 -4376 -3410 -4364
rect -3380 -4304 -3246 -4292
rect -3380 -4338 -3368 -4304
rect -3334 -4338 -3290 -4304
rect -3256 -4338 -3246 -4304
rect -3380 -4376 -3246 -4338
rect -3841 -4460 -3787 -4376
rect -3296 -4492 -3246 -4376
rect -3216 -4312 -3160 -4292
rect -3216 -4346 -3206 -4312
rect -3172 -4346 -3160 -4312
rect -3216 -4380 -3160 -4346
rect -3216 -4414 -3206 -4380
rect -3172 -4414 -3160 -4380
rect -3216 -4448 -3160 -4414
rect -3079 -4304 -3027 -4292
rect -3079 -4338 -3071 -4304
rect -3037 -4338 -3027 -4304
rect -3079 -4372 -3027 -4338
rect -3079 -4406 -3071 -4372
rect -3037 -4406 -3027 -4372
rect -3079 -4420 -3027 -4406
rect -2997 -4304 -2930 -4292
rect -2997 -4338 -2974 -4304
rect -2940 -4338 -2930 -4304
rect -2997 -4372 -2930 -4338
rect -2997 -4406 -2974 -4372
rect -2940 -4406 -2930 -4372
rect -2997 -4420 -2930 -4406
rect -3216 -4482 -3206 -4448
rect -3172 -4482 -3160 -4448
rect -3216 -4492 -3160 -4482
rect -2982 -4440 -2930 -4420
rect -2982 -4474 -2974 -4440
rect -2940 -4474 -2930 -4440
rect -2982 -4492 -2930 -4474
rect -2900 -4340 -2848 -4292
rect -2900 -4374 -2890 -4340
rect -2856 -4374 -2848 -4340
rect -2900 -4408 -2848 -4374
rect -2900 -4442 -2890 -4408
rect -2856 -4442 -2848 -4408
rect -2783 -4312 -2731 -4298
rect -2783 -4346 -2775 -4312
rect -2741 -4346 -2731 -4312
rect -2783 -4380 -2731 -4346
rect -2783 -4414 -2775 -4380
rect -2741 -4414 -2731 -4380
rect -2783 -4426 -2731 -4414
rect -2701 -4328 -2647 -4298
rect -2701 -4362 -2691 -4328
rect -2657 -4362 -2647 -4328
rect -2701 -4426 -2647 -4362
rect -2617 -4312 -2565 -4298
rect -2617 -4346 -2607 -4312
rect -2573 -4346 -2565 -4312
rect -2617 -4380 -2565 -4346
rect -2432 -4304 -2380 -4292
rect -2432 -4338 -2424 -4304
rect -2390 -4338 -2380 -4304
rect -2432 -4376 -2380 -4338
rect -2350 -4312 -2288 -4292
rect -2350 -4346 -2340 -4312
rect -2306 -4346 -2288 -4312
rect -2350 -4376 -2288 -4346
rect -2258 -4306 -2189 -4292
rect -2258 -4340 -2247 -4306
rect -2213 -4340 -2189 -4306
rect -2258 -4376 -2189 -4340
rect -2159 -4330 -2049 -4292
rect -2159 -4364 -2093 -4330
rect -2059 -4364 -2049 -4330
rect -2159 -4376 -2049 -4364
rect -2019 -4314 -1952 -4292
rect -2019 -4348 -1996 -4314
rect -1962 -4348 -1952 -4314
rect -2019 -4376 -1952 -4348
rect -1922 -4330 -1870 -4292
rect -1922 -4364 -1912 -4330
rect -1878 -4364 -1870 -4330
rect -1922 -4376 -1870 -4364
rect -1807 -4304 -1755 -4292
rect -1807 -4338 -1799 -4304
rect -1765 -4338 -1755 -4304
rect -2617 -4414 -2607 -4380
rect -2573 -4414 -2565 -4380
rect -2617 -4426 -2565 -4414
rect -2900 -4492 -2848 -4442
rect -1807 -4460 -1755 -4338
rect -1725 -4312 -1656 -4292
rect -1725 -4346 -1711 -4312
rect -1677 -4346 -1656 -4312
rect -1725 -4376 -1656 -4346
rect -1626 -4305 -1570 -4292
rect -1626 -4339 -1614 -4305
rect -1580 -4339 -1570 -4305
rect -1626 -4376 -1570 -4339
rect -1540 -4376 -1486 -4292
rect -1456 -4304 -1378 -4292
rect -1456 -4338 -1422 -4304
rect -1388 -4338 -1378 -4304
rect -1456 -4376 -1378 -4338
rect -1348 -4330 -1294 -4292
rect -1348 -4364 -1338 -4330
rect -1304 -4364 -1294 -4330
rect -1348 -4376 -1294 -4364
rect -1264 -4304 -1130 -4292
rect -1264 -4338 -1252 -4304
rect -1218 -4338 -1174 -4304
rect -1140 -4338 -1130 -4304
rect -1264 -4376 -1130 -4338
rect -1725 -4460 -1671 -4376
rect -1180 -4492 -1130 -4376
rect -1100 -4312 -1044 -4292
rect -1100 -4346 -1090 -4312
rect -1056 -4346 -1044 -4312
rect -1100 -4380 -1044 -4346
rect -1100 -4414 -1090 -4380
rect -1056 -4414 -1044 -4380
rect -1100 -4448 -1044 -4414
rect -963 -4304 -911 -4292
rect -963 -4338 -955 -4304
rect -921 -4338 -911 -4304
rect -963 -4372 -911 -4338
rect -963 -4406 -955 -4372
rect -921 -4406 -911 -4372
rect -963 -4420 -911 -4406
rect -881 -4304 -814 -4292
rect -881 -4338 -858 -4304
rect -824 -4338 -814 -4304
rect -881 -4372 -814 -4338
rect -881 -4406 -858 -4372
rect -824 -4406 -814 -4372
rect -881 -4420 -814 -4406
rect -1100 -4482 -1090 -4448
rect -1056 -4482 -1044 -4448
rect -1100 -4492 -1044 -4482
rect -866 -4440 -814 -4420
rect -866 -4474 -858 -4440
rect -824 -4474 -814 -4440
rect -866 -4492 -814 -4474
rect -784 -4340 -732 -4292
rect -784 -4374 -774 -4340
rect -740 -4374 -732 -4340
rect -784 -4408 -732 -4374
rect -784 -4442 -774 -4408
rect -740 -4442 -732 -4408
rect -667 -4312 -615 -4298
rect -667 -4346 -659 -4312
rect -625 -4346 -615 -4312
rect -667 -4380 -615 -4346
rect -667 -4414 -659 -4380
rect -625 -4414 -615 -4380
rect -667 -4426 -615 -4414
rect -585 -4328 -531 -4298
rect -585 -4362 -575 -4328
rect -541 -4362 -531 -4328
rect -585 -4426 -531 -4362
rect -501 -4312 -449 -4298
rect -501 -4346 -491 -4312
rect -457 -4346 -449 -4312
rect -501 -4380 -449 -4346
rect -316 -4304 -264 -4292
rect -316 -4338 -308 -4304
rect -274 -4338 -264 -4304
rect -316 -4376 -264 -4338
rect -234 -4312 -172 -4292
rect -234 -4346 -224 -4312
rect -190 -4346 -172 -4312
rect -234 -4376 -172 -4346
rect -142 -4306 -73 -4292
rect -142 -4340 -131 -4306
rect -97 -4340 -73 -4306
rect -142 -4376 -73 -4340
rect -43 -4330 67 -4292
rect -43 -4364 23 -4330
rect 57 -4364 67 -4330
rect -43 -4376 67 -4364
rect 97 -4314 164 -4292
rect 97 -4348 120 -4314
rect 154 -4348 164 -4314
rect 97 -4376 164 -4348
rect 194 -4330 246 -4292
rect 194 -4364 204 -4330
rect 238 -4364 246 -4330
rect 194 -4376 246 -4364
rect 309 -4304 361 -4292
rect 309 -4338 317 -4304
rect 351 -4338 361 -4304
rect -501 -4414 -491 -4380
rect -457 -4414 -449 -4380
rect -501 -4426 -449 -4414
rect -784 -4492 -732 -4442
rect 309 -4460 361 -4338
rect 391 -4312 460 -4292
rect 391 -4346 405 -4312
rect 439 -4346 460 -4312
rect 391 -4376 460 -4346
rect 490 -4305 546 -4292
rect 490 -4339 502 -4305
rect 536 -4339 546 -4305
rect 490 -4376 546 -4339
rect 576 -4376 630 -4292
rect 660 -4304 738 -4292
rect 660 -4338 694 -4304
rect 728 -4338 738 -4304
rect 660 -4376 738 -4338
rect 768 -4330 822 -4292
rect 768 -4364 778 -4330
rect 812 -4364 822 -4330
rect 768 -4376 822 -4364
rect 852 -4304 986 -4292
rect 852 -4338 864 -4304
rect 898 -4338 942 -4304
rect 976 -4338 986 -4304
rect 852 -4376 986 -4338
rect 391 -4460 445 -4376
rect 936 -4492 986 -4376
rect 1016 -4312 1072 -4292
rect 1016 -4346 1026 -4312
rect 1060 -4346 1072 -4312
rect 1016 -4380 1072 -4346
rect 1016 -4414 1026 -4380
rect 1060 -4414 1072 -4380
rect 1016 -4448 1072 -4414
rect 1153 -4304 1205 -4292
rect 1153 -4338 1161 -4304
rect 1195 -4338 1205 -4304
rect 1153 -4372 1205 -4338
rect 1153 -4406 1161 -4372
rect 1195 -4406 1205 -4372
rect 1153 -4420 1205 -4406
rect 1235 -4304 1302 -4292
rect 1235 -4338 1258 -4304
rect 1292 -4338 1302 -4304
rect 1235 -4372 1302 -4338
rect 1235 -4406 1258 -4372
rect 1292 -4406 1302 -4372
rect 1235 -4420 1302 -4406
rect 1016 -4482 1026 -4448
rect 1060 -4482 1072 -4448
rect 1016 -4492 1072 -4482
rect 1250 -4440 1302 -4420
rect 1250 -4474 1258 -4440
rect 1292 -4474 1302 -4440
rect 1250 -4492 1302 -4474
rect 1332 -4340 1384 -4292
rect 1332 -4374 1342 -4340
rect 1376 -4374 1384 -4340
rect 1332 -4408 1384 -4374
rect 1332 -4442 1342 -4408
rect 1376 -4442 1384 -4408
rect 1449 -4312 1501 -4298
rect 1449 -4346 1457 -4312
rect 1491 -4346 1501 -4312
rect 1449 -4380 1501 -4346
rect 1449 -4414 1457 -4380
rect 1491 -4414 1501 -4380
rect 1449 -4426 1501 -4414
rect 1531 -4328 1585 -4298
rect 1531 -4362 1541 -4328
rect 1575 -4362 1585 -4328
rect 1531 -4426 1585 -4362
rect 1615 -4312 1667 -4298
rect 1615 -4346 1625 -4312
rect 1659 -4346 1667 -4312
rect 1615 -4380 1667 -4346
rect 1800 -4304 1852 -4292
rect 1800 -4338 1808 -4304
rect 1842 -4338 1852 -4304
rect 1800 -4376 1852 -4338
rect 1882 -4312 1944 -4292
rect 1882 -4346 1892 -4312
rect 1926 -4346 1944 -4312
rect 1882 -4376 1944 -4346
rect 1974 -4306 2043 -4292
rect 1974 -4340 1985 -4306
rect 2019 -4340 2043 -4306
rect 1974 -4376 2043 -4340
rect 2073 -4330 2183 -4292
rect 2073 -4364 2139 -4330
rect 2173 -4364 2183 -4330
rect 2073 -4376 2183 -4364
rect 2213 -4314 2280 -4292
rect 2213 -4348 2236 -4314
rect 2270 -4348 2280 -4314
rect 2213 -4376 2280 -4348
rect 2310 -4330 2362 -4292
rect 2310 -4364 2320 -4330
rect 2354 -4364 2362 -4330
rect 2310 -4376 2362 -4364
rect 2425 -4304 2477 -4292
rect 2425 -4338 2433 -4304
rect 2467 -4338 2477 -4304
rect 1615 -4414 1625 -4380
rect 1659 -4414 1667 -4380
rect 1615 -4426 1667 -4414
rect 1332 -4492 1384 -4442
rect 2425 -4460 2477 -4338
rect 2507 -4312 2576 -4292
rect 2507 -4346 2521 -4312
rect 2555 -4346 2576 -4312
rect 2507 -4376 2576 -4346
rect 2606 -4305 2662 -4292
rect 2606 -4339 2618 -4305
rect 2652 -4339 2662 -4305
rect 2606 -4376 2662 -4339
rect 2692 -4376 2746 -4292
rect 2776 -4304 2854 -4292
rect 2776 -4338 2810 -4304
rect 2844 -4338 2854 -4304
rect 2776 -4376 2854 -4338
rect 2884 -4330 2938 -4292
rect 2884 -4364 2894 -4330
rect 2928 -4364 2938 -4330
rect 2884 -4376 2938 -4364
rect 2968 -4304 3102 -4292
rect 2968 -4338 2980 -4304
rect 3014 -4338 3058 -4304
rect 3092 -4338 3102 -4304
rect 2968 -4376 3102 -4338
rect 2507 -4460 2561 -4376
rect 3052 -4492 3102 -4376
rect 3132 -4312 3188 -4292
rect 3132 -4346 3142 -4312
rect 3176 -4346 3188 -4312
rect 3132 -4380 3188 -4346
rect 3132 -4414 3142 -4380
rect 3176 -4414 3188 -4380
rect 3132 -4448 3188 -4414
rect 3269 -4304 3321 -4292
rect 3269 -4338 3277 -4304
rect 3311 -4338 3321 -4304
rect 3269 -4372 3321 -4338
rect 3269 -4406 3277 -4372
rect 3311 -4406 3321 -4372
rect 3269 -4420 3321 -4406
rect 3351 -4304 3418 -4292
rect 3351 -4338 3374 -4304
rect 3408 -4338 3418 -4304
rect 3351 -4372 3418 -4338
rect 3351 -4406 3374 -4372
rect 3408 -4406 3418 -4372
rect 3351 -4420 3418 -4406
rect 3132 -4482 3142 -4448
rect 3176 -4482 3188 -4448
rect 3132 -4492 3188 -4482
rect 3366 -4440 3418 -4420
rect 3366 -4474 3374 -4440
rect 3408 -4474 3418 -4440
rect 3366 -4492 3418 -4474
rect 3448 -4340 3500 -4292
rect 3448 -4374 3458 -4340
rect 3492 -4374 3500 -4340
rect 3448 -4408 3500 -4374
rect 3448 -4442 3458 -4408
rect 3492 -4442 3500 -4408
rect 3565 -4312 3617 -4298
rect 3565 -4346 3573 -4312
rect 3607 -4346 3617 -4312
rect 3565 -4380 3617 -4346
rect 3565 -4414 3573 -4380
rect 3607 -4414 3617 -4380
rect 3565 -4426 3617 -4414
rect 3647 -4328 3701 -4298
rect 3647 -4362 3657 -4328
rect 3691 -4362 3701 -4328
rect 3647 -4426 3701 -4362
rect 3731 -4312 3783 -4298
rect 3731 -4346 3741 -4312
rect 3775 -4346 3783 -4312
rect 3731 -4380 3783 -4346
rect 3916 -4304 3968 -4292
rect 3916 -4338 3924 -4304
rect 3958 -4338 3968 -4304
rect 3916 -4376 3968 -4338
rect 3998 -4312 4060 -4292
rect 3998 -4346 4008 -4312
rect 4042 -4346 4060 -4312
rect 3998 -4376 4060 -4346
rect 4090 -4306 4159 -4292
rect 4090 -4340 4101 -4306
rect 4135 -4340 4159 -4306
rect 4090 -4376 4159 -4340
rect 4189 -4330 4299 -4292
rect 4189 -4364 4255 -4330
rect 4289 -4364 4299 -4330
rect 4189 -4376 4299 -4364
rect 4329 -4314 4396 -4292
rect 4329 -4348 4352 -4314
rect 4386 -4348 4396 -4314
rect 4329 -4376 4396 -4348
rect 4426 -4330 4478 -4292
rect 4426 -4364 4436 -4330
rect 4470 -4364 4478 -4330
rect 4426 -4376 4478 -4364
rect 4541 -4304 4593 -4292
rect 4541 -4338 4549 -4304
rect 4583 -4338 4593 -4304
rect 3731 -4414 3741 -4380
rect 3775 -4414 3783 -4380
rect 3731 -4426 3783 -4414
rect 3448 -4492 3500 -4442
rect 4541 -4460 4593 -4338
rect 4623 -4312 4692 -4292
rect 4623 -4346 4637 -4312
rect 4671 -4346 4692 -4312
rect 4623 -4376 4692 -4346
rect 4722 -4305 4778 -4292
rect 4722 -4339 4734 -4305
rect 4768 -4339 4778 -4305
rect 4722 -4376 4778 -4339
rect 4808 -4376 4862 -4292
rect 4892 -4304 4970 -4292
rect 4892 -4338 4926 -4304
rect 4960 -4338 4970 -4304
rect 4892 -4376 4970 -4338
rect 5000 -4330 5054 -4292
rect 5000 -4364 5010 -4330
rect 5044 -4364 5054 -4330
rect 5000 -4376 5054 -4364
rect 5084 -4304 5218 -4292
rect 5084 -4338 5096 -4304
rect 5130 -4338 5174 -4304
rect 5208 -4338 5218 -4304
rect 5084 -4376 5218 -4338
rect 4623 -4460 4677 -4376
rect 5168 -4492 5218 -4376
rect 5248 -4312 5304 -4292
rect 5248 -4346 5258 -4312
rect 5292 -4346 5304 -4312
rect 5248 -4380 5304 -4346
rect 5248 -4414 5258 -4380
rect 5292 -4414 5304 -4380
rect 5248 -4448 5304 -4414
rect 5385 -4304 5437 -4292
rect 5385 -4338 5393 -4304
rect 5427 -4338 5437 -4304
rect 5385 -4372 5437 -4338
rect 5385 -4406 5393 -4372
rect 5427 -4406 5437 -4372
rect 5385 -4420 5437 -4406
rect 5467 -4304 5534 -4292
rect 5467 -4338 5490 -4304
rect 5524 -4338 5534 -4304
rect 5467 -4372 5534 -4338
rect 5467 -4406 5490 -4372
rect 5524 -4406 5534 -4372
rect 5467 -4420 5534 -4406
rect 5248 -4482 5258 -4448
rect 5292 -4482 5304 -4448
rect 5248 -4492 5304 -4482
rect 5482 -4440 5534 -4420
rect 5482 -4474 5490 -4440
rect 5524 -4474 5534 -4440
rect 5482 -4492 5534 -4474
rect 5564 -4340 5616 -4292
rect 5564 -4374 5574 -4340
rect 5608 -4374 5616 -4340
rect 5564 -4408 5616 -4374
rect 5564 -4442 5574 -4408
rect 5608 -4442 5616 -4408
rect 5681 -4312 5733 -4298
rect 5681 -4346 5689 -4312
rect 5723 -4346 5733 -4312
rect 5681 -4380 5733 -4346
rect 5681 -4414 5689 -4380
rect 5723 -4414 5733 -4380
rect 5681 -4426 5733 -4414
rect 5763 -4328 5817 -4298
rect 5763 -4362 5773 -4328
rect 5807 -4362 5817 -4328
rect 5763 -4426 5817 -4362
rect 5847 -4312 5899 -4298
rect 5847 -4346 5857 -4312
rect 5891 -4346 5899 -4312
rect 5847 -4380 5899 -4346
rect 6032 -4304 6084 -4292
rect 6032 -4338 6040 -4304
rect 6074 -4338 6084 -4304
rect 6032 -4376 6084 -4338
rect 6114 -4312 6176 -4292
rect 6114 -4346 6124 -4312
rect 6158 -4346 6176 -4312
rect 6114 -4376 6176 -4346
rect 6206 -4306 6275 -4292
rect 6206 -4340 6217 -4306
rect 6251 -4340 6275 -4306
rect 6206 -4376 6275 -4340
rect 6305 -4330 6415 -4292
rect 6305 -4364 6371 -4330
rect 6405 -4364 6415 -4330
rect 6305 -4376 6415 -4364
rect 6445 -4314 6512 -4292
rect 6445 -4348 6468 -4314
rect 6502 -4348 6512 -4314
rect 6445 -4376 6512 -4348
rect 6542 -4330 6594 -4292
rect 6542 -4364 6552 -4330
rect 6586 -4364 6594 -4330
rect 6542 -4376 6594 -4364
rect 6657 -4304 6709 -4292
rect 6657 -4338 6665 -4304
rect 6699 -4338 6709 -4304
rect 5847 -4414 5857 -4380
rect 5891 -4414 5899 -4380
rect 5847 -4426 5899 -4414
rect 5564 -4492 5616 -4442
rect 6657 -4460 6709 -4338
rect 6739 -4312 6808 -4292
rect 6739 -4346 6753 -4312
rect 6787 -4346 6808 -4312
rect 6739 -4376 6808 -4346
rect 6838 -4305 6894 -4292
rect 6838 -4339 6850 -4305
rect 6884 -4339 6894 -4305
rect 6838 -4376 6894 -4339
rect 6924 -4376 6978 -4292
rect 7008 -4304 7086 -4292
rect 7008 -4338 7042 -4304
rect 7076 -4338 7086 -4304
rect 7008 -4376 7086 -4338
rect 7116 -4330 7170 -4292
rect 7116 -4364 7126 -4330
rect 7160 -4364 7170 -4330
rect 7116 -4376 7170 -4364
rect 7200 -4304 7334 -4292
rect 7200 -4338 7212 -4304
rect 7246 -4338 7290 -4304
rect 7324 -4338 7334 -4304
rect 7200 -4376 7334 -4338
rect 6739 -4460 6793 -4376
rect 7284 -4492 7334 -4376
rect 7364 -4312 7420 -4292
rect 7364 -4346 7374 -4312
rect 7408 -4346 7420 -4312
rect 7364 -4380 7420 -4346
rect 7364 -4414 7374 -4380
rect 7408 -4414 7420 -4380
rect 7364 -4448 7420 -4414
rect 7501 -4304 7553 -4292
rect 7501 -4338 7509 -4304
rect 7543 -4338 7553 -4304
rect 7501 -4372 7553 -4338
rect 7501 -4406 7509 -4372
rect 7543 -4406 7553 -4372
rect 7501 -4420 7553 -4406
rect 7583 -4304 7650 -4292
rect 7583 -4338 7606 -4304
rect 7640 -4338 7650 -4304
rect 7583 -4372 7650 -4338
rect 7583 -4406 7606 -4372
rect 7640 -4406 7650 -4372
rect 7583 -4420 7650 -4406
rect 7364 -4482 7374 -4448
rect 7408 -4482 7420 -4448
rect 7364 -4492 7420 -4482
rect 7598 -4440 7650 -4420
rect 7598 -4474 7606 -4440
rect 7640 -4474 7650 -4440
rect 7598 -4492 7650 -4474
rect 7680 -4340 7732 -4292
rect 7680 -4374 7690 -4340
rect 7724 -4374 7732 -4340
rect 7680 -4408 7732 -4374
rect 7680 -4442 7690 -4408
rect 7724 -4442 7732 -4408
rect 7797 -4312 7849 -4298
rect 7797 -4346 7805 -4312
rect 7839 -4346 7849 -4312
rect 7797 -4380 7849 -4346
rect 7797 -4414 7805 -4380
rect 7839 -4414 7849 -4380
rect 7797 -4426 7849 -4414
rect 7879 -4328 7933 -4298
rect 7879 -4362 7889 -4328
rect 7923 -4362 7933 -4328
rect 7879 -4426 7933 -4362
rect 7963 -4312 8015 -4298
rect 7963 -4346 7973 -4312
rect 8007 -4346 8015 -4312
rect 7963 -4380 8015 -4346
rect 8148 -4304 8200 -4292
rect 8148 -4338 8156 -4304
rect 8190 -4338 8200 -4304
rect 8148 -4376 8200 -4338
rect 8230 -4312 8292 -4292
rect 8230 -4346 8240 -4312
rect 8274 -4346 8292 -4312
rect 8230 -4376 8292 -4346
rect 8322 -4306 8391 -4292
rect 8322 -4340 8333 -4306
rect 8367 -4340 8391 -4306
rect 8322 -4376 8391 -4340
rect 8421 -4330 8531 -4292
rect 8421 -4364 8487 -4330
rect 8521 -4364 8531 -4330
rect 8421 -4376 8531 -4364
rect 8561 -4314 8628 -4292
rect 8561 -4348 8584 -4314
rect 8618 -4348 8628 -4314
rect 8561 -4376 8628 -4348
rect 8658 -4330 8710 -4292
rect 8658 -4364 8668 -4330
rect 8702 -4364 8710 -4330
rect 8658 -4376 8710 -4364
rect 8773 -4304 8825 -4292
rect 8773 -4338 8781 -4304
rect 8815 -4338 8825 -4304
rect 7963 -4414 7973 -4380
rect 8007 -4414 8015 -4380
rect 7963 -4426 8015 -4414
rect 7680 -4492 7732 -4442
rect 8773 -4460 8825 -4338
rect 8855 -4312 8924 -4292
rect 8855 -4346 8869 -4312
rect 8903 -4346 8924 -4312
rect 8855 -4376 8924 -4346
rect 8954 -4305 9010 -4292
rect 8954 -4339 8966 -4305
rect 9000 -4339 9010 -4305
rect 8954 -4376 9010 -4339
rect 9040 -4376 9094 -4292
rect 9124 -4304 9202 -4292
rect 9124 -4338 9158 -4304
rect 9192 -4338 9202 -4304
rect 9124 -4376 9202 -4338
rect 9232 -4330 9286 -4292
rect 9232 -4364 9242 -4330
rect 9276 -4364 9286 -4330
rect 9232 -4376 9286 -4364
rect 9316 -4304 9450 -4292
rect 9316 -4338 9328 -4304
rect 9362 -4338 9406 -4304
rect 9440 -4338 9450 -4304
rect 9316 -4376 9450 -4338
rect 8855 -4460 8909 -4376
rect 9400 -4492 9450 -4376
rect 9480 -4312 9536 -4292
rect 9480 -4346 9490 -4312
rect 9524 -4346 9536 -4312
rect 9480 -4380 9536 -4346
rect 9480 -4414 9490 -4380
rect 9524 -4414 9536 -4380
rect 9480 -4448 9536 -4414
rect 9617 -4304 9669 -4292
rect 9617 -4338 9625 -4304
rect 9659 -4338 9669 -4304
rect 9617 -4372 9669 -4338
rect 9617 -4406 9625 -4372
rect 9659 -4406 9669 -4372
rect 9617 -4420 9669 -4406
rect 9699 -4304 9766 -4292
rect 9699 -4338 9722 -4304
rect 9756 -4338 9766 -4304
rect 9699 -4372 9766 -4338
rect 9699 -4406 9722 -4372
rect 9756 -4406 9766 -4372
rect 9699 -4420 9766 -4406
rect 9480 -4482 9490 -4448
rect 9524 -4482 9536 -4448
rect 9480 -4492 9536 -4482
rect 9714 -4440 9766 -4420
rect 9714 -4474 9722 -4440
rect 9756 -4474 9766 -4440
rect 9714 -4492 9766 -4474
rect 9796 -4340 9848 -4292
rect 9796 -4374 9806 -4340
rect 9840 -4374 9848 -4340
rect 9796 -4408 9848 -4374
rect 9796 -4442 9806 -4408
rect 9840 -4442 9848 -4408
rect 9913 -4312 9965 -4298
rect 9913 -4346 9921 -4312
rect 9955 -4346 9965 -4312
rect 9913 -4380 9965 -4346
rect 9913 -4414 9921 -4380
rect 9955 -4414 9965 -4380
rect 9913 -4426 9965 -4414
rect 9995 -4328 10049 -4298
rect 9995 -4362 10005 -4328
rect 10039 -4362 10049 -4328
rect 9995 -4426 10049 -4362
rect 10079 -4312 10131 -4298
rect 10079 -4346 10089 -4312
rect 10123 -4346 10131 -4312
rect 10079 -4380 10131 -4346
rect 10264 -4304 10316 -4292
rect 10264 -4338 10272 -4304
rect 10306 -4338 10316 -4304
rect 10264 -4376 10316 -4338
rect 10346 -4312 10408 -4292
rect 10346 -4346 10356 -4312
rect 10390 -4346 10408 -4312
rect 10346 -4376 10408 -4346
rect 10438 -4306 10507 -4292
rect 10438 -4340 10449 -4306
rect 10483 -4340 10507 -4306
rect 10438 -4376 10507 -4340
rect 10537 -4330 10647 -4292
rect 10537 -4364 10603 -4330
rect 10637 -4364 10647 -4330
rect 10537 -4376 10647 -4364
rect 10677 -4314 10744 -4292
rect 10677 -4348 10700 -4314
rect 10734 -4348 10744 -4314
rect 10677 -4376 10744 -4348
rect 10774 -4330 10826 -4292
rect 10774 -4364 10784 -4330
rect 10818 -4364 10826 -4330
rect 10774 -4376 10826 -4364
rect 10889 -4304 10941 -4292
rect 10889 -4338 10897 -4304
rect 10931 -4338 10941 -4304
rect 10079 -4414 10089 -4380
rect 10123 -4414 10131 -4380
rect 10079 -4426 10131 -4414
rect 9796 -4492 9848 -4442
rect 10889 -4460 10941 -4338
rect 10971 -4312 11040 -4292
rect 10971 -4346 10985 -4312
rect 11019 -4346 11040 -4312
rect 10971 -4376 11040 -4346
rect 11070 -4305 11126 -4292
rect 11070 -4339 11082 -4305
rect 11116 -4339 11126 -4305
rect 11070 -4376 11126 -4339
rect 11156 -4376 11210 -4292
rect 11240 -4304 11318 -4292
rect 11240 -4338 11274 -4304
rect 11308 -4338 11318 -4304
rect 11240 -4376 11318 -4338
rect 11348 -4330 11402 -4292
rect 11348 -4364 11358 -4330
rect 11392 -4364 11402 -4330
rect 11348 -4376 11402 -4364
rect 11432 -4304 11566 -4292
rect 11432 -4338 11444 -4304
rect 11478 -4338 11522 -4304
rect 11556 -4338 11566 -4304
rect 11432 -4376 11566 -4338
rect 10971 -4460 11025 -4376
rect 11516 -4492 11566 -4376
rect 11596 -4312 11652 -4292
rect 11596 -4346 11606 -4312
rect 11640 -4346 11652 -4312
rect 11596 -4380 11652 -4346
rect 11596 -4414 11606 -4380
rect 11640 -4414 11652 -4380
rect 11596 -4448 11652 -4414
rect 11733 -4304 11785 -4292
rect 11733 -4338 11741 -4304
rect 11775 -4338 11785 -4304
rect 11733 -4372 11785 -4338
rect 11733 -4406 11741 -4372
rect 11775 -4406 11785 -4372
rect 11733 -4420 11785 -4406
rect 11815 -4304 11882 -4292
rect 11815 -4338 11838 -4304
rect 11872 -4338 11882 -4304
rect 11815 -4372 11882 -4338
rect 11815 -4406 11838 -4372
rect 11872 -4406 11882 -4372
rect 11815 -4420 11882 -4406
rect 11596 -4482 11606 -4448
rect 11640 -4482 11652 -4448
rect 11596 -4492 11652 -4482
rect 11830 -4440 11882 -4420
rect 11830 -4474 11838 -4440
rect 11872 -4474 11882 -4440
rect 11830 -4492 11882 -4474
rect 11912 -4340 11964 -4292
rect 11912 -4374 11922 -4340
rect 11956 -4374 11964 -4340
rect 11912 -4408 11964 -4374
rect 11912 -4442 11922 -4408
rect 11956 -4442 11964 -4408
rect 12029 -4312 12081 -4298
rect 12029 -4346 12037 -4312
rect 12071 -4346 12081 -4312
rect 12029 -4380 12081 -4346
rect 12029 -4414 12037 -4380
rect 12071 -4414 12081 -4380
rect 12029 -4426 12081 -4414
rect 12111 -4328 12165 -4298
rect 12111 -4362 12121 -4328
rect 12155 -4362 12165 -4328
rect 12111 -4426 12165 -4362
rect 12195 -4312 12247 -4298
rect 12195 -4346 12205 -4312
rect 12239 -4346 12247 -4312
rect 12195 -4380 12247 -4346
rect 12380 -4304 12432 -4292
rect 12380 -4338 12388 -4304
rect 12422 -4338 12432 -4304
rect 12380 -4376 12432 -4338
rect 12462 -4312 12524 -4292
rect 12462 -4346 12472 -4312
rect 12506 -4346 12524 -4312
rect 12462 -4376 12524 -4346
rect 12554 -4306 12623 -4292
rect 12554 -4340 12565 -4306
rect 12599 -4340 12623 -4306
rect 12554 -4376 12623 -4340
rect 12653 -4330 12763 -4292
rect 12653 -4364 12719 -4330
rect 12753 -4364 12763 -4330
rect 12653 -4376 12763 -4364
rect 12793 -4314 12860 -4292
rect 12793 -4348 12816 -4314
rect 12850 -4348 12860 -4314
rect 12793 -4376 12860 -4348
rect 12890 -4330 12942 -4292
rect 12890 -4364 12900 -4330
rect 12934 -4364 12942 -4330
rect 12890 -4376 12942 -4364
rect 13005 -4304 13057 -4292
rect 13005 -4338 13013 -4304
rect 13047 -4338 13057 -4304
rect 12195 -4414 12205 -4380
rect 12239 -4414 12247 -4380
rect 12195 -4426 12247 -4414
rect 11912 -4492 11964 -4442
rect 13005 -4460 13057 -4338
rect 13087 -4312 13156 -4292
rect 13087 -4346 13101 -4312
rect 13135 -4346 13156 -4312
rect 13087 -4376 13156 -4346
rect 13186 -4305 13242 -4292
rect 13186 -4339 13198 -4305
rect 13232 -4339 13242 -4305
rect 13186 -4376 13242 -4339
rect 13272 -4376 13326 -4292
rect 13356 -4304 13434 -4292
rect 13356 -4338 13390 -4304
rect 13424 -4338 13434 -4304
rect 13356 -4376 13434 -4338
rect 13464 -4330 13518 -4292
rect 13464 -4364 13474 -4330
rect 13508 -4364 13518 -4330
rect 13464 -4376 13518 -4364
rect 13548 -4304 13682 -4292
rect 13548 -4338 13560 -4304
rect 13594 -4338 13638 -4304
rect 13672 -4338 13682 -4304
rect 13548 -4376 13682 -4338
rect 13087 -4460 13141 -4376
rect 13632 -4492 13682 -4376
rect 13712 -4312 13768 -4292
rect 13712 -4346 13722 -4312
rect 13756 -4346 13768 -4312
rect 13712 -4380 13768 -4346
rect 13712 -4414 13722 -4380
rect 13756 -4414 13768 -4380
rect 13712 -4448 13768 -4414
rect 13849 -4304 13901 -4292
rect 13849 -4338 13857 -4304
rect 13891 -4338 13901 -4304
rect 13849 -4372 13901 -4338
rect 13849 -4406 13857 -4372
rect 13891 -4406 13901 -4372
rect 13849 -4420 13901 -4406
rect 13931 -4304 13998 -4292
rect 13931 -4338 13954 -4304
rect 13988 -4338 13998 -4304
rect 13931 -4372 13998 -4338
rect 13931 -4406 13954 -4372
rect 13988 -4406 13998 -4372
rect 13931 -4420 13998 -4406
rect 13712 -4482 13722 -4448
rect 13756 -4482 13768 -4448
rect 13712 -4492 13768 -4482
rect 13946 -4440 13998 -4420
rect 13946 -4474 13954 -4440
rect 13988 -4474 13998 -4440
rect 13946 -4492 13998 -4474
rect 14028 -4340 14080 -4292
rect 14028 -4374 14038 -4340
rect 14072 -4374 14080 -4340
rect 14028 -4408 14080 -4374
rect 14028 -4442 14038 -4408
rect 14072 -4442 14080 -4408
rect 14145 -4312 14197 -4298
rect 14145 -4346 14153 -4312
rect 14187 -4346 14197 -4312
rect 14145 -4380 14197 -4346
rect 14145 -4414 14153 -4380
rect 14187 -4414 14197 -4380
rect 14145 -4426 14197 -4414
rect 14227 -4328 14281 -4298
rect 14227 -4362 14237 -4328
rect 14271 -4362 14281 -4328
rect 14227 -4426 14281 -4362
rect 14311 -4312 14363 -4298
rect 14311 -4346 14321 -4312
rect 14355 -4346 14363 -4312
rect 14311 -4380 14363 -4346
rect 14496 -4304 14548 -4292
rect 14496 -4338 14504 -4304
rect 14538 -4338 14548 -4304
rect 14496 -4376 14548 -4338
rect 14578 -4312 14640 -4292
rect 14578 -4346 14588 -4312
rect 14622 -4346 14640 -4312
rect 14578 -4376 14640 -4346
rect 14670 -4306 14739 -4292
rect 14670 -4340 14681 -4306
rect 14715 -4340 14739 -4306
rect 14670 -4376 14739 -4340
rect 14769 -4330 14879 -4292
rect 14769 -4364 14835 -4330
rect 14869 -4364 14879 -4330
rect 14769 -4376 14879 -4364
rect 14909 -4314 14976 -4292
rect 14909 -4348 14932 -4314
rect 14966 -4348 14976 -4314
rect 14909 -4376 14976 -4348
rect 15006 -4330 15058 -4292
rect 15006 -4364 15016 -4330
rect 15050 -4364 15058 -4330
rect 15006 -4376 15058 -4364
rect 15121 -4304 15173 -4292
rect 15121 -4338 15129 -4304
rect 15163 -4338 15173 -4304
rect 14311 -4414 14321 -4380
rect 14355 -4414 14363 -4380
rect 14311 -4426 14363 -4414
rect 14028 -4492 14080 -4442
rect 15121 -4460 15173 -4338
rect 15203 -4312 15272 -4292
rect 15203 -4346 15217 -4312
rect 15251 -4346 15272 -4312
rect 15203 -4376 15272 -4346
rect 15302 -4305 15358 -4292
rect 15302 -4339 15314 -4305
rect 15348 -4339 15358 -4305
rect 15302 -4376 15358 -4339
rect 15388 -4376 15442 -4292
rect 15472 -4304 15550 -4292
rect 15472 -4338 15506 -4304
rect 15540 -4338 15550 -4304
rect 15472 -4376 15550 -4338
rect 15580 -4330 15634 -4292
rect 15580 -4364 15590 -4330
rect 15624 -4364 15634 -4330
rect 15580 -4376 15634 -4364
rect 15664 -4304 15798 -4292
rect 15664 -4338 15676 -4304
rect 15710 -4338 15754 -4304
rect 15788 -4338 15798 -4304
rect 15664 -4376 15798 -4338
rect 15203 -4460 15257 -4376
rect 15748 -4492 15798 -4376
rect 15828 -4312 15884 -4292
rect 15828 -4346 15838 -4312
rect 15872 -4346 15884 -4312
rect 15828 -4380 15884 -4346
rect 15828 -4414 15838 -4380
rect 15872 -4414 15884 -4380
rect 15828 -4448 15884 -4414
rect 15965 -4304 16017 -4292
rect 15965 -4338 15973 -4304
rect 16007 -4338 16017 -4304
rect 15965 -4372 16017 -4338
rect 15965 -4406 15973 -4372
rect 16007 -4406 16017 -4372
rect 15965 -4420 16017 -4406
rect 16047 -4304 16114 -4292
rect 16047 -4338 16070 -4304
rect 16104 -4338 16114 -4304
rect 16047 -4372 16114 -4338
rect 16047 -4406 16070 -4372
rect 16104 -4406 16114 -4372
rect 16047 -4420 16114 -4406
rect 15828 -4482 15838 -4448
rect 15872 -4482 15884 -4448
rect 15828 -4492 15884 -4482
rect 16062 -4440 16114 -4420
rect 16062 -4474 16070 -4440
rect 16104 -4474 16114 -4440
rect 16062 -4492 16114 -4474
rect 16144 -4340 16196 -4292
rect 16144 -4374 16154 -4340
rect 16188 -4374 16196 -4340
rect 16144 -4408 16196 -4374
rect 16144 -4442 16154 -4408
rect 16188 -4442 16196 -4408
rect 16261 -4312 16313 -4298
rect 16261 -4346 16269 -4312
rect 16303 -4346 16313 -4312
rect 16261 -4380 16313 -4346
rect 16261 -4414 16269 -4380
rect 16303 -4414 16313 -4380
rect 16261 -4426 16313 -4414
rect 16343 -4328 16397 -4298
rect 16343 -4362 16353 -4328
rect 16387 -4362 16397 -4328
rect 16343 -4426 16397 -4362
rect 16427 -4312 16479 -4298
rect 16427 -4346 16437 -4312
rect 16471 -4346 16479 -4312
rect 16427 -4380 16479 -4346
rect 16612 -4304 16664 -4292
rect 16612 -4338 16620 -4304
rect 16654 -4338 16664 -4304
rect 16612 -4376 16664 -4338
rect 16694 -4312 16756 -4292
rect 16694 -4346 16704 -4312
rect 16738 -4346 16756 -4312
rect 16694 -4376 16756 -4346
rect 16786 -4306 16855 -4292
rect 16786 -4340 16797 -4306
rect 16831 -4340 16855 -4306
rect 16786 -4376 16855 -4340
rect 16885 -4330 16995 -4292
rect 16885 -4364 16951 -4330
rect 16985 -4364 16995 -4330
rect 16885 -4376 16995 -4364
rect 17025 -4314 17092 -4292
rect 17025 -4348 17048 -4314
rect 17082 -4348 17092 -4314
rect 17025 -4376 17092 -4348
rect 17122 -4330 17174 -4292
rect 17122 -4364 17132 -4330
rect 17166 -4364 17174 -4330
rect 17122 -4376 17174 -4364
rect 17237 -4304 17289 -4292
rect 17237 -4338 17245 -4304
rect 17279 -4338 17289 -4304
rect 16427 -4414 16437 -4380
rect 16471 -4414 16479 -4380
rect 16427 -4426 16479 -4414
rect 16144 -4492 16196 -4442
rect 17237 -4460 17289 -4338
rect 17319 -4312 17388 -4292
rect 17319 -4346 17333 -4312
rect 17367 -4346 17388 -4312
rect 17319 -4376 17388 -4346
rect 17418 -4305 17474 -4292
rect 17418 -4339 17430 -4305
rect 17464 -4339 17474 -4305
rect 17418 -4376 17474 -4339
rect 17504 -4376 17558 -4292
rect 17588 -4304 17666 -4292
rect 17588 -4338 17622 -4304
rect 17656 -4338 17666 -4304
rect 17588 -4376 17666 -4338
rect 17696 -4330 17750 -4292
rect 17696 -4364 17706 -4330
rect 17740 -4364 17750 -4330
rect 17696 -4376 17750 -4364
rect 17780 -4304 17914 -4292
rect 17780 -4338 17792 -4304
rect 17826 -4338 17870 -4304
rect 17904 -4338 17914 -4304
rect 17780 -4376 17914 -4338
rect 17319 -4460 17373 -4376
rect 17864 -4492 17914 -4376
rect 17944 -4312 18000 -4292
rect 17944 -4346 17954 -4312
rect 17988 -4346 18000 -4312
rect 17944 -4380 18000 -4346
rect 17944 -4414 17954 -4380
rect 17988 -4414 18000 -4380
rect 17944 -4448 18000 -4414
rect 18081 -4304 18133 -4292
rect 18081 -4338 18089 -4304
rect 18123 -4338 18133 -4304
rect 18081 -4372 18133 -4338
rect 18081 -4406 18089 -4372
rect 18123 -4406 18133 -4372
rect 18081 -4420 18133 -4406
rect 18163 -4304 18230 -4292
rect 18163 -4338 18186 -4304
rect 18220 -4338 18230 -4304
rect 18163 -4372 18230 -4338
rect 18163 -4406 18186 -4372
rect 18220 -4406 18230 -4372
rect 18163 -4420 18230 -4406
rect 17944 -4482 17954 -4448
rect 17988 -4482 18000 -4448
rect 17944 -4492 18000 -4482
rect 18178 -4440 18230 -4420
rect 18178 -4474 18186 -4440
rect 18220 -4474 18230 -4440
rect 18178 -4492 18230 -4474
rect 18260 -4340 18312 -4292
rect 18260 -4374 18270 -4340
rect 18304 -4374 18312 -4340
rect 18260 -4408 18312 -4374
rect 18260 -4442 18270 -4408
rect 18304 -4442 18312 -4408
rect 18377 -4312 18429 -4298
rect 18377 -4346 18385 -4312
rect 18419 -4346 18429 -4312
rect 18377 -4380 18429 -4346
rect 18377 -4414 18385 -4380
rect 18419 -4414 18429 -4380
rect 18377 -4426 18429 -4414
rect 18459 -4328 18513 -4298
rect 18459 -4362 18469 -4328
rect 18503 -4362 18513 -4328
rect 18459 -4426 18513 -4362
rect 18543 -4312 18595 -4298
rect 18543 -4346 18553 -4312
rect 18587 -4346 18595 -4312
rect 18543 -4380 18595 -4346
rect 18728 -4304 18780 -4292
rect 18728 -4338 18736 -4304
rect 18770 -4338 18780 -4304
rect 18728 -4376 18780 -4338
rect 18810 -4312 18872 -4292
rect 18810 -4346 18820 -4312
rect 18854 -4346 18872 -4312
rect 18810 -4376 18872 -4346
rect 18902 -4306 18971 -4292
rect 18902 -4340 18913 -4306
rect 18947 -4340 18971 -4306
rect 18902 -4376 18971 -4340
rect 19001 -4330 19111 -4292
rect 19001 -4364 19067 -4330
rect 19101 -4364 19111 -4330
rect 19001 -4376 19111 -4364
rect 19141 -4314 19208 -4292
rect 19141 -4348 19164 -4314
rect 19198 -4348 19208 -4314
rect 19141 -4376 19208 -4348
rect 19238 -4330 19290 -4292
rect 19238 -4364 19248 -4330
rect 19282 -4364 19290 -4330
rect 19238 -4376 19290 -4364
rect 19353 -4304 19405 -4292
rect 19353 -4338 19361 -4304
rect 19395 -4338 19405 -4304
rect 18543 -4414 18553 -4380
rect 18587 -4414 18595 -4380
rect 18543 -4426 18595 -4414
rect 18260 -4492 18312 -4442
rect 19353 -4460 19405 -4338
rect 19435 -4312 19504 -4292
rect 19435 -4346 19449 -4312
rect 19483 -4346 19504 -4312
rect 19435 -4376 19504 -4346
rect 19534 -4305 19590 -4292
rect 19534 -4339 19546 -4305
rect 19580 -4339 19590 -4305
rect 19534 -4376 19590 -4339
rect 19620 -4376 19674 -4292
rect 19704 -4304 19782 -4292
rect 19704 -4338 19738 -4304
rect 19772 -4338 19782 -4304
rect 19704 -4376 19782 -4338
rect 19812 -4330 19866 -4292
rect 19812 -4364 19822 -4330
rect 19856 -4364 19866 -4330
rect 19812 -4376 19866 -4364
rect 19896 -4304 20030 -4292
rect 19896 -4338 19908 -4304
rect 19942 -4338 19986 -4304
rect 20020 -4338 20030 -4304
rect 19896 -4376 20030 -4338
rect 19435 -4460 19489 -4376
rect 19980 -4492 20030 -4376
rect 20060 -4312 20116 -4292
rect 20060 -4346 20070 -4312
rect 20104 -4346 20116 -4312
rect 20060 -4380 20116 -4346
rect 20060 -4414 20070 -4380
rect 20104 -4414 20116 -4380
rect 20060 -4448 20116 -4414
rect 20197 -4304 20249 -4292
rect 20197 -4338 20205 -4304
rect 20239 -4338 20249 -4304
rect 20197 -4372 20249 -4338
rect 20197 -4406 20205 -4372
rect 20239 -4406 20249 -4372
rect 20197 -4420 20249 -4406
rect 20279 -4304 20346 -4292
rect 20279 -4338 20302 -4304
rect 20336 -4338 20346 -4304
rect 20279 -4372 20346 -4338
rect 20279 -4406 20302 -4372
rect 20336 -4406 20346 -4372
rect 20279 -4420 20346 -4406
rect 20060 -4482 20070 -4448
rect 20104 -4482 20116 -4448
rect 20060 -4492 20116 -4482
rect 20294 -4440 20346 -4420
rect 20294 -4474 20302 -4440
rect 20336 -4474 20346 -4440
rect 20294 -4492 20346 -4474
rect 20376 -4340 20428 -4292
rect 20376 -4374 20386 -4340
rect 20420 -4374 20428 -4340
rect 20376 -4408 20428 -4374
rect 20376 -4442 20386 -4408
rect 20420 -4442 20428 -4408
rect 20493 -4312 20545 -4298
rect 20493 -4346 20501 -4312
rect 20535 -4346 20545 -4312
rect 20493 -4380 20545 -4346
rect 20493 -4414 20501 -4380
rect 20535 -4414 20545 -4380
rect 20493 -4426 20545 -4414
rect 20575 -4328 20629 -4298
rect 20575 -4362 20585 -4328
rect 20619 -4362 20629 -4328
rect 20575 -4426 20629 -4362
rect 20659 -4312 20711 -4298
rect 20659 -4346 20669 -4312
rect 20703 -4346 20711 -4312
rect 20659 -4380 20711 -4346
rect 20844 -4304 20896 -4292
rect 20844 -4338 20852 -4304
rect 20886 -4338 20896 -4304
rect 20844 -4376 20896 -4338
rect 20926 -4312 20988 -4292
rect 20926 -4346 20936 -4312
rect 20970 -4346 20988 -4312
rect 20926 -4376 20988 -4346
rect 21018 -4306 21087 -4292
rect 21018 -4340 21029 -4306
rect 21063 -4340 21087 -4306
rect 21018 -4376 21087 -4340
rect 21117 -4330 21227 -4292
rect 21117 -4364 21183 -4330
rect 21217 -4364 21227 -4330
rect 21117 -4376 21227 -4364
rect 21257 -4314 21324 -4292
rect 21257 -4348 21280 -4314
rect 21314 -4348 21324 -4314
rect 21257 -4376 21324 -4348
rect 21354 -4330 21406 -4292
rect 21354 -4364 21364 -4330
rect 21398 -4364 21406 -4330
rect 21354 -4376 21406 -4364
rect 21469 -4304 21521 -4292
rect 21469 -4338 21477 -4304
rect 21511 -4338 21521 -4304
rect 20659 -4414 20669 -4380
rect 20703 -4414 20711 -4380
rect 20659 -4426 20711 -4414
rect 20376 -4492 20428 -4442
rect 21469 -4460 21521 -4338
rect 21551 -4312 21620 -4292
rect 21551 -4346 21565 -4312
rect 21599 -4346 21620 -4312
rect 21551 -4376 21620 -4346
rect 21650 -4305 21706 -4292
rect 21650 -4339 21662 -4305
rect 21696 -4339 21706 -4305
rect 21650 -4376 21706 -4339
rect 21736 -4376 21790 -4292
rect 21820 -4304 21898 -4292
rect 21820 -4338 21854 -4304
rect 21888 -4338 21898 -4304
rect 21820 -4376 21898 -4338
rect 21928 -4330 21982 -4292
rect 21928 -4364 21938 -4330
rect 21972 -4364 21982 -4330
rect 21928 -4376 21982 -4364
rect 22012 -4304 22146 -4292
rect 22012 -4338 22024 -4304
rect 22058 -4338 22102 -4304
rect 22136 -4338 22146 -4304
rect 22012 -4376 22146 -4338
rect 21551 -4460 21605 -4376
rect 22096 -4492 22146 -4376
rect 22176 -4312 22232 -4292
rect 22176 -4346 22186 -4312
rect 22220 -4346 22232 -4312
rect 22176 -4380 22232 -4346
rect 22176 -4414 22186 -4380
rect 22220 -4414 22232 -4380
rect 22176 -4448 22232 -4414
rect 22313 -4304 22365 -4292
rect 22313 -4338 22321 -4304
rect 22355 -4338 22365 -4304
rect 22313 -4372 22365 -4338
rect 22313 -4406 22321 -4372
rect 22355 -4406 22365 -4372
rect 22313 -4420 22365 -4406
rect 22395 -4304 22462 -4292
rect 22395 -4338 22418 -4304
rect 22452 -4338 22462 -4304
rect 22395 -4372 22462 -4338
rect 22395 -4406 22418 -4372
rect 22452 -4406 22462 -4372
rect 22395 -4420 22462 -4406
rect 22176 -4482 22186 -4448
rect 22220 -4482 22232 -4448
rect 22176 -4492 22232 -4482
rect 22410 -4440 22462 -4420
rect 22410 -4474 22418 -4440
rect 22452 -4474 22462 -4440
rect 22410 -4492 22462 -4474
rect 22492 -4340 22544 -4292
rect 22492 -4374 22502 -4340
rect 22536 -4374 22544 -4340
rect 22492 -4408 22544 -4374
rect 22492 -4442 22502 -4408
rect 22536 -4442 22544 -4408
rect 22609 -4312 22661 -4298
rect 22609 -4346 22617 -4312
rect 22651 -4346 22661 -4312
rect 22609 -4380 22661 -4346
rect 22609 -4414 22617 -4380
rect 22651 -4414 22661 -4380
rect 22609 -4426 22661 -4414
rect 22691 -4328 22745 -4298
rect 22691 -4362 22701 -4328
rect 22735 -4362 22745 -4328
rect 22691 -4426 22745 -4362
rect 22775 -4312 22827 -4298
rect 22775 -4346 22785 -4312
rect 22819 -4346 22827 -4312
rect 22775 -4380 22827 -4346
rect 22960 -4304 23012 -4292
rect 22960 -4338 22968 -4304
rect 23002 -4338 23012 -4304
rect 22960 -4376 23012 -4338
rect 23042 -4312 23104 -4292
rect 23042 -4346 23052 -4312
rect 23086 -4346 23104 -4312
rect 23042 -4376 23104 -4346
rect 23134 -4306 23203 -4292
rect 23134 -4340 23145 -4306
rect 23179 -4340 23203 -4306
rect 23134 -4376 23203 -4340
rect 23233 -4330 23343 -4292
rect 23233 -4364 23299 -4330
rect 23333 -4364 23343 -4330
rect 23233 -4376 23343 -4364
rect 23373 -4314 23440 -4292
rect 23373 -4348 23396 -4314
rect 23430 -4348 23440 -4314
rect 23373 -4376 23440 -4348
rect 23470 -4330 23522 -4292
rect 23470 -4364 23480 -4330
rect 23514 -4364 23522 -4330
rect 23470 -4376 23522 -4364
rect 23585 -4304 23637 -4292
rect 23585 -4338 23593 -4304
rect 23627 -4338 23637 -4304
rect 22775 -4414 22785 -4380
rect 22819 -4414 22827 -4380
rect 22775 -4426 22827 -4414
rect 22492 -4492 22544 -4442
rect 23585 -4460 23637 -4338
rect 23667 -4312 23736 -4292
rect 23667 -4346 23681 -4312
rect 23715 -4346 23736 -4312
rect 23667 -4376 23736 -4346
rect 23766 -4305 23822 -4292
rect 23766 -4339 23778 -4305
rect 23812 -4339 23822 -4305
rect 23766 -4376 23822 -4339
rect 23852 -4376 23906 -4292
rect 23936 -4304 24014 -4292
rect 23936 -4338 23970 -4304
rect 24004 -4338 24014 -4304
rect 23936 -4376 24014 -4338
rect 24044 -4330 24098 -4292
rect 24044 -4364 24054 -4330
rect 24088 -4364 24098 -4330
rect 24044 -4376 24098 -4364
rect 24128 -4304 24262 -4292
rect 24128 -4338 24140 -4304
rect 24174 -4338 24218 -4304
rect 24252 -4338 24262 -4304
rect 24128 -4376 24262 -4338
rect 23667 -4460 23721 -4376
rect 24212 -4492 24262 -4376
rect 24292 -4312 24348 -4292
rect 24292 -4346 24302 -4312
rect 24336 -4346 24348 -4312
rect 24292 -4380 24348 -4346
rect 24292 -4414 24302 -4380
rect 24336 -4414 24348 -4380
rect 24292 -4448 24348 -4414
rect 24429 -4304 24481 -4292
rect 24429 -4338 24437 -4304
rect 24471 -4338 24481 -4304
rect 24429 -4372 24481 -4338
rect 24429 -4406 24437 -4372
rect 24471 -4406 24481 -4372
rect 24429 -4420 24481 -4406
rect 24511 -4304 24578 -4292
rect 24511 -4338 24534 -4304
rect 24568 -4338 24578 -4304
rect 24511 -4372 24578 -4338
rect 24511 -4406 24534 -4372
rect 24568 -4406 24578 -4372
rect 24511 -4420 24578 -4406
rect 24292 -4482 24302 -4448
rect 24336 -4482 24348 -4448
rect 24292 -4492 24348 -4482
rect 24526 -4440 24578 -4420
rect 24526 -4474 24534 -4440
rect 24568 -4474 24578 -4440
rect 24526 -4492 24578 -4474
rect 24608 -4340 24660 -4292
rect 24608 -4374 24618 -4340
rect 24652 -4374 24660 -4340
rect 24608 -4408 24660 -4374
rect 24608 -4442 24618 -4408
rect 24652 -4442 24660 -4408
rect 24725 -4312 24777 -4298
rect 24725 -4346 24733 -4312
rect 24767 -4346 24777 -4312
rect 24725 -4380 24777 -4346
rect 24725 -4414 24733 -4380
rect 24767 -4414 24777 -4380
rect 24725 -4426 24777 -4414
rect 24807 -4328 24861 -4298
rect 24807 -4362 24817 -4328
rect 24851 -4362 24861 -4328
rect 24807 -4426 24861 -4362
rect 24891 -4312 24943 -4298
rect 24891 -4346 24901 -4312
rect 24935 -4346 24943 -4312
rect 24891 -4380 24943 -4346
rect 25076 -4304 25128 -4292
rect 25076 -4338 25084 -4304
rect 25118 -4338 25128 -4304
rect 25076 -4376 25128 -4338
rect 25158 -4312 25220 -4292
rect 25158 -4346 25168 -4312
rect 25202 -4346 25220 -4312
rect 25158 -4376 25220 -4346
rect 25250 -4306 25319 -4292
rect 25250 -4340 25261 -4306
rect 25295 -4340 25319 -4306
rect 25250 -4376 25319 -4340
rect 25349 -4330 25459 -4292
rect 25349 -4364 25415 -4330
rect 25449 -4364 25459 -4330
rect 25349 -4376 25459 -4364
rect 25489 -4314 25556 -4292
rect 25489 -4348 25512 -4314
rect 25546 -4348 25556 -4314
rect 25489 -4376 25556 -4348
rect 25586 -4330 25638 -4292
rect 25586 -4364 25596 -4330
rect 25630 -4364 25638 -4330
rect 25586 -4376 25638 -4364
rect 25701 -4304 25753 -4292
rect 25701 -4338 25709 -4304
rect 25743 -4338 25753 -4304
rect 24891 -4414 24901 -4380
rect 24935 -4414 24943 -4380
rect 24891 -4426 24943 -4414
rect 24608 -4492 24660 -4442
rect 25701 -4460 25753 -4338
rect 25783 -4312 25852 -4292
rect 25783 -4346 25797 -4312
rect 25831 -4346 25852 -4312
rect 25783 -4376 25852 -4346
rect 25882 -4305 25938 -4292
rect 25882 -4339 25894 -4305
rect 25928 -4339 25938 -4305
rect 25882 -4376 25938 -4339
rect 25968 -4376 26022 -4292
rect 26052 -4304 26130 -4292
rect 26052 -4338 26086 -4304
rect 26120 -4338 26130 -4304
rect 26052 -4376 26130 -4338
rect 26160 -4330 26214 -4292
rect 26160 -4364 26170 -4330
rect 26204 -4364 26214 -4330
rect 26160 -4376 26214 -4364
rect 26244 -4304 26378 -4292
rect 26244 -4338 26256 -4304
rect 26290 -4338 26334 -4304
rect 26368 -4338 26378 -4304
rect 26244 -4376 26378 -4338
rect 25783 -4460 25837 -4376
rect 26328 -4492 26378 -4376
rect 26408 -4312 26464 -4292
rect 26408 -4346 26418 -4312
rect 26452 -4346 26464 -4312
rect 26408 -4380 26464 -4346
rect 26408 -4414 26418 -4380
rect 26452 -4414 26464 -4380
rect 26408 -4448 26464 -4414
rect 26545 -4304 26597 -4292
rect 26545 -4338 26553 -4304
rect 26587 -4338 26597 -4304
rect 26545 -4372 26597 -4338
rect 26545 -4406 26553 -4372
rect 26587 -4406 26597 -4372
rect 26545 -4420 26597 -4406
rect 26627 -4304 26694 -4292
rect 26627 -4338 26650 -4304
rect 26684 -4338 26694 -4304
rect 26627 -4372 26694 -4338
rect 26627 -4406 26650 -4372
rect 26684 -4406 26694 -4372
rect 26627 -4420 26694 -4406
rect 26408 -4482 26418 -4448
rect 26452 -4482 26464 -4448
rect 26408 -4492 26464 -4482
rect 26642 -4440 26694 -4420
rect 26642 -4474 26650 -4440
rect 26684 -4474 26694 -4440
rect 26642 -4492 26694 -4474
rect 26724 -4340 26776 -4292
rect 26724 -4374 26734 -4340
rect 26768 -4374 26776 -4340
rect 26724 -4408 26776 -4374
rect 26724 -4442 26734 -4408
rect 26768 -4442 26776 -4408
rect 26841 -4312 26893 -4298
rect 26841 -4346 26849 -4312
rect 26883 -4346 26893 -4312
rect 26841 -4380 26893 -4346
rect 26841 -4414 26849 -4380
rect 26883 -4414 26893 -4380
rect 26841 -4426 26893 -4414
rect 26923 -4328 26977 -4298
rect 26923 -4362 26933 -4328
rect 26967 -4362 26977 -4328
rect 26923 -4426 26977 -4362
rect 27007 -4312 27059 -4298
rect 27007 -4346 27017 -4312
rect 27051 -4346 27059 -4312
rect 27007 -4380 27059 -4346
rect 27192 -4304 27244 -4292
rect 27192 -4338 27200 -4304
rect 27234 -4338 27244 -4304
rect 27192 -4376 27244 -4338
rect 27274 -4312 27336 -4292
rect 27274 -4346 27284 -4312
rect 27318 -4346 27336 -4312
rect 27274 -4376 27336 -4346
rect 27366 -4306 27435 -4292
rect 27366 -4340 27377 -4306
rect 27411 -4340 27435 -4306
rect 27366 -4376 27435 -4340
rect 27465 -4330 27575 -4292
rect 27465 -4364 27531 -4330
rect 27565 -4364 27575 -4330
rect 27465 -4376 27575 -4364
rect 27605 -4314 27672 -4292
rect 27605 -4348 27628 -4314
rect 27662 -4348 27672 -4314
rect 27605 -4376 27672 -4348
rect 27702 -4330 27754 -4292
rect 27702 -4364 27712 -4330
rect 27746 -4364 27754 -4330
rect 27702 -4376 27754 -4364
rect 27817 -4304 27869 -4292
rect 27817 -4338 27825 -4304
rect 27859 -4338 27869 -4304
rect 27007 -4414 27017 -4380
rect 27051 -4414 27059 -4380
rect 27007 -4426 27059 -4414
rect 26724 -4492 26776 -4442
rect 27817 -4460 27869 -4338
rect 27899 -4312 27968 -4292
rect 27899 -4346 27913 -4312
rect 27947 -4346 27968 -4312
rect 27899 -4376 27968 -4346
rect 27998 -4305 28054 -4292
rect 27998 -4339 28010 -4305
rect 28044 -4339 28054 -4305
rect 27998 -4376 28054 -4339
rect 28084 -4376 28138 -4292
rect 28168 -4304 28246 -4292
rect 28168 -4338 28202 -4304
rect 28236 -4338 28246 -4304
rect 28168 -4376 28246 -4338
rect 28276 -4330 28330 -4292
rect 28276 -4364 28286 -4330
rect 28320 -4364 28330 -4330
rect 28276 -4376 28330 -4364
rect 28360 -4304 28494 -4292
rect 28360 -4338 28372 -4304
rect 28406 -4338 28450 -4304
rect 28484 -4338 28494 -4304
rect 28360 -4376 28494 -4338
rect 27899 -4460 27953 -4376
rect 28444 -4492 28494 -4376
rect 28524 -4312 28580 -4292
rect 28524 -4346 28534 -4312
rect 28568 -4346 28580 -4312
rect 28524 -4380 28580 -4346
rect 28524 -4414 28534 -4380
rect 28568 -4414 28580 -4380
rect 28524 -4448 28580 -4414
rect 28661 -4304 28713 -4292
rect 28661 -4338 28669 -4304
rect 28703 -4338 28713 -4304
rect 28661 -4372 28713 -4338
rect 28661 -4406 28669 -4372
rect 28703 -4406 28713 -4372
rect 28661 -4420 28713 -4406
rect 28743 -4304 28810 -4292
rect 28743 -4338 28766 -4304
rect 28800 -4338 28810 -4304
rect 28743 -4372 28810 -4338
rect 28743 -4406 28766 -4372
rect 28800 -4406 28810 -4372
rect 28743 -4420 28810 -4406
rect 28524 -4482 28534 -4448
rect 28568 -4482 28580 -4448
rect 28524 -4492 28580 -4482
rect 28758 -4440 28810 -4420
rect 28758 -4474 28766 -4440
rect 28800 -4474 28810 -4440
rect 28758 -4492 28810 -4474
rect 28840 -4340 28892 -4292
rect 28840 -4374 28850 -4340
rect 28884 -4374 28892 -4340
rect 28840 -4408 28892 -4374
rect 28840 -4442 28850 -4408
rect 28884 -4442 28892 -4408
rect 28957 -4312 29009 -4298
rect 28957 -4346 28965 -4312
rect 28999 -4346 29009 -4312
rect 28957 -4380 29009 -4346
rect 28957 -4414 28965 -4380
rect 28999 -4414 29009 -4380
rect 28957 -4426 29009 -4414
rect 29039 -4328 29093 -4298
rect 29039 -4362 29049 -4328
rect 29083 -4362 29093 -4328
rect 29039 -4426 29093 -4362
rect 29123 -4312 29175 -4298
rect 29123 -4346 29133 -4312
rect 29167 -4346 29175 -4312
rect 29123 -4380 29175 -4346
rect 29308 -4304 29360 -4292
rect 29308 -4338 29316 -4304
rect 29350 -4338 29360 -4304
rect 29308 -4376 29360 -4338
rect 29390 -4312 29452 -4292
rect 29390 -4346 29400 -4312
rect 29434 -4346 29452 -4312
rect 29390 -4376 29452 -4346
rect 29482 -4306 29551 -4292
rect 29482 -4340 29493 -4306
rect 29527 -4340 29551 -4306
rect 29482 -4376 29551 -4340
rect 29581 -4330 29691 -4292
rect 29581 -4364 29647 -4330
rect 29681 -4364 29691 -4330
rect 29581 -4376 29691 -4364
rect 29721 -4314 29788 -4292
rect 29721 -4348 29744 -4314
rect 29778 -4348 29788 -4314
rect 29721 -4376 29788 -4348
rect 29818 -4330 29870 -4292
rect 29818 -4364 29828 -4330
rect 29862 -4364 29870 -4330
rect 29818 -4376 29870 -4364
rect 29933 -4304 29985 -4292
rect 29933 -4338 29941 -4304
rect 29975 -4338 29985 -4304
rect 29123 -4414 29133 -4380
rect 29167 -4414 29175 -4380
rect 29123 -4426 29175 -4414
rect 28840 -4492 28892 -4442
rect 29933 -4460 29985 -4338
rect 30015 -4312 30084 -4292
rect 30015 -4346 30029 -4312
rect 30063 -4346 30084 -4312
rect 30015 -4376 30084 -4346
rect 30114 -4305 30170 -4292
rect 30114 -4339 30126 -4305
rect 30160 -4339 30170 -4305
rect 30114 -4376 30170 -4339
rect 30200 -4376 30254 -4292
rect 30284 -4304 30362 -4292
rect 30284 -4338 30318 -4304
rect 30352 -4338 30362 -4304
rect 30284 -4376 30362 -4338
rect 30392 -4330 30446 -4292
rect 30392 -4364 30402 -4330
rect 30436 -4364 30446 -4330
rect 30392 -4376 30446 -4364
rect 30476 -4304 30610 -4292
rect 30476 -4338 30488 -4304
rect 30522 -4338 30566 -4304
rect 30600 -4338 30610 -4304
rect 30476 -4376 30610 -4338
rect 30015 -4460 30069 -4376
rect 30560 -4492 30610 -4376
rect 30640 -4312 30696 -4292
rect 30640 -4346 30650 -4312
rect 30684 -4346 30696 -4312
rect 30640 -4380 30696 -4346
rect 30640 -4414 30650 -4380
rect 30684 -4414 30696 -4380
rect 30640 -4448 30696 -4414
rect 30777 -4304 30829 -4292
rect 30777 -4338 30785 -4304
rect 30819 -4338 30829 -4304
rect 30777 -4372 30829 -4338
rect 30777 -4406 30785 -4372
rect 30819 -4406 30829 -4372
rect 30777 -4420 30829 -4406
rect 30859 -4304 30926 -4292
rect 30859 -4338 30882 -4304
rect 30916 -4338 30926 -4304
rect 30859 -4372 30926 -4338
rect 30859 -4406 30882 -4372
rect 30916 -4406 30926 -4372
rect 30859 -4420 30926 -4406
rect 30640 -4482 30650 -4448
rect 30684 -4482 30696 -4448
rect 30640 -4492 30696 -4482
rect 30874 -4440 30926 -4420
rect 30874 -4474 30882 -4440
rect 30916 -4474 30926 -4440
rect 30874 -4492 30926 -4474
rect 30956 -4340 31008 -4292
rect 30956 -4374 30966 -4340
rect 31000 -4374 31008 -4340
rect 30956 -4408 31008 -4374
rect 30956 -4442 30966 -4408
rect 31000 -4442 31008 -4408
rect 31073 -4312 31125 -4298
rect 31073 -4346 31081 -4312
rect 31115 -4346 31125 -4312
rect 31073 -4380 31125 -4346
rect 31073 -4414 31081 -4380
rect 31115 -4414 31125 -4380
rect 31073 -4426 31125 -4414
rect 31155 -4328 31209 -4298
rect 31155 -4362 31165 -4328
rect 31199 -4362 31209 -4328
rect 31155 -4426 31209 -4362
rect 31239 -4312 31291 -4298
rect 31239 -4346 31249 -4312
rect 31283 -4346 31291 -4312
rect 31239 -4380 31291 -4346
rect 31424 -4304 31476 -4292
rect 31424 -4338 31432 -4304
rect 31466 -4338 31476 -4304
rect 31424 -4376 31476 -4338
rect 31506 -4312 31568 -4292
rect 31506 -4346 31516 -4312
rect 31550 -4346 31568 -4312
rect 31506 -4376 31568 -4346
rect 31598 -4306 31667 -4292
rect 31598 -4340 31609 -4306
rect 31643 -4340 31667 -4306
rect 31598 -4376 31667 -4340
rect 31697 -4330 31807 -4292
rect 31697 -4364 31763 -4330
rect 31797 -4364 31807 -4330
rect 31697 -4376 31807 -4364
rect 31837 -4314 31904 -4292
rect 31837 -4348 31860 -4314
rect 31894 -4348 31904 -4314
rect 31837 -4376 31904 -4348
rect 31934 -4330 31986 -4292
rect 31934 -4364 31944 -4330
rect 31978 -4364 31986 -4330
rect 31934 -4376 31986 -4364
rect 32049 -4304 32101 -4292
rect 32049 -4338 32057 -4304
rect 32091 -4338 32101 -4304
rect 31239 -4414 31249 -4380
rect 31283 -4414 31291 -4380
rect 31239 -4426 31291 -4414
rect 30956 -4492 31008 -4442
rect 32049 -4460 32101 -4338
rect 32131 -4312 32200 -4292
rect 32131 -4346 32145 -4312
rect 32179 -4346 32200 -4312
rect 32131 -4376 32200 -4346
rect 32230 -4305 32286 -4292
rect 32230 -4339 32242 -4305
rect 32276 -4339 32286 -4305
rect 32230 -4376 32286 -4339
rect 32316 -4376 32370 -4292
rect 32400 -4304 32478 -4292
rect 32400 -4338 32434 -4304
rect 32468 -4338 32478 -4304
rect 32400 -4376 32478 -4338
rect 32508 -4330 32562 -4292
rect 32508 -4364 32518 -4330
rect 32552 -4364 32562 -4330
rect 32508 -4376 32562 -4364
rect 32592 -4304 32726 -4292
rect 32592 -4338 32604 -4304
rect 32638 -4338 32682 -4304
rect 32716 -4338 32726 -4304
rect 32592 -4376 32726 -4338
rect 32131 -4460 32185 -4376
rect 32676 -4492 32726 -4376
rect 32756 -4312 32812 -4292
rect 32756 -4346 32766 -4312
rect 32800 -4346 32812 -4312
rect 32756 -4380 32812 -4346
rect 32756 -4414 32766 -4380
rect 32800 -4414 32812 -4380
rect 32756 -4448 32812 -4414
rect 32893 -4304 32945 -4292
rect 32893 -4338 32901 -4304
rect 32935 -4338 32945 -4304
rect 32893 -4372 32945 -4338
rect 32893 -4406 32901 -4372
rect 32935 -4406 32945 -4372
rect 32893 -4420 32945 -4406
rect 32975 -4304 33042 -4292
rect 32975 -4338 32998 -4304
rect 33032 -4338 33042 -4304
rect 32975 -4372 33042 -4338
rect 32975 -4406 32998 -4372
rect 33032 -4406 33042 -4372
rect 32975 -4420 33042 -4406
rect 32756 -4482 32766 -4448
rect 32800 -4482 32812 -4448
rect 32756 -4492 32812 -4482
rect 32990 -4440 33042 -4420
rect 32990 -4474 32998 -4440
rect 33032 -4474 33042 -4440
rect 32990 -4492 33042 -4474
rect 33072 -4340 33124 -4292
rect 33072 -4374 33082 -4340
rect 33116 -4374 33124 -4340
rect 33072 -4408 33124 -4374
rect 33072 -4442 33082 -4408
rect 33116 -4442 33124 -4408
rect 33072 -4492 33124 -4442
rect 9375 -7683 9433 -7675
rect 9375 -7719 9388 -7683
rect 9422 -7719 9433 -7683
rect 9375 -7757 9433 -7719
rect 9375 -7793 9387 -7757
rect 9421 -7793 9433 -7757
rect 9375 -7830 9433 -7793
rect 9375 -7866 9387 -7830
rect 9421 -7866 9433 -7830
rect 9375 -7875 9433 -7866
rect 9633 -7687 9691 -7675
rect 9633 -7723 9645 -7687
rect 9679 -7723 9691 -7687
rect 9633 -7757 9691 -7723
rect 9633 -7793 9645 -7757
rect 9679 -7793 9691 -7757
rect 9633 -7830 9691 -7793
rect 9633 -7866 9644 -7830
rect 9678 -7866 9691 -7830
rect 9633 -7875 9691 -7866
rect 10035 -7683 10093 -7675
rect 10035 -7719 10048 -7683
rect 10082 -7719 10093 -7683
rect 10035 -7757 10093 -7719
rect 10035 -7793 10047 -7757
rect 10081 -7793 10093 -7757
rect 10035 -7830 10093 -7793
rect 10035 -7866 10047 -7830
rect 10081 -7866 10093 -7830
rect 10035 -7875 10093 -7866
rect 10293 -7687 10351 -7675
rect 10293 -7723 10305 -7687
rect 10339 -7723 10351 -7687
rect 10293 -7757 10351 -7723
rect 10293 -7793 10305 -7757
rect 10339 -7793 10351 -7757
rect 10293 -7830 10351 -7793
rect 10293 -7866 10304 -7830
rect 10338 -7866 10351 -7830
rect 10293 -7875 10351 -7866
rect 10505 -7683 10563 -7675
rect 10505 -7719 10518 -7683
rect 10552 -7719 10563 -7683
rect 10505 -7757 10563 -7719
rect 10505 -7793 10517 -7757
rect 10551 -7793 10563 -7757
rect 10505 -7830 10563 -7793
rect 10505 -7866 10517 -7830
rect 10551 -7866 10563 -7830
rect 10505 -7875 10563 -7866
rect 10763 -7687 10821 -7675
rect 10763 -7723 10775 -7687
rect 10809 -7723 10821 -7687
rect 10763 -7757 10821 -7723
rect 10763 -7793 10775 -7757
rect 10809 -7793 10821 -7757
rect 10763 -7830 10821 -7793
rect 10763 -7866 10774 -7830
rect 10808 -7866 10821 -7830
rect 10763 -7875 10821 -7866
rect 11108 -7687 11166 -7676
rect 11108 -7723 11120 -7687
rect 11154 -7723 11166 -7687
rect 11108 -7758 11166 -7723
rect 11108 -7794 11120 -7758
rect 11154 -7794 11166 -7758
rect 11108 -7829 11166 -7794
rect 11108 -7865 11120 -7829
rect 11154 -7865 11166 -7829
rect 11108 -7876 11166 -7865
rect 11366 -7687 11424 -7676
rect 11366 -7723 11378 -7687
rect 11412 -7723 11424 -7687
rect 11366 -7758 11424 -7723
rect 11366 -7794 11378 -7758
rect 11412 -7794 11424 -7758
rect 11366 -7829 11424 -7794
rect 11366 -7865 11378 -7829
rect 11412 -7865 11424 -7829
rect 11366 -7876 11424 -7865
rect 11624 -7687 11682 -7676
rect 11624 -7723 11636 -7687
rect 11670 -7723 11682 -7687
rect 11624 -7758 11682 -7723
rect 11624 -7794 11636 -7758
rect 11670 -7794 11682 -7758
rect 11624 -7829 11682 -7794
rect 11624 -7865 11636 -7829
rect 11670 -7865 11682 -7829
rect 11624 -7876 11682 -7865
rect 11882 -7687 11940 -7676
rect 11882 -7723 11894 -7687
rect 11928 -7723 11940 -7687
rect 11882 -7758 11940 -7723
rect 11882 -7794 11894 -7758
rect 11928 -7794 11940 -7758
rect 11882 -7829 11940 -7794
rect 11882 -7865 11894 -7829
rect 11928 -7865 11940 -7829
rect 11882 -7876 11940 -7865
rect 12140 -7687 12198 -7676
rect 12140 -7723 12152 -7687
rect 12186 -7723 12198 -7687
rect 12140 -7758 12198 -7723
rect 12140 -7794 12152 -7758
rect 12186 -7794 12198 -7758
rect 12140 -7829 12198 -7794
rect 12140 -7865 12152 -7829
rect 12186 -7865 12198 -7829
rect 12140 -7876 12198 -7865
rect 12398 -7687 12456 -7676
rect 12398 -7723 12410 -7687
rect 12444 -7723 12456 -7687
rect 12398 -7758 12456 -7723
rect 12398 -7794 12410 -7758
rect 12444 -7794 12456 -7758
rect 12398 -7829 12456 -7794
rect 12398 -7865 12410 -7829
rect 12444 -7865 12456 -7829
rect 12398 -7876 12456 -7865
rect 12923 -7687 12981 -7676
rect 12923 -7723 12935 -7687
rect 12969 -7723 12981 -7687
rect 12923 -7758 12981 -7723
rect 12923 -7794 12935 -7758
rect 12969 -7794 12981 -7758
rect 12923 -7829 12981 -7794
rect 12923 -7865 12935 -7829
rect 12969 -7865 12981 -7829
rect 12923 -7876 12981 -7865
rect 13181 -7687 13239 -7676
rect 13181 -7723 13193 -7687
rect 13227 -7723 13239 -7687
rect 13181 -7758 13239 -7723
rect 13181 -7794 13193 -7758
rect 13227 -7794 13239 -7758
rect 13181 -7829 13239 -7794
rect 13181 -7865 13193 -7829
rect 13227 -7865 13239 -7829
rect 13181 -7876 13239 -7865
rect 13439 -7687 13497 -7676
rect 13439 -7723 13451 -7687
rect 13485 -7723 13497 -7687
rect 13439 -7758 13497 -7723
rect 13439 -7794 13451 -7758
rect 13485 -7794 13497 -7758
rect 13439 -7829 13497 -7794
rect 13439 -7865 13451 -7829
rect 13485 -7865 13497 -7829
rect 13439 -7876 13497 -7865
rect 13697 -7687 13755 -7676
rect 13697 -7723 13709 -7687
rect 13743 -7723 13755 -7687
rect 13697 -7758 13755 -7723
rect 13697 -7794 13709 -7758
rect 13743 -7794 13755 -7758
rect 13697 -7829 13755 -7794
rect 13697 -7865 13709 -7829
rect 13743 -7865 13755 -7829
rect 13697 -7876 13755 -7865
rect 13955 -7687 14013 -7676
rect 13955 -7723 13967 -7687
rect 14001 -7723 14013 -7687
rect 13955 -7758 14013 -7723
rect 13955 -7794 13967 -7758
rect 14001 -7794 14013 -7758
rect 13955 -7829 14013 -7794
rect 13955 -7865 13967 -7829
rect 14001 -7865 14013 -7829
rect 13955 -7876 14013 -7865
rect 14213 -7687 14271 -7676
rect 14213 -7723 14225 -7687
rect 14259 -7723 14271 -7687
rect 14213 -7758 14271 -7723
rect 14213 -7794 14225 -7758
rect 14259 -7794 14271 -7758
rect 14213 -7829 14271 -7794
rect 14213 -7865 14225 -7829
rect 14259 -7865 14271 -7829
rect 14213 -7876 14271 -7865
rect 14729 -7687 14787 -7676
rect 14729 -7723 14741 -7687
rect 14775 -7723 14787 -7687
rect 14729 -7758 14787 -7723
rect 14729 -7794 14741 -7758
rect 14775 -7794 14787 -7758
rect 14729 -7829 14787 -7794
rect 14729 -7865 14741 -7829
rect 14775 -7865 14787 -7829
rect 14729 -7876 14787 -7865
rect 14987 -7687 15045 -7676
rect 14987 -7723 14999 -7687
rect 15033 -7723 15045 -7687
rect 14987 -7758 15045 -7723
rect 14987 -7794 14999 -7758
rect 15033 -7794 15045 -7758
rect 14987 -7829 15045 -7794
rect 14987 -7865 14999 -7829
rect 15033 -7865 15045 -7829
rect 14987 -7876 15045 -7865
rect 15245 -7687 15303 -7676
rect 15245 -7723 15257 -7687
rect 15291 -7723 15303 -7687
rect 15245 -7758 15303 -7723
rect 15245 -7794 15257 -7758
rect 15291 -7794 15303 -7758
rect 15245 -7829 15303 -7794
rect 15245 -7865 15257 -7829
rect 15291 -7865 15303 -7829
rect 15245 -7876 15303 -7865
rect 15503 -7687 15561 -7676
rect 15503 -7723 15515 -7687
rect 15549 -7723 15561 -7687
rect 15503 -7758 15561 -7723
rect 15503 -7794 15515 -7758
rect 15549 -7794 15561 -7758
rect 15503 -7829 15561 -7794
rect 15503 -7865 15515 -7829
rect 15549 -7865 15561 -7829
rect 15503 -7876 15561 -7865
rect 15761 -7687 15819 -7676
rect 15761 -7723 15773 -7687
rect 15807 -7723 15819 -7687
rect 15761 -7758 15819 -7723
rect 15761 -7794 15773 -7758
rect 15807 -7794 15819 -7758
rect 15761 -7829 15819 -7794
rect 15761 -7865 15773 -7829
rect 15807 -7865 15819 -7829
rect 15761 -7876 15819 -7865
rect 16019 -7687 16077 -7676
rect 16019 -7723 16031 -7687
rect 16065 -7723 16077 -7687
rect 16019 -7758 16077 -7723
rect 16019 -7794 16031 -7758
rect 16065 -7794 16077 -7758
rect 16019 -7829 16077 -7794
rect 16019 -7865 16031 -7829
rect 16065 -7865 16077 -7829
rect 16019 -7876 16077 -7865
rect 9310 -8687 9384 -8649
rect 9310 -8723 9330 -8687
rect 9368 -8723 9384 -8687
rect 9310 -8759 9384 -8723
rect 9500 -8685 9574 -8649
rect 9500 -8721 9516 -8685
rect 9554 -8721 9574 -8685
rect 9500 -8759 9574 -8721
rect 9679 -8687 9737 -8649
rect 9679 -8721 9691 -8687
rect 9725 -8721 9737 -8687
rect 9679 -8759 9737 -8721
rect 10537 -8687 10595 -8649
rect 10537 -8721 10549 -8687
rect 10583 -8721 10595 -8687
rect 10537 -8759 10595 -8721
rect 10696 -8687 10770 -8649
rect 10696 -8723 10716 -8687
rect 10754 -8723 10770 -8687
rect 10696 -8759 10770 -8723
rect 10886 -8685 10960 -8649
rect 10886 -8721 10902 -8685
rect 10940 -8721 10960 -8685
rect 10886 -8759 10960 -8721
rect 11066 -8687 11140 -8649
rect 11066 -8723 11086 -8687
rect 11124 -8723 11140 -8687
rect 11066 -8759 11140 -8723
rect 11256 -8685 11330 -8649
rect 11256 -8721 11272 -8685
rect 11310 -8721 11330 -8685
rect 11256 -8759 11330 -8721
rect 11488 -8687 11562 -8649
rect 11488 -8723 11508 -8687
rect 11546 -8723 11562 -8687
rect 11488 -8759 11562 -8723
rect 11678 -8685 11752 -8649
rect 11678 -8721 11694 -8685
rect 11732 -8721 11752 -8685
rect 11678 -8759 11752 -8721
rect 11910 -8687 11984 -8649
rect 11910 -8723 11930 -8687
rect 11968 -8723 11984 -8687
rect 11910 -8759 11984 -8723
rect 12100 -8685 12174 -8649
rect 12100 -8721 12116 -8685
rect 12154 -8721 12174 -8685
rect 12100 -8759 12174 -8721
rect 12349 -8687 12407 -8649
rect 12349 -8721 12361 -8687
rect 12395 -8721 12407 -8687
rect 12349 -8759 12407 -8721
rect 13207 -8687 13265 -8649
rect 13207 -8721 13219 -8687
rect 13253 -8721 13265 -8687
rect 13207 -8759 13265 -8721
rect 13410 -8687 13484 -8649
rect 13410 -8723 13430 -8687
rect 13468 -8723 13484 -8687
rect 13410 -8759 13484 -8723
rect 13600 -8685 13674 -8649
rect 13600 -8721 13616 -8685
rect 13654 -8721 13674 -8685
rect 13600 -8759 13674 -8721
rect 13780 -8687 13854 -8649
rect 13780 -8723 13800 -8687
rect 13838 -8723 13854 -8687
rect 13780 -8759 13854 -8723
rect 13970 -8685 14044 -8649
rect 13970 -8721 13986 -8685
rect 14024 -8721 14044 -8685
rect 13970 -8759 14044 -8721
rect 14202 -8687 14276 -8649
rect 14202 -8723 14222 -8687
rect 14260 -8723 14276 -8687
rect 14202 -8759 14276 -8723
rect 14392 -8685 14466 -8649
rect 14392 -8721 14408 -8685
rect 14446 -8721 14466 -8685
rect 14392 -8759 14466 -8721
rect 14624 -8687 14698 -8649
rect 14624 -8723 14644 -8687
rect 14682 -8723 14698 -8687
rect 14624 -8759 14698 -8723
rect 14814 -8685 14888 -8649
rect 14814 -8721 14830 -8685
rect 14868 -8721 14888 -8685
rect 14814 -8759 14888 -8721
rect 15012 -8686 15070 -8648
rect 15012 -8720 15024 -8686
rect 15058 -8720 15070 -8686
rect 15012 -8758 15070 -8720
rect 15870 -8686 15928 -8648
rect 15870 -8720 15882 -8686
rect 15916 -8720 15928 -8686
rect 15870 -8758 15928 -8720
rect 16064 -8687 16138 -8649
rect 16064 -8723 16084 -8687
rect 16122 -8723 16138 -8687
rect 16064 -8759 16138 -8723
rect 16254 -8685 16328 -8649
rect 16254 -8721 16270 -8685
rect 16308 -8721 16328 -8685
rect 16254 -8759 16328 -8721
rect 9310 -14369 9384 -14331
rect 9310 -14405 9330 -14369
rect 9368 -14405 9384 -14369
rect 9310 -14441 9384 -14405
rect 9500 -14367 9574 -14331
rect 9500 -14403 9516 -14367
rect 9554 -14403 9574 -14367
rect 9500 -14441 9574 -14403
rect 9671 -14369 9729 -14331
rect 9671 -14403 9683 -14369
rect 9717 -14403 9729 -14369
rect 9671 -14441 9729 -14403
rect 10529 -14369 10587 -14331
rect 10529 -14403 10541 -14369
rect 10575 -14403 10587 -14369
rect 10529 -14441 10587 -14403
rect 10696 -14370 10770 -14332
rect 10696 -14406 10716 -14370
rect 10754 -14406 10770 -14370
rect 10696 -14442 10770 -14406
rect 10886 -14368 10960 -14332
rect 10886 -14404 10902 -14368
rect 10940 -14404 10960 -14368
rect 10886 -14442 10960 -14404
rect 11066 -14370 11140 -14332
rect 11066 -14406 11086 -14370
rect 11124 -14406 11140 -14370
rect 11066 -14442 11140 -14406
rect 11256 -14368 11330 -14332
rect 11256 -14404 11272 -14368
rect 11310 -14404 11330 -14368
rect 11256 -14442 11330 -14404
rect 11488 -14370 11562 -14332
rect 11488 -14406 11508 -14370
rect 11546 -14406 11562 -14370
rect 11488 -14442 11562 -14406
rect 11678 -14368 11752 -14332
rect 11678 -14404 11694 -14368
rect 11732 -14404 11752 -14368
rect 11678 -14442 11752 -14404
rect 11910 -14370 11984 -14332
rect 11910 -14406 11930 -14370
rect 11968 -14406 11984 -14370
rect 11910 -14442 11984 -14406
rect 12100 -14368 12174 -14332
rect 12100 -14404 12116 -14368
rect 12154 -14404 12174 -14368
rect 12100 -14442 12174 -14404
rect 12347 -14369 12406 -14331
rect 12347 -14403 12360 -14369
rect 12394 -14403 12406 -14369
rect 12347 -14438 12406 -14403
rect 12348 -14441 12406 -14438
rect 13206 -14369 13264 -14331
rect 13206 -14403 13218 -14369
rect 13252 -14403 13264 -14369
rect 13206 -14441 13264 -14403
rect 13410 -14366 13484 -14328
rect 13410 -14402 13430 -14366
rect 13468 -14402 13484 -14366
rect 13410 -14438 13484 -14402
rect 13600 -14364 13674 -14328
rect 13600 -14400 13616 -14364
rect 13654 -14400 13674 -14364
rect 13600 -14438 13674 -14400
rect 13780 -14366 13854 -14328
rect 13780 -14402 13800 -14366
rect 13838 -14402 13854 -14366
rect 13780 -14438 13854 -14402
rect 13970 -14364 14044 -14328
rect 13970 -14400 13986 -14364
rect 14024 -14400 14044 -14364
rect 13970 -14438 14044 -14400
rect 14202 -14366 14276 -14328
rect 14202 -14402 14222 -14366
rect 14260 -14402 14276 -14366
rect 14202 -14438 14276 -14402
rect 14392 -14364 14466 -14328
rect 14392 -14400 14408 -14364
rect 14446 -14400 14466 -14364
rect 14392 -14438 14466 -14400
rect 14624 -14366 14698 -14328
rect 14624 -14402 14644 -14366
rect 14682 -14402 14698 -14366
rect 14624 -14438 14698 -14402
rect 14814 -14364 14888 -14328
rect 14814 -14400 14830 -14364
rect 14868 -14400 14888 -14364
rect 14814 -14438 14888 -14400
rect 15012 -14368 15070 -14330
rect 15012 -14402 15024 -14368
rect 15058 -14402 15070 -14368
rect 15012 -14440 15070 -14402
rect 15870 -14368 15928 -14330
rect 15870 -14402 15882 -14368
rect 15916 -14402 15928 -14368
rect 15870 -14440 15928 -14402
rect 16008 -14369 16082 -14331
rect 16008 -14405 16028 -14369
rect 16066 -14405 16082 -14369
rect 16008 -14441 16082 -14405
rect 16198 -14367 16272 -14331
rect 16198 -14403 16214 -14367
rect 16252 -14403 16272 -14367
rect 16198 -14441 16272 -14403
rect 16642 -19634 16700 -19622
rect 9355 -20293 9429 -20255
rect 9355 -20329 9375 -20293
rect 9413 -20329 9429 -20293
rect 9355 -20365 9429 -20329
rect 9545 -20291 9619 -20255
rect 9545 -20327 9561 -20291
rect 9599 -20327 9619 -20291
rect 9545 -20365 9619 -20327
rect 9679 -20294 9737 -20256
rect 9679 -20328 9691 -20294
rect 9725 -20328 9737 -20294
rect 9679 -20366 9737 -20328
rect 10537 -20294 10595 -20256
rect 10537 -20328 10549 -20294
rect 10583 -20328 10595 -20294
rect 10537 -20366 10595 -20328
rect 10696 -20295 10770 -20257
rect 10696 -20331 10716 -20295
rect 10754 -20331 10770 -20295
rect 10696 -20367 10770 -20331
rect 10886 -20293 10960 -20257
rect 10886 -20329 10902 -20293
rect 10940 -20329 10960 -20293
rect 10886 -20367 10960 -20329
rect 11066 -20295 11140 -20257
rect 11066 -20331 11086 -20295
rect 11124 -20331 11140 -20295
rect 11066 -20367 11140 -20331
rect 11256 -20293 11330 -20257
rect 11256 -20329 11272 -20293
rect 11310 -20329 11330 -20293
rect 11256 -20367 11330 -20329
rect 11488 -20295 11562 -20257
rect 11488 -20331 11508 -20295
rect 11546 -20331 11562 -20295
rect 11488 -20367 11562 -20331
rect 11678 -20293 11752 -20257
rect 11678 -20329 11694 -20293
rect 11732 -20329 11752 -20293
rect 11678 -20367 11752 -20329
rect 11910 -20295 11984 -20257
rect 11910 -20331 11930 -20295
rect 11968 -20331 11984 -20295
rect 11910 -20367 11984 -20331
rect 12100 -20293 12174 -20257
rect 12100 -20329 12116 -20293
rect 12154 -20329 12174 -20293
rect 12100 -20367 12174 -20329
rect 12349 -20294 12407 -20256
rect 12349 -20328 12361 -20294
rect 12395 -20328 12407 -20294
rect 12349 -20366 12407 -20328
rect 13207 -20294 13265 -20256
rect 13207 -20328 13219 -20294
rect 13253 -20328 13265 -20294
rect 13207 -20366 13265 -20328
rect 13397 -20295 13471 -20257
rect 13397 -20331 13417 -20295
rect 13455 -20331 13471 -20295
rect 13397 -20367 13471 -20331
rect 13587 -20293 13661 -20257
rect 13587 -20329 13603 -20293
rect 13641 -20329 13661 -20293
rect 13587 -20367 13661 -20329
rect 13767 -20295 13841 -20257
rect 13767 -20331 13787 -20295
rect 13825 -20331 13841 -20295
rect 13767 -20367 13841 -20331
rect 13957 -20293 14031 -20257
rect 13957 -20329 13973 -20293
rect 14011 -20329 14031 -20293
rect 13957 -20367 14031 -20329
rect 14189 -20295 14263 -20257
rect 14189 -20331 14209 -20295
rect 14247 -20331 14263 -20295
rect 14189 -20367 14263 -20331
rect 14379 -20293 14453 -20257
rect 14379 -20329 14395 -20293
rect 14433 -20329 14453 -20293
rect 14379 -20367 14453 -20329
rect 14611 -20295 14685 -20257
rect 14611 -20331 14631 -20295
rect 14669 -20331 14685 -20295
rect 14611 -20367 14685 -20331
rect 14801 -20293 14875 -20257
rect 14801 -20329 14817 -20293
rect 14855 -20329 14875 -20293
rect 14801 -20367 14875 -20329
rect 15012 -20293 15070 -20255
rect 15012 -20327 15024 -20293
rect 15058 -20327 15070 -20293
rect 15012 -20365 15070 -20327
rect 15870 -20293 15928 -20255
rect 15870 -20327 15882 -20293
rect 15916 -20327 15928 -20293
rect 15870 -20365 15928 -20327
rect 16642 -19946 16654 -19634
rect 16688 -19946 16700 -19634
rect 16642 -19958 16700 -19946
rect 16730 -19634 16788 -19622
rect 16730 -19946 16742 -19634
rect 16776 -19946 16788 -19634
rect 16730 -19958 16788 -19946
rect 17032 -19636 17090 -19624
rect 17032 -19948 17044 -19636
rect 17078 -19948 17090 -19636
rect 17032 -19960 17090 -19948
rect 17120 -19636 17178 -19624
rect 17120 -19948 17132 -19636
rect 17166 -19948 17178 -19636
rect 17120 -19960 17178 -19948
<< ndiffc >>
rect 1098 4256 1132 4344
rect 1186 4256 1220 4344
rect 1314 4258 1348 4346
rect 1402 4258 1436 4346
rect 1532 4258 1566 4346
rect 1620 4258 1654 4346
rect 1754 4256 1788 4344
rect 1842 4256 1876 4344
rect 6284 4274 6318 4362
rect 6372 4274 6406 4362
rect 6500 4276 6534 4364
rect 6588 4276 6622 4364
rect 6718 4276 6752 4364
rect 6806 4276 6840 4364
rect 6940 4274 6974 4362
rect 7028 4274 7062 4362
rect 11460 4286 11494 4374
rect 11548 4286 11582 4374
rect 11676 4288 11710 4376
rect 11764 4288 11798 4376
rect 11894 4288 11928 4376
rect 11982 4288 12016 4376
rect 12116 4286 12150 4374
rect 12204 4286 12238 4374
rect 17116 4078 17150 4166
rect 17204 4078 17238 4166
rect 17332 4080 17366 4168
rect 17420 4080 17454 4168
rect 17550 4080 17584 4168
rect 17638 4080 17672 4168
rect 17772 4078 17806 4166
rect 17860 4078 17894 4166
rect 8786 3409 8820 3559
rect 9044 3409 9078 3559
rect 9302 3409 9336 3559
rect 9560 3409 9594 3559
rect 9800 3409 9834 3559
rect 10058 3409 10092 3559
rect 10316 3409 10350 3559
rect 10574 3409 10608 3559
rect -61818 3102 -61784 3190
rect -61722 3102 -61688 3190
rect -61626 3102 -61592 3190
rect -61530 3102 -61496 3190
rect -61434 3102 -61400 3190
rect 8786 2853 8820 3003
rect 9044 2853 9078 3003
rect 9302 2853 9336 3003
rect 9560 2853 9594 3003
rect 9800 2853 9834 3003
rect 10058 2853 10092 3003
rect 10316 2853 10350 3003
rect 10574 2853 10608 3003
rect 2626 2388 2660 2476
rect 2884 2388 2918 2476
rect 3102 2390 3136 2478
rect 3960 2390 3994 2478
rect 4074 2390 4108 2478
rect 4932 2390 4966 2478
rect 5160 2388 5194 2476
rect 5418 2388 5452 2476
rect 9107 1740 9141 1828
rect 9565 1740 9599 1828
rect 9702 1740 9736 1828
rect 10160 1740 10194 1828
rect 13318 1020 13352 2408
rect 13576 1020 13610 2408
rect 13868 2386 13902 2774
rect 14126 2386 14160 2774
rect 14384 2386 14418 2774
rect 14642 2386 14676 2774
rect 14868 2386 14902 2774
rect 15126 2386 15160 2774
rect 15384 2386 15418 2774
rect 15642 2386 15676 2774
rect 13868 1430 13902 1818
rect 14126 1430 14160 1818
rect 14384 1430 14418 1818
rect 14642 1430 14676 1818
rect 14868 1430 14902 1818
rect 15126 1430 15160 1818
rect 15384 1430 15418 1818
rect 15642 1430 15676 1818
rect 13868 474 13902 862
rect 14126 474 14160 862
rect 14384 474 14418 862
rect 14642 474 14676 862
rect 14868 474 14902 862
rect 15126 474 15160 862
rect 15384 474 15418 862
rect 15642 474 15676 862
rect 15916 970 15950 2358
rect 16174 970 16208 2358
rect 26886 2072 26920 2196
rect 26982 2072 27016 2196
rect 27078 2072 27112 2196
rect 27498 2080 27532 2204
rect 27594 2080 27628 2204
rect 27690 2080 27724 2204
rect 28076 2076 28110 2200
rect 28172 2076 28206 2200
rect 28268 2076 28302 2200
rect 28650 2084 28684 2208
rect 28746 2084 28780 2208
rect 28842 2084 28876 2208
rect 29228 2084 29262 2208
rect 29324 2084 29358 2208
rect 29420 2084 29454 2208
rect 29806 2084 29840 2208
rect 29902 2084 29936 2208
rect 29998 2084 30032 2208
rect 30388 2088 30422 2212
rect 30484 2088 30518 2212
rect 30580 2088 30614 2212
rect 30964 2084 30998 2208
rect 31060 2084 31094 2208
rect 31156 2084 31190 2208
rect 31534 2080 31568 2204
rect 31630 2080 31664 2204
rect 31726 2080 31760 2204
rect 28944 -266 28978 358
rect 29040 -266 29074 358
rect 29136 -266 29170 358
rect 29232 -266 29266 358
rect 29328 -266 29362 358
rect 29424 -266 29458 358
rect 29520 -266 29554 358
rect 29616 -266 29650 358
rect 29712 -266 29746 358
rect 29808 -266 29842 358
rect 8769 -1434 8803 -1400
rect 8853 -1460 8887 -1426
rect 8937 -1434 8971 -1400
rect 9059 -1464 9093 -1430
rect 9192 -1458 9226 -1424
rect 9299 -1458 9333 -1424
rect 9645 -1460 9679 -1426
rect 9757 -1464 9791 -1430
rect 9867 -1460 9901 -1426
rect 10079 -1464 10113 -1430
rect 10297 -1444 10331 -1410
rect 10401 -1421 10435 -1387
rect 10485 -1388 10519 -1354
rect 10485 -1456 10519 -1422
rect 10589 -1434 10623 -1400
rect 10686 -1440 10720 -1406
rect 10770 -1410 10804 -1376
rect 11235 -1434 11269 -1400
rect 11319 -1460 11353 -1426
rect 11403 -1434 11437 -1400
rect 11525 -1464 11559 -1430
rect 11658 -1458 11692 -1424
rect 11765 -1458 11799 -1424
rect 12111 -1460 12145 -1426
rect 12223 -1464 12257 -1430
rect 12333 -1460 12367 -1426
rect 12545 -1464 12579 -1430
rect 12763 -1444 12797 -1410
rect 12867 -1421 12901 -1387
rect 12951 -1388 12985 -1354
rect 12951 -1456 12985 -1422
rect 13055 -1434 13089 -1400
rect 13152 -1440 13186 -1406
rect 13236 -1410 13270 -1376
rect 10189 -2190 10223 -2156
rect 10189 -2262 10223 -2228
rect 10273 -2190 10307 -2156
rect 10273 -2262 10307 -2228
rect 10357 -2190 10391 -2156
rect 10357 -2262 10391 -2228
rect 11235 -2236 11269 -2202
rect 11319 -2262 11353 -2228
rect 11403 -2236 11437 -2202
rect 11525 -2266 11559 -2232
rect 11658 -2260 11692 -2226
rect 11765 -2260 11799 -2226
rect 12111 -2262 12145 -2228
rect 12223 -2266 12257 -2232
rect 12333 -2262 12367 -2228
rect 12545 -2266 12579 -2232
rect 12763 -2246 12797 -2212
rect 12867 -2223 12901 -2189
rect 12951 -2190 12985 -2156
rect 12951 -2258 12985 -2224
rect 13055 -2236 13089 -2202
rect 13152 -2242 13186 -2208
rect 13236 -2212 13270 -2178
rect -9123 -4704 -9089 -4670
rect -9039 -4730 -9005 -4696
rect -8955 -4704 -8921 -4670
rect -8833 -4734 -8799 -4700
rect -8700 -4728 -8666 -4694
rect -8593 -4728 -8559 -4694
rect -8247 -4730 -8213 -4696
rect -8135 -4734 -8101 -4700
rect -8025 -4730 -7991 -4696
rect -7813 -4734 -7779 -4700
rect -7595 -4714 -7561 -4680
rect -7491 -4691 -7457 -4657
rect -7407 -4658 -7373 -4624
rect -7407 -4726 -7373 -4692
rect -7303 -4704 -7269 -4670
rect -7206 -4710 -7172 -4676
rect -7122 -4680 -7088 -4646
rect -7007 -4704 -6973 -4670
rect -6923 -4730 -6889 -4696
rect -6839 -4704 -6805 -4670
rect -6717 -4734 -6683 -4700
rect -6584 -4728 -6550 -4694
rect -6477 -4728 -6443 -4694
rect -6131 -4730 -6097 -4696
rect -6019 -4734 -5985 -4700
rect -5909 -4730 -5875 -4696
rect -5697 -4734 -5663 -4700
rect -5479 -4714 -5445 -4680
rect -5375 -4691 -5341 -4657
rect -5291 -4658 -5257 -4624
rect -5291 -4726 -5257 -4692
rect -5187 -4704 -5153 -4670
rect -5090 -4710 -5056 -4676
rect -5006 -4680 -4972 -4646
rect -4891 -4704 -4857 -4670
rect -4807 -4730 -4773 -4696
rect -4723 -4704 -4689 -4670
rect -4601 -4734 -4567 -4700
rect -4468 -4728 -4434 -4694
rect -4361 -4728 -4327 -4694
rect -4015 -4730 -3981 -4696
rect -3903 -4734 -3869 -4700
rect -3793 -4730 -3759 -4696
rect -3581 -4734 -3547 -4700
rect -3363 -4714 -3329 -4680
rect -3259 -4691 -3225 -4657
rect -3175 -4658 -3141 -4624
rect -3175 -4726 -3141 -4692
rect -3071 -4704 -3037 -4670
rect -2974 -4710 -2940 -4676
rect -2890 -4680 -2856 -4646
rect -2775 -4704 -2741 -4670
rect -2691 -4730 -2657 -4696
rect -2607 -4704 -2573 -4670
rect -2485 -4734 -2451 -4700
rect -2352 -4728 -2318 -4694
rect -2245 -4728 -2211 -4694
rect -1899 -4730 -1865 -4696
rect -1787 -4734 -1753 -4700
rect -1677 -4730 -1643 -4696
rect -1465 -4734 -1431 -4700
rect -1247 -4714 -1213 -4680
rect -1143 -4691 -1109 -4657
rect -1059 -4658 -1025 -4624
rect -1059 -4726 -1025 -4692
rect -955 -4704 -921 -4670
rect -858 -4710 -824 -4676
rect -774 -4680 -740 -4646
rect -659 -4704 -625 -4670
rect -575 -4730 -541 -4696
rect -491 -4704 -457 -4670
rect -369 -4734 -335 -4700
rect -236 -4728 -202 -4694
rect -129 -4728 -95 -4694
rect 217 -4730 251 -4696
rect 329 -4734 363 -4700
rect 439 -4730 473 -4696
rect 651 -4734 685 -4700
rect 869 -4714 903 -4680
rect 973 -4691 1007 -4657
rect 1057 -4658 1091 -4624
rect 1057 -4726 1091 -4692
rect 1161 -4704 1195 -4670
rect 1258 -4710 1292 -4676
rect 1342 -4680 1376 -4646
rect 1457 -4704 1491 -4670
rect 1541 -4730 1575 -4696
rect 1625 -4704 1659 -4670
rect 1747 -4734 1781 -4700
rect 1880 -4728 1914 -4694
rect 1987 -4728 2021 -4694
rect 2333 -4730 2367 -4696
rect 2445 -4734 2479 -4700
rect 2555 -4730 2589 -4696
rect 2767 -4734 2801 -4700
rect 2985 -4714 3019 -4680
rect 3089 -4691 3123 -4657
rect 3173 -4658 3207 -4624
rect 3173 -4726 3207 -4692
rect 3277 -4704 3311 -4670
rect 3374 -4710 3408 -4676
rect 3458 -4680 3492 -4646
rect 3573 -4704 3607 -4670
rect 3657 -4730 3691 -4696
rect 3741 -4704 3775 -4670
rect 3863 -4734 3897 -4700
rect 3996 -4728 4030 -4694
rect 4103 -4728 4137 -4694
rect 4449 -4730 4483 -4696
rect 4561 -4734 4595 -4700
rect 4671 -4730 4705 -4696
rect 4883 -4734 4917 -4700
rect 5101 -4714 5135 -4680
rect 5205 -4691 5239 -4657
rect 5289 -4658 5323 -4624
rect 5289 -4726 5323 -4692
rect 5393 -4704 5427 -4670
rect 5490 -4710 5524 -4676
rect 5574 -4680 5608 -4646
rect 5689 -4704 5723 -4670
rect 5773 -4730 5807 -4696
rect 5857 -4704 5891 -4670
rect 5979 -4734 6013 -4700
rect 6112 -4728 6146 -4694
rect 6219 -4728 6253 -4694
rect 6565 -4730 6599 -4696
rect 6677 -4734 6711 -4700
rect 6787 -4730 6821 -4696
rect 6999 -4734 7033 -4700
rect 7217 -4714 7251 -4680
rect 7321 -4691 7355 -4657
rect 7405 -4658 7439 -4624
rect 7405 -4726 7439 -4692
rect 7509 -4704 7543 -4670
rect 7606 -4710 7640 -4676
rect 7690 -4680 7724 -4646
rect 7805 -4704 7839 -4670
rect 7889 -4730 7923 -4696
rect 7973 -4704 8007 -4670
rect 8095 -4734 8129 -4700
rect 8228 -4728 8262 -4694
rect 8335 -4728 8369 -4694
rect 8681 -4730 8715 -4696
rect 8793 -4734 8827 -4700
rect 8903 -4730 8937 -4696
rect 9115 -4734 9149 -4700
rect 9333 -4714 9367 -4680
rect 9437 -4691 9471 -4657
rect 9521 -4658 9555 -4624
rect 9521 -4726 9555 -4692
rect 9625 -4704 9659 -4670
rect 9722 -4710 9756 -4676
rect 9806 -4680 9840 -4646
rect 9921 -4704 9955 -4670
rect 10005 -4730 10039 -4696
rect 10089 -4704 10123 -4670
rect 10211 -4734 10245 -4700
rect 10344 -4728 10378 -4694
rect 10451 -4728 10485 -4694
rect 10797 -4730 10831 -4696
rect 10909 -4734 10943 -4700
rect 11019 -4730 11053 -4696
rect 11231 -4734 11265 -4700
rect 11449 -4714 11483 -4680
rect 11553 -4691 11587 -4657
rect 11637 -4658 11671 -4624
rect 11637 -4726 11671 -4692
rect 11741 -4704 11775 -4670
rect 11838 -4710 11872 -4676
rect 11922 -4680 11956 -4646
rect 12037 -4704 12071 -4670
rect 12121 -4730 12155 -4696
rect 12205 -4704 12239 -4670
rect 12327 -4734 12361 -4700
rect 12460 -4728 12494 -4694
rect 12567 -4728 12601 -4694
rect 12913 -4730 12947 -4696
rect 13025 -4734 13059 -4700
rect 13135 -4730 13169 -4696
rect 13347 -4734 13381 -4700
rect 13565 -4714 13599 -4680
rect 13669 -4691 13703 -4657
rect 13753 -4658 13787 -4624
rect 13753 -4726 13787 -4692
rect 13857 -4704 13891 -4670
rect 13954 -4710 13988 -4676
rect 14038 -4680 14072 -4646
rect 14153 -4704 14187 -4670
rect 14237 -4730 14271 -4696
rect 14321 -4704 14355 -4670
rect 14443 -4734 14477 -4700
rect 14576 -4728 14610 -4694
rect 14683 -4728 14717 -4694
rect 15029 -4730 15063 -4696
rect 15141 -4734 15175 -4700
rect 15251 -4730 15285 -4696
rect 15463 -4734 15497 -4700
rect 15681 -4714 15715 -4680
rect 15785 -4691 15819 -4657
rect 15869 -4658 15903 -4624
rect 15869 -4726 15903 -4692
rect 15973 -4704 16007 -4670
rect 16070 -4710 16104 -4676
rect 16154 -4680 16188 -4646
rect 16269 -4704 16303 -4670
rect 16353 -4730 16387 -4696
rect 16437 -4704 16471 -4670
rect 16559 -4734 16593 -4700
rect 16692 -4728 16726 -4694
rect 16799 -4728 16833 -4694
rect 17145 -4730 17179 -4696
rect 17257 -4734 17291 -4700
rect 17367 -4730 17401 -4696
rect 17579 -4734 17613 -4700
rect 17797 -4714 17831 -4680
rect 17901 -4691 17935 -4657
rect 17985 -4658 18019 -4624
rect 17985 -4726 18019 -4692
rect 18089 -4704 18123 -4670
rect 18186 -4710 18220 -4676
rect 18270 -4680 18304 -4646
rect 18385 -4704 18419 -4670
rect 18469 -4730 18503 -4696
rect 18553 -4704 18587 -4670
rect 18675 -4734 18709 -4700
rect 18808 -4728 18842 -4694
rect 18915 -4728 18949 -4694
rect 19261 -4730 19295 -4696
rect 19373 -4734 19407 -4700
rect 19483 -4730 19517 -4696
rect 19695 -4734 19729 -4700
rect 19913 -4714 19947 -4680
rect 20017 -4691 20051 -4657
rect 20101 -4658 20135 -4624
rect 20101 -4726 20135 -4692
rect 20205 -4704 20239 -4670
rect 20302 -4710 20336 -4676
rect 20386 -4680 20420 -4646
rect 20501 -4704 20535 -4670
rect 20585 -4730 20619 -4696
rect 20669 -4704 20703 -4670
rect 20791 -4734 20825 -4700
rect 20924 -4728 20958 -4694
rect 21031 -4728 21065 -4694
rect 21377 -4730 21411 -4696
rect 21489 -4734 21523 -4700
rect 21599 -4730 21633 -4696
rect 21811 -4734 21845 -4700
rect 22029 -4714 22063 -4680
rect 22133 -4691 22167 -4657
rect 22217 -4658 22251 -4624
rect 22217 -4726 22251 -4692
rect 22321 -4704 22355 -4670
rect 22418 -4710 22452 -4676
rect 22502 -4680 22536 -4646
rect 22617 -4704 22651 -4670
rect 22701 -4730 22735 -4696
rect 22785 -4704 22819 -4670
rect 22907 -4734 22941 -4700
rect 23040 -4728 23074 -4694
rect 23147 -4728 23181 -4694
rect 23493 -4730 23527 -4696
rect 23605 -4734 23639 -4700
rect 23715 -4730 23749 -4696
rect 23927 -4734 23961 -4700
rect 24145 -4714 24179 -4680
rect 24249 -4691 24283 -4657
rect 24333 -4658 24367 -4624
rect 24333 -4726 24367 -4692
rect 24437 -4704 24471 -4670
rect 24534 -4710 24568 -4676
rect 24618 -4680 24652 -4646
rect 24733 -4704 24767 -4670
rect 24817 -4730 24851 -4696
rect 24901 -4704 24935 -4670
rect 25023 -4734 25057 -4700
rect 25156 -4728 25190 -4694
rect 25263 -4728 25297 -4694
rect 25609 -4730 25643 -4696
rect 25721 -4734 25755 -4700
rect 25831 -4730 25865 -4696
rect 26043 -4734 26077 -4700
rect 26261 -4714 26295 -4680
rect 26365 -4691 26399 -4657
rect 26449 -4658 26483 -4624
rect 26449 -4726 26483 -4692
rect 26553 -4704 26587 -4670
rect 26650 -4710 26684 -4676
rect 26734 -4680 26768 -4646
rect 26849 -4704 26883 -4670
rect 26933 -4730 26967 -4696
rect 27017 -4704 27051 -4670
rect 27139 -4734 27173 -4700
rect 27272 -4728 27306 -4694
rect 27379 -4728 27413 -4694
rect 27725 -4730 27759 -4696
rect 27837 -4734 27871 -4700
rect 27947 -4730 27981 -4696
rect 28159 -4734 28193 -4700
rect 28377 -4714 28411 -4680
rect 28481 -4691 28515 -4657
rect 28565 -4658 28599 -4624
rect 28565 -4726 28599 -4692
rect 28669 -4704 28703 -4670
rect 28766 -4710 28800 -4676
rect 28850 -4680 28884 -4646
rect 28965 -4704 28999 -4670
rect 29049 -4730 29083 -4696
rect 29133 -4704 29167 -4670
rect 29255 -4734 29289 -4700
rect 29388 -4728 29422 -4694
rect 29495 -4728 29529 -4694
rect 29841 -4730 29875 -4696
rect 29953 -4734 29987 -4700
rect 30063 -4730 30097 -4696
rect 30275 -4734 30309 -4700
rect 30493 -4714 30527 -4680
rect 30597 -4691 30631 -4657
rect 30681 -4658 30715 -4624
rect 30681 -4726 30715 -4692
rect 30785 -4704 30819 -4670
rect 30882 -4710 30916 -4676
rect 30966 -4680 31000 -4646
rect 31081 -4704 31115 -4670
rect 31165 -4730 31199 -4696
rect 31249 -4704 31283 -4670
rect 31371 -4734 31405 -4700
rect 31504 -4728 31538 -4694
rect 31611 -4728 31645 -4694
rect 31957 -4730 31991 -4696
rect 32069 -4734 32103 -4700
rect 32179 -4730 32213 -4696
rect 32391 -4734 32425 -4700
rect 32609 -4714 32643 -4680
rect 32713 -4691 32747 -4657
rect 32797 -4658 32831 -4624
rect 32797 -4726 32831 -4692
rect 32901 -4704 32935 -4670
rect 32998 -4710 33032 -4676
rect 33082 -4680 33116 -4646
rect 4369 -9011 4403 -7635
rect 6027 -9011 6061 -7635
rect 7685 -9011 7719 -7635
rect 4369 -10521 4403 -9145
rect 6027 -10521 6061 -9145
rect 7685 -10521 7719 -9145
rect 4369 -12031 4403 -10655
rect 6027 -12031 6061 -10655
rect 7685 -12031 7719 -10655
rect 4369 -13541 4403 -12165
rect 6027 -13541 6061 -12165
rect 7685 -13541 7719 -12165
rect 4369 -15051 4403 -13675
rect 6027 -15051 6061 -13675
rect 7685 -15051 7719 -13675
rect 4369 -16561 4403 -15185
rect 6027 -16561 6061 -15185
rect 7685 -16561 7719 -15185
rect 4369 -18071 4403 -16695
rect 6027 -18071 6061 -16695
rect 7685 -18071 7719 -16695
rect 4369 -19581 4403 -18205
rect 6027 -19581 6061 -18205
rect 7685 -19581 7719 -18205
rect 4369 -21091 4403 -19715
rect 6027 -21091 6061 -19715
rect 7685 -21091 7719 -19715
rect 4369 -22601 4403 -21225
rect 6027 -22601 6061 -21225
rect 7685 -22601 7719 -21225
rect 4369 -24111 4403 -22735
rect 6027 -24111 6061 -22735
rect 7685 -24111 7719 -22735
rect 4369 -25621 4403 -24245
rect 6027 -25621 6061 -24245
rect 7685 -25621 7719 -24245
rect 9113 -9684 9147 -9648
rect 9113 -9754 9147 -9718
rect 9113 -9824 9147 -9788
rect 9371 -9684 9405 -9648
rect 9371 -9754 9405 -9718
rect 9371 -9824 9405 -9788
rect 9629 -9684 9663 -9648
rect 9629 -9754 9663 -9718
rect 9629 -9825 9663 -9789
rect 9887 -9684 9921 -9648
rect 9887 -9754 9921 -9718
rect 9887 -9824 9921 -9788
rect 10145 -9684 10179 -9648
rect 10145 -9754 10179 -9718
rect 10145 -9824 10179 -9788
rect 10403 -9684 10437 -9648
rect 10403 -9754 10437 -9718
rect 10403 -9824 10437 -9788
rect 10661 -9684 10695 -9648
rect 10661 -9754 10695 -9718
rect 10661 -9824 10695 -9788
rect 10919 -9684 10953 -9648
rect 10919 -9754 10953 -9718
rect 10919 -9824 10953 -9788
rect 11177 -9684 11211 -9648
rect 11177 -9754 11211 -9718
rect 11177 -9824 11211 -9788
rect 11783 -9684 11817 -9648
rect 11783 -9754 11817 -9718
rect 11783 -9824 11817 -9788
rect 12041 -9684 12075 -9648
rect 12041 -9754 12075 -9718
rect 12041 -9824 12075 -9788
rect 12299 -9684 12333 -9648
rect 12299 -9754 12333 -9718
rect 12299 -9825 12333 -9789
rect 12557 -9684 12591 -9648
rect 12557 -9754 12591 -9718
rect 12557 -9824 12591 -9788
rect 12815 -9684 12849 -9648
rect 12815 -9754 12849 -9718
rect 12815 -9824 12849 -9788
rect 13073 -9684 13107 -9648
rect 13073 -9754 13107 -9718
rect 13073 -9824 13107 -9788
rect 13331 -9684 13365 -9648
rect 13331 -9754 13365 -9718
rect 13331 -9824 13365 -9788
rect 13589 -9684 13623 -9648
rect 13589 -9754 13623 -9718
rect 13589 -9824 13623 -9788
rect 13847 -9684 13881 -9648
rect 13847 -9754 13881 -9718
rect 13847 -9824 13881 -9788
rect 14446 -9683 14480 -9647
rect 14446 -9753 14480 -9717
rect 14446 -9823 14480 -9787
rect 14704 -9683 14738 -9647
rect 14704 -9753 14738 -9717
rect 14704 -9823 14738 -9787
rect 14962 -9683 14996 -9647
rect 14962 -9753 14996 -9717
rect 14962 -9824 14996 -9788
rect 15220 -9683 15254 -9647
rect 15220 -9753 15254 -9717
rect 15220 -9823 15254 -9787
rect 15478 -9683 15512 -9647
rect 15478 -9753 15512 -9717
rect 15478 -9823 15512 -9787
rect 15736 -9683 15770 -9647
rect 15736 -9753 15770 -9717
rect 15736 -9823 15770 -9787
rect 15994 -9683 16028 -9647
rect 15994 -9753 16028 -9717
rect 15994 -9823 16028 -9787
rect 16252 -9683 16286 -9647
rect 16252 -9753 16286 -9717
rect 16252 -9823 16286 -9787
rect 16510 -9683 16544 -9647
rect 16510 -9753 16544 -9717
rect 16510 -9823 16544 -9787
rect 9113 -10102 9147 -10066
rect 9113 -10172 9147 -10136
rect 9113 -10242 9147 -10206
rect 9371 -10102 9405 -10066
rect 9371 -10172 9405 -10136
rect 9371 -10242 9405 -10206
rect 9629 -10102 9663 -10066
rect 9629 -10172 9663 -10136
rect 9629 -10243 9663 -10207
rect 9887 -10102 9921 -10066
rect 9887 -10172 9921 -10136
rect 9887 -10242 9921 -10206
rect 10145 -10102 10179 -10066
rect 10145 -10172 10179 -10136
rect 10145 -10242 10179 -10206
rect 10403 -10102 10437 -10066
rect 10403 -10172 10437 -10136
rect 10403 -10242 10437 -10206
rect 10661 -10102 10695 -10066
rect 10661 -10172 10695 -10136
rect 10661 -10242 10695 -10206
rect 10919 -10102 10953 -10066
rect 10919 -10172 10953 -10136
rect 10919 -10242 10953 -10206
rect 11177 -10102 11211 -10066
rect 11177 -10172 11211 -10136
rect 11177 -10242 11211 -10206
rect 11783 -10102 11817 -10066
rect 11783 -10172 11817 -10136
rect 11783 -10242 11817 -10206
rect 12041 -10102 12075 -10066
rect 12041 -10172 12075 -10136
rect 12041 -10242 12075 -10206
rect 12299 -10102 12333 -10066
rect 12299 -10172 12333 -10136
rect 12299 -10243 12333 -10207
rect 12557 -10102 12591 -10066
rect 12557 -10172 12591 -10136
rect 12557 -10242 12591 -10206
rect 12815 -10102 12849 -10066
rect 12815 -10172 12849 -10136
rect 12815 -10242 12849 -10206
rect 13073 -10102 13107 -10066
rect 13073 -10172 13107 -10136
rect 13073 -10242 13107 -10206
rect 13331 -10102 13365 -10066
rect 13331 -10172 13365 -10136
rect 13331 -10242 13365 -10206
rect 13589 -10102 13623 -10066
rect 13589 -10172 13623 -10136
rect 13589 -10242 13623 -10206
rect 13847 -10102 13881 -10066
rect 13847 -10172 13881 -10136
rect 13847 -10242 13881 -10206
rect 14446 -10101 14480 -10065
rect 14446 -10171 14480 -10135
rect 14446 -10241 14480 -10205
rect 14704 -10101 14738 -10065
rect 14704 -10171 14738 -10135
rect 14704 -10241 14738 -10205
rect 14962 -10101 14996 -10065
rect 14962 -10171 14996 -10135
rect 14962 -10242 14996 -10206
rect 15220 -10101 15254 -10065
rect 15220 -10171 15254 -10135
rect 15220 -10241 15254 -10205
rect 15478 -10101 15512 -10065
rect 15478 -10171 15512 -10135
rect 15478 -10241 15512 -10205
rect 15736 -10101 15770 -10065
rect 15736 -10171 15770 -10135
rect 15736 -10241 15770 -10205
rect 15994 -10101 16028 -10065
rect 15994 -10171 16028 -10135
rect 15994 -10241 16028 -10205
rect 16252 -10101 16286 -10065
rect 16252 -10171 16286 -10135
rect 16252 -10241 16286 -10205
rect 16510 -10101 16544 -10065
rect 16510 -10171 16544 -10135
rect 16510 -10241 16544 -10205
rect 9113 -10520 9147 -10484
rect 9113 -10590 9147 -10554
rect 9113 -10660 9147 -10624
rect 9371 -10520 9405 -10484
rect 9371 -10590 9405 -10554
rect 9371 -10660 9405 -10624
rect 9629 -10520 9663 -10484
rect 9629 -10590 9663 -10554
rect 9629 -10661 9663 -10625
rect 9887 -10520 9921 -10484
rect 9887 -10590 9921 -10554
rect 9887 -10660 9921 -10624
rect 10145 -10520 10179 -10484
rect 10145 -10590 10179 -10554
rect 10145 -10660 10179 -10624
rect 10403 -10520 10437 -10484
rect 10403 -10590 10437 -10554
rect 10403 -10660 10437 -10624
rect 10661 -10520 10695 -10484
rect 10661 -10590 10695 -10554
rect 10661 -10660 10695 -10624
rect 10919 -10520 10953 -10484
rect 10919 -10590 10953 -10554
rect 10919 -10660 10953 -10624
rect 11177 -10520 11211 -10484
rect 11177 -10590 11211 -10554
rect 11177 -10660 11211 -10624
rect 11783 -10520 11817 -10484
rect 11783 -10590 11817 -10554
rect 11783 -10660 11817 -10624
rect 12041 -10520 12075 -10484
rect 12041 -10590 12075 -10554
rect 12041 -10660 12075 -10624
rect 12299 -10520 12333 -10484
rect 12299 -10590 12333 -10554
rect 12299 -10661 12333 -10625
rect 12557 -10520 12591 -10484
rect 12557 -10590 12591 -10554
rect 12557 -10660 12591 -10624
rect 12815 -10520 12849 -10484
rect 12815 -10590 12849 -10554
rect 12815 -10660 12849 -10624
rect 13073 -10520 13107 -10484
rect 13073 -10590 13107 -10554
rect 13073 -10660 13107 -10624
rect 13331 -10520 13365 -10484
rect 13331 -10590 13365 -10554
rect 13331 -10660 13365 -10624
rect 13589 -10520 13623 -10484
rect 13589 -10590 13623 -10554
rect 13589 -10660 13623 -10624
rect 13847 -10520 13881 -10484
rect 13847 -10590 13881 -10554
rect 13847 -10660 13881 -10624
rect 14446 -10519 14480 -10483
rect 14446 -10589 14480 -10553
rect 14446 -10659 14480 -10623
rect 14704 -10519 14738 -10483
rect 14704 -10589 14738 -10553
rect 14704 -10659 14738 -10623
rect 14962 -10519 14996 -10483
rect 14962 -10589 14996 -10553
rect 14962 -10660 14996 -10624
rect 15220 -10519 15254 -10483
rect 15220 -10589 15254 -10553
rect 15220 -10659 15254 -10623
rect 15478 -10519 15512 -10483
rect 15478 -10589 15512 -10553
rect 15478 -10659 15512 -10623
rect 15736 -10519 15770 -10483
rect 15736 -10589 15770 -10553
rect 15736 -10659 15770 -10623
rect 15994 -10519 16028 -10483
rect 15994 -10589 16028 -10553
rect 15994 -10659 16028 -10623
rect 16252 -10519 16286 -10483
rect 16252 -10589 16286 -10553
rect 16252 -10659 16286 -10623
rect 16510 -10519 16544 -10483
rect 16510 -10589 16544 -10553
rect 16510 -10659 16544 -10623
rect 9113 -10938 9147 -10902
rect 9113 -11008 9147 -10972
rect 9113 -11078 9147 -11042
rect 9371 -10938 9405 -10902
rect 9371 -11008 9405 -10972
rect 9371 -11078 9405 -11042
rect 9629 -10938 9663 -10902
rect 9629 -11008 9663 -10972
rect 9629 -11079 9663 -11043
rect 9887 -10938 9921 -10902
rect 9887 -11008 9921 -10972
rect 9887 -11078 9921 -11042
rect 10145 -10938 10179 -10902
rect 10145 -11008 10179 -10972
rect 10145 -11078 10179 -11042
rect 10403 -10938 10437 -10902
rect 10403 -11008 10437 -10972
rect 10403 -11078 10437 -11042
rect 10661 -10938 10695 -10902
rect 10661 -11008 10695 -10972
rect 10661 -11078 10695 -11042
rect 10919 -10938 10953 -10902
rect 10919 -11008 10953 -10972
rect 10919 -11078 10953 -11042
rect 11177 -10938 11211 -10902
rect 11177 -11008 11211 -10972
rect 11177 -11078 11211 -11042
rect 11783 -10938 11817 -10902
rect 11783 -11008 11817 -10972
rect 11783 -11078 11817 -11042
rect 12041 -10938 12075 -10902
rect 12041 -11008 12075 -10972
rect 12041 -11078 12075 -11042
rect 12299 -10938 12333 -10902
rect 12299 -11008 12333 -10972
rect 12299 -11079 12333 -11043
rect 12557 -10938 12591 -10902
rect 12557 -11008 12591 -10972
rect 12557 -11078 12591 -11042
rect 12815 -10938 12849 -10902
rect 12815 -11008 12849 -10972
rect 12815 -11078 12849 -11042
rect 13073 -10938 13107 -10902
rect 13073 -11008 13107 -10972
rect 13073 -11078 13107 -11042
rect 13331 -10938 13365 -10902
rect 13331 -11008 13365 -10972
rect 13331 -11078 13365 -11042
rect 13589 -10938 13623 -10902
rect 13589 -11008 13623 -10972
rect 13589 -11078 13623 -11042
rect 13847 -10938 13881 -10902
rect 13847 -11008 13881 -10972
rect 13847 -11078 13881 -11042
rect 14446 -10937 14480 -10901
rect 14446 -11007 14480 -10971
rect 14446 -11077 14480 -11041
rect 14704 -10937 14738 -10901
rect 14704 -11007 14738 -10971
rect 14704 -11077 14738 -11041
rect 14962 -10937 14996 -10901
rect 14962 -11007 14996 -10971
rect 14962 -11078 14996 -11042
rect 15220 -10937 15254 -10901
rect 15220 -11007 15254 -10971
rect 15220 -11077 15254 -11041
rect 15478 -10937 15512 -10901
rect 15478 -11007 15512 -10971
rect 15478 -11077 15512 -11041
rect 15736 -10937 15770 -10901
rect 15736 -11007 15770 -10971
rect 15736 -11077 15770 -11041
rect 15994 -10937 16028 -10901
rect 15994 -11007 16028 -10971
rect 15994 -11077 16028 -11041
rect 16252 -10937 16286 -10901
rect 16252 -11007 16286 -10971
rect 16252 -11077 16286 -11041
rect 16510 -10937 16544 -10901
rect 16510 -11007 16544 -10971
rect 16510 -11077 16544 -11041
rect 9113 -11356 9147 -11320
rect 9113 -11426 9147 -11390
rect 9113 -11496 9147 -11460
rect 9371 -11356 9405 -11320
rect 9371 -11426 9405 -11390
rect 9371 -11496 9405 -11460
rect 9629 -11356 9663 -11320
rect 9629 -11426 9663 -11390
rect 9629 -11497 9663 -11461
rect 9887 -11356 9921 -11320
rect 9887 -11426 9921 -11390
rect 9887 -11496 9921 -11460
rect 10145 -11356 10179 -11320
rect 10145 -11426 10179 -11390
rect 10145 -11496 10179 -11460
rect 10403 -11356 10437 -11320
rect 10403 -11426 10437 -11390
rect 10403 -11496 10437 -11460
rect 10661 -11356 10695 -11320
rect 10661 -11426 10695 -11390
rect 10661 -11496 10695 -11460
rect 10919 -11356 10953 -11320
rect 10919 -11426 10953 -11390
rect 10919 -11496 10953 -11460
rect 11177 -11356 11211 -11320
rect 11177 -11426 11211 -11390
rect 11177 -11496 11211 -11460
rect 11783 -11356 11817 -11320
rect 11783 -11426 11817 -11390
rect 11783 -11496 11817 -11460
rect 12041 -11356 12075 -11320
rect 12041 -11426 12075 -11390
rect 12041 -11496 12075 -11460
rect 12299 -11356 12333 -11320
rect 12299 -11426 12333 -11390
rect 12299 -11497 12333 -11461
rect 12557 -11356 12591 -11320
rect 12557 -11426 12591 -11390
rect 12557 -11496 12591 -11460
rect 12815 -11356 12849 -11320
rect 12815 -11426 12849 -11390
rect 12815 -11496 12849 -11460
rect 13073 -11356 13107 -11320
rect 13073 -11426 13107 -11390
rect 13073 -11496 13107 -11460
rect 13331 -11356 13365 -11320
rect 13331 -11426 13365 -11390
rect 13331 -11496 13365 -11460
rect 13589 -11356 13623 -11320
rect 13589 -11426 13623 -11390
rect 13589 -11496 13623 -11460
rect 13847 -11356 13881 -11320
rect 13847 -11426 13881 -11390
rect 13847 -11496 13881 -11460
rect 14446 -11355 14480 -11319
rect 14446 -11425 14480 -11389
rect 14446 -11495 14480 -11459
rect 14704 -11355 14738 -11319
rect 14704 -11425 14738 -11389
rect 14704 -11495 14738 -11459
rect 14962 -11355 14996 -11319
rect 14962 -11425 14996 -11389
rect 14962 -11496 14996 -11460
rect 15220 -11355 15254 -11319
rect 15220 -11425 15254 -11389
rect 15220 -11495 15254 -11459
rect 15478 -11355 15512 -11319
rect 15478 -11425 15512 -11389
rect 15478 -11495 15512 -11459
rect 15736 -11355 15770 -11319
rect 15736 -11425 15770 -11389
rect 15736 -11495 15770 -11459
rect 15994 -11355 16028 -11319
rect 15994 -11425 16028 -11389
rect 15994 -11495 16028 -11459
rect 16252 -11355 16286 -11319
rect 16252 -11425 16286 -11389
rect 16252 -11495 16286 -11459
rect 16510 -11355 16544 -11319
rect 16510 -11425 16544 -11389
rect 16510 -11495 16544 -11459
rect 9113 -11774 9147 -11738
rect 9113 -11844 9147 -11808
rect 9113 -11914 9147 -11878
rect 9371 -11774 9405 -11738
rect 9371 -11844 9405 -11808
rect 9371 -11914 9405 -11878
rect 9629 -11774 9663 -11738
rect 9629 -11844 9663 -11808
rect 9629 -11915 9663 -11879
rect 9887 -11774 9921 -11738
rect 9887 -11844 9921 -11808
rect 9887 -11914 9921 -11878
rect 10145 -11774 10179 -11738
rect 10145 -11844 10179 -11808
rect 10145 -11914 10179 -11878
rect 10403 -11774 10437 -11738
rect 10403 -11844 10437 -11808
rect 10403 -11914 10437 -11878
rect 10661 -11774 10695 -11738
rect 10661 -11844 10695 -11808
rect 10661 -11914 10695 -11878
rect 10919 -11774 10953 -11738
rect 10919 -11844 10953 -11808
rect 10919 -11914 10953 -11878
rect 11177 -11774 11211 -11738
rect 11177 -11844 11211 -11808
rect 11177 -11914 11211 -11878
rect 11783 -11774 11817 -11738
rect 11783 -11844 11817 -11808
rect 11783 -11914 11817 -11878
rect 12041 -11774 12075 -11738
rect 12041 -11844 12075 -11808
rect 12041 -11914 12075 -11878
rect 12299 -11774 12333 -11738
rect 12299 -11844 12333 -11808
rect 12299 -11915 12333 -11879
rect 12557 -11774 12591 -11738
rect 12557 -11844 12591 -11808
rect 12557 -11914 12591 -11878
rect 12815 -11774 12849 -11738
rect 12815 -11844 12849 -11808
rect 12815 -11914 12849 -11878
rect 13073 -11774 13107 -11738
rect 13073 -11844 13107 -11808
rect 13073 -11914 13107 -11878
rect 13331 -11774 13365 -11738
rect 13331 -11844 13365 -11808
rect 13331 -11914 13365 -11878
rect 13589 -11774 13623 -11738
rect 13589 -11844 13623 -11808
rect 13589 -11914 13623 -11878
rect 13847 -11774 13881 -11738
rect 13847 -11844 13881 -11808
rect 13847 -11914 13881 -11878
rect 14446 -11773 14480 -11737
rect 14446 -11843 14480 -11807
rect 14446 -11913 14480 -11877
rect 14704 -11773 14738 -11737
rect 14704 -11843 14738 -11807
rect 14704 -11913 14738 -11877
rect 14962 -11773 14996 -11737
rect 14962 -11843 14996 -11807
rect 14962 -11914 14996 -11878
rect 15220 -11773 15254 -11737
rect 15220 -11843 15254 -11807
rect 15220 -11913 15254 -11877
rect 15478 -11773 15512 -11737
rect 15478 -11843 15512 -11807
rect 15478 -11913 15512 -11877
rect 15736 -11773 15770 -11737
rect 15736 -11843 15770 -11807
rect 15736 -11913 15770 -11877
rect 15994 -11773 16028 -11737
rect 15994 -11843 16028 -11807
rect 15994 -11913 16028 -11877
rect 16252 -11773 16286 -11737
rect 16252 -11843 16286 -11807
rect 16252 -11913 16286 -11877
rect 16510 -11773 16544 -11737
rect 16510 -11843 16544 -11807
rect 16510 -11913 16544 -11877
rect 9113 -12192 9147 -12156
rect 9113 -12262 9147 -12226
rect 9113 -12332 9147 -12296
rect 9371 -12192 9405 -12156
rect 9371 -12262 9405 -12226
rect 9371 -12332 9405 -12296
rect 9629 -12192 9663 -12156
rect 9629 -12262 9663 -12226
rect 9629 -12333 9663 -12297
rect 9887 -12192 9921 -12156
rect 9887 -12262 9921 -12226
rect 9887 -12332 9921 -12296
rect 10145 -12192 10179 -12156
rect 10145 -12262 10179 -12226
rect 10145 -12332 10179 -12296
rect 10403 -12192 10437 -12156
rect 10403 -12262 10437 -12226
rect 10403 -12332 10437 -12296
rect 10661 -12192 10695 -12156
rect 10661 -12262 10695 -12226
rect 10661 -12332 10695 -12296
rect 10919 -12192 10953 -12156
rect 10919 -12262 10953 -12226
rect 10919 -12332 10953 -12296
rect 11177 -12192 11211 -12156
rect 11177 -12262 11211 -12226
rect 11177 -12332 11211 -12296
rect 11783 -12192 11817 -12156
rect 11783 -12262 11817 -12226
rect 11783 -12332 11817 -12296
rect 12041 -12192 12075 -12156
rect 12041 -12262 12075 -12226
rect 12041 -12332 12075 -12296
rect 12299 -12192 12333 -12156
rect 12299 -12262 12333 -12226
rect 12299 -12333 12333 -12297
rect 12557 -12192 12591 -12156
rect 12557 -12262 12591 -12226
rect 12557 -12332 12591 -12296
rect 12815 -12192 12849 -12156
rect 12815 -12262 12849 -12226
rect 12815 -12332 12849 -12296
rect 13073 -12192 13107 -12156
rect 13073 -12262 13107 -12226
rect 13073 -12332 13107 -12296
rect 13331 -12192 13365 -12156
rect 13331 -12262 13365 -12226
rect 13331 -12332 13365 -12296
rect 13589 -12192 13623 -12156
rect 13589 -12262 13623 -12226
rect 13589 -12332 13623 -12296
rect 13847 -12192 13881 -12156
rect 13847 -12262 13881 -12226
rect 13847 -12332 13881 -12296
rect 14446 -12191 14480 -12155
rect 14446 -12261 14480 -12225
rect 14446 -12331 14480 -12295
rect 14704 -12191 14738 -12155
rect 14704 -12261 14738 -12225
rect 14704 -12331 14738 -12295
rect 14962 -12191 14996 -12155
rect 14962 -12261 14996 -12225
rect 14962 -12332 14996 -12296
rect 15220 -12191 15254 -12155
rect 15220 -12261 15254 -12225
rect 15220 -12331 15254 -12295
rect 15478 -12191 15512 -12155
rect 15478 -12261 15512 -12225
rect 15478 -12331 15512 -12295
rect 15736 -12191 15770 -12155
rect 15736 -12261 15770 -12225
rect 15736 -12331 15770 -12295
rect 15994 -12191 16028 -12155
rect 15994 -12261 16028 -12225
rect 15994 -12331 16028 -12295
rect 16252 -12191 16286 -12155
rect 16252 -12261 16286 -12225
rect 16252 -12331 16286 -12295
rect 16510 -12191 16544 -12155
rect 16510 -12261 16544 -12225
rect 16510 -12331 16544 -12295
rect 8993 -12844 9027 -12810
rect 8993 -12914 9027 -12878
rect 8993 -12982 9027 -12948
rect 9251 -12844 9285 -12810
rect 9251 -12914 9285 -12878
rect 9251 -12982 9285 -12948
rect 9533 -12844 9567 -12810
rect 9533 -12914 9567 -12878
rect 9533 -12982 9567 -12948
rect 9791 -12844 9825 -12810
rect 9791 -12914 9825 -12878
rect 9791 -12982 9825 -12948
rect 10013 -12844 10047 -12810
rect 10013 -12914 10047 -12878
rect 10013 -12982 10047 -12948
rect 10271 -12844 10305 -12810
rect 10271 -12914 10305 -12878
rect 10271 -12982 10305 -12948
rect 10516 -12842 10550 -12808
rect 10516 -12912 10550 -12876
rect 10516 -12980 10550 -12946
rect 10774 -12842 10808 -12808
rect 10774 -12912 10808 -12876
rect 10774 -12980 10808 -12946
rect 11026 -12832 11060 -12798
rect 11026 -12902 11060 -12866
rect 11026 -12970 11060 -12936
rect 11284 -12832 11318 -12798
rect 11284 -12902 11318 -12866
rect 11284 -12970 11318 -12936
rect 11663 -12844 11697 -12810
rect 11663 -12914 11697 -12878
rect 11663 -12982 11697 -12948
rect 11921 -12844 11955 -12810
rect 11921 -12914 11955 -12878
rect 11921 -12982 11955 -12948
rect 12203 -12844 12237 -12810
rect 12203 -12914 12237 -12878
rect 12203 -12982 12237 -12948
rect 12461 -12844 12495 -12810
rect 12461 -12914 12495 -12878
rect 12461 -12982 12495 -12948
rect 12683 -12844 12717 -12810
rect 12683 -12914 12717 -12878
rect 12683 -12982 12717 -12948
rect 12941 -12844 12975 -12810
rect 12941 -12914 12975 -12878
rect 12941 -12982 12975 -12948
rect 13186 -12842 13220 -12808
rect 13186 -12912 13220 -12876
rect 13186 -12980 13220 -12946
rect 13444 -12842 13478 -12808
rect 13444 -12912 13478 -12876
rect 13444 -12980 13478 -12946
rect 13696 -12832 13730 -12798
rect 13696 -12902 13730 -12866
rect 13696 -12970 13730 -12936
rect 13954 -12832 13988 -12798
rect 13954 -12902 13988 -12866
rect 13954 -12970 13988 -12936
rect 14326 -12843 14360 -12809
rect 14326 -12913 14360 -12877
rect 14326 -12981 14360 -12947
rect 14584 -12843 14618 -12809
rect 14584 -12913 14618 -12877
rect 14584 -12981 14618 -12947
rect 14866 -12843 14900 -12809
rect 14866 -12913 14900 -12877
rect 14866 -12981 14900 -12947
rect 15124 -12843 15158 -12809
rect 15124 -12913 15158 -12877
rect 15124 -12981 15158 -12947
rect 15346 -12843 15380 -12809
rect 15346 -12913 15380 -12877
rect 15346 -12981 15380 -12947
rect 15604 -12843 15638 -12809
rect 15604 -12913 15638 -12877
rect 15604 -12981 15638 -12947
rect 15849 -12841 15883 -12807
rect 15849 -12911 15883 -12875
rect 15849 -12979 15883 -12945
rect 16107 -12841 16141 -12807
rect 16107 -12911 16141 -12875
rect 16107 -12979 16141 -12945
rect 16359 -12831 16393 -12797
rect 16359 -12901 16393 -12865
rect 16359 -12969 16393 -12935
rect 16617 -12831 16651 -12797
rect 16617 -12901 16651 -12865
rect 16617 -12969 16651 -12935
rect 9113 -15401 9147 -15365
rect 9113 -15471 9147 -15435
rect 9113 -15541 9147 -15505
rect 9371 -15401 9405 -15365
rect 9371 -15471 9405 -15435
rect 9371 -15541 9405 -15505
rect 9629 -15401 9663 -15365
rect 9629 -15471 9663 -15435
rect 9629 -15542 9663 -15506
rect 9887 -15401 9921 -15365
rect 9887 -15471 9921 -15435
rect 9887 -15541 9921 -15505
rect 10145 -15401 10179 -15365
rect 10145 -15471 10179 -15435
rect 10145 -15541 10179 -15505
rect 10403 -15401 10437 -15365
rect 10403 -15471 10437 -15435
rect 10403 -15541 10437 -15505
rect 10661 -15401 10695 -15365
rect 10661 -15471 10695 -15435
rect 10661 -15541 10695 -15505
rect 10919 -15401 10953 -15365
rect 10919 -15471 10953 -15435
rect 10919 -15541 10953 -15505
rect 11177 -15401 11211 -15365
rect 11177 -15471 11211 -15435
rect 11177 -15541 11211 -15505
rect 11783 -15401 11817 -15365
rect 11783 -15471 11817 -15435
rect 11783 -15541 11817 -15505
rect 12041 -15401 12075 -15365
rect 12041 -15471 12075 -15435
rect 12041 -15541 12075 -15505
rect 12299 -15401 12333 -15365
rect 12299 -15471 12333 -15435
rect 12299 -15542 12333 -15506
rect 12557 -15401 12591 -15365
rect 12557 -15471 12591 -15435
rect 12557 -15541 12591 -15505
rect 12815 -15401 12849 -15365
rect 12815 -15471 12849 -15435
rect 12815 -15541 12849 -15505
rect 13073 -15401 13107 -15365
rect 13073 -15471 13107 -15435
rect 13073 -15541 13107 -15505
rect 13331 -15401 13365 -15365
rect 13331 -15471 13365 -15435
rect 13331 -15541 13365 -15505
rect 13589 -15401 13623 -15365
rect 13589 -15471 13623 -15435
rect 13589 -15541 13623 -15505
rect 13847 -15401 13881 -15365
rect 13847 -15471 13881 -15435
rect 13847 -15541 13881 -15505
rect 14446 -15400 14480 -15364
rect 14446 -15470 14480 -15434
rect 14446 -15540 14480 -15504
rect 14704 -15400 14738 -15364
rect 14704 -15470 14738 -15434
rect 14704 -15540 14738 -15504
rect 14962 -15400 14996 -15364
rect 14962 -15470 14996 -15434
rect 14962 -15541 14996 -15505
rect 15220 -15400 15254 -15364
rect 15220 -15470 15254 -15434
rect 15220 -15540 15254 -15504
rect 15478 -15400 15512 -15364
rect 15478 -15470 15512 -15434
rect 15478 -15540 15512 -15504
rect 15736 -15400 15770 -15364
rect 15736 -15470 15770 -15434
rect 15736 -15540 15770 -15504
rect 15994 -15400 16028 -15364
rect 15994 -15470 16028 -15434
rect 15994 -15540 16028 -15504
rect 16252 -15400 16286 -15364
rect 16252 -15470 16286 -15434
rect 16252 -15540 16286 -15504
rect 16510 -15400 16544 -15364
rect 16510 -15470 16544 -15434
rect 16510 -15540 16544 -15504
rect 9113 -15819 9147 -15783
rect 9113 -15889 9147 -15853
rect 9113 -15959 9147 -15923
rect 9371 -15819 9405 -15783
rect 9371 -15889 9405 -15853
rect 9371 -15959 9405 -15923
rect 9629 -15819 9663 -15783
rect 9629 -15889 9663 -15853
rect 9629 -15960 9663 -15924
rect 9887 -15819 9921 -15783
rect 9887 -15889 9921 -15853
rect 9887 -15959 9921 -15923
rect 10145 -15819 10179 -15783
rect 10145 -15889 10179 -15853
rect 10145 -15959 10179 -15923
rect 10403 -15819 10437 -15783
rect 10403 -15889 10437 -15853
rect 10403 -15959 10437 -15923
rect 10661 -15819 10695 -15783
rect 10661 -15889 10695 -15853
rect 10661 -15959 10695 -15923
rect 10919 -15819 10953 -15783
rect 10919 -15889 10953 -15853
rect 10919 -15959 10953 -15923
rect 11177 -15819 11211 -15783
rect 11177 -15889 11211 -15853
rect 11177 -15959 11211 -15923
rect 11783 -15819 11817 -15783
rect 11783 -15889 11817 -15853
rect 11783 -15959 11817 -15923
rect 12041 -15819 12075 -15783
rect 12041 -15889 12075 -15853
rect 12041 -15959 12075 -15923
rect 12299 -15819 12333 -15783
rect 12299 -15889 12333 -15853
rect 12299 -15960 12333 -15924
rect 12557 -15819 12591 -15783
rect 12557 -15889 12591 -15853
rect 12557 -15959 12591 -15923
rect 12815 -15819 12849 -15783
rect 12815 -15889 12849 -15853
rect 12815 -15959 12849 -15923
rect 13073 -15819 13107 -15783
rect 13073 -15889 13107 -15853
rect 13073 -15959 13107 -15923
rect 13331 -15819 13365 -15783
rect 13331 -15889 13365 -15853
rect 13331 -15959 13365 -15923
rect 13589 -15819 13623 -15783
rect 13589 -15889 13623 -15853
rect 13589 -15959 13623 -15923
rect 13847 -15819 13881 -15783
rect 13847 -15889 13881 -15853
rect 13847 -15959 13881 -15923
rect 14446 -15818 14480 -15782
rect 14446 -15888 14480 -15852
rect 14446 -15958 14480 -15922
rect 14704 -15818 14738 -15782
rect 14704 -15888 14738 -15852
rect 14704 -15958 14738 -15922
rect 14962 -15818 14996 -15782
rect 14962 -15888 14996 -15852
rect 14962 -15959 14996 -15923
rect 15220 -15818 15254 -15782
rect 15220 -15888 15254 -15852
rect 15220 -15958 15254 -15922
rect 15478 -15818 15512 -15782
rect 15478 -15888 15512 -15852
rect 15478 -15958 15512 -15922
rect 15736 -15818 15770 -15782
rect 15736 -15888 15770 -15852
rect 15736 -15958 15770 -15922
rect 15994 -15818 16028 -15782
rect 15994 -15888 16028 -15852
rect 15994 -15958 16028 -15922
rect 16252 -15818 16286 -15782
rect 16252 -15888 16286 -15852
rect 16252 -15958 16286 -15922
rect 16510 -15818 16544 -15782
rect 16510 -15888 16544 -15852
rect 16510 -15958 16544 -15922
rect 9113 -16237 9147 -16201
rect 9113 -16307 9147 -16271
rect 9113 -16377 9147 -16341
rect 9371 -16237 9405 -16201
rect 9371 -16307 9405 -16271
rect 9371 -16377 9405 -16341
rect 9629 -16237 9663 -16201
rect 9629 -16307 9663 -16271
rect 9629 -16378 9663 -16342
rect 9887 -16237 9921 -16201
rect 9887 -16307 9921 -16271
rect 9887 -16377 9921 -16341
rect 10145 -16237 10179 -16201
rect 10145 -16307 10179 -16271
rect 10145 -16377 10179 -16341
rect 10403 -16237 10437 -16201
rect 10403 -16307 10437 -16271
rect 10403 -16377 10437 -16341
rect 10661 -16237 10695 -16201
rect 10661 -16307 10695 -16271
rect 10661 -16377 10695 -16341
rect 10919 -16237 10953 -16201
rect 10919 -16307 10953 -16271
rect 10919 -16377 10953 -16341
rect 11177 -16237 11211 -16201
rect 11177 -16307 11211 -16271
rect 11177 -16377 11211 -16341
rect 11783 -16237 11817 -16201
rect 11783 -16307 11817 -16271
rect 11783 -16377 11817 -16341
rect 12041 -16237 12075 -16201
rect 12041 -16307 12075 -16271
rect 12041 -16377 12075 -16341
rect 12299 -16237 12333 -16201
rect 12299 -16307 12333 -16271
rect 12299 -16378 12333 -16342
rect 12557 -16237 12591 -16201
rect 12557 -16307 12591 -16271
rect 12557 -16377 12591 -16341
rect 12815 -16237 12849 -16201
rect 12815 -16307 12849 -16271
rect 12815 -16377 12849 -16341
rect 13073 -16237 13107 -16201
rect 13073 -16307 13107 -16271
rect 13073 -16377 13107 -16341
rect 13331 -16237 13365 -16201
rect 13331 -16307 13365 -16271
rect 13331 -16377 13365 -16341
rect 13589 -16237 13623 -16201
rect 13589 -16307 13623 -16271
rect 13589 -16377 13623 -16341
rect 13847 -16237 13881 -16201
rect 13847 -16307 13881 -16271
rect 13847 -16377 13881 -16341
rect 14446 -16236 14480 -16200
rect 14446 -16306 14480 -16270
rect 14446 -16376 14480 -16340
rect 14704 -16236 14738 -16200
rect 14704 -16306 14738 -16270
rect 14704 -16376 14738 -16340
rect 14962 -16236 14996 -16200
rect 14962 -16306 14996 -16270
rect 14962 -16377 14996 -16341
rect 15220 -16236 15254 -16200
rect 15220 -16306 15254 -16270
rect 15220 -16376 15254 -16340
rect 15478 -16236 15512 -16200
rect 15478 -16306 15512 -16270
rect 15478 -16376 15512 -16340
rect 15736 -16236 15770 -16200
rect 15736 -16306 15770 -16270
rect 15736 -16376 15770 -16340
rect 15994 -16236 16028 -16200
rect 15994 -16306 16028 -16270
rect 15994 -16376 16028 -16340
rect 16252 -16236 16286 -16200
rect 16252 -16306 16286 -16270
rect 16252 -16376 16286 -16340
rect 16510 -16236 16544 -16200
rect 16510 -16306 16544 -16270
rect 16510 -16376 16544 -16340
rect 9113 -16655 9147 -16619
rect 9113 -16725 9147 -16689
rect 9113 -16795 9147 -16759
rect 9371 -16655 9405 -16619
rect 9371 -16725 9405 -16689
rect 9371 -16795 9405 -16759
rect 9629 -16655 9663 -16619
rect 9629 -16725 9663 -16689
rect 9629 -16796 9663 -16760
rect 9887 -16655 9921 -16619
rect 9887 -16725 9921 -16689
rect 9887 -16795 9921 -16759
rect 10145 -16655 10179 -16619
rect 10145 -16725 10179 -16689
rect 10145 -16795 10179 -16759
rect 10403 -16655 10437 -16619
rect 10403 -16725 10437 -16689
rect 10403 -16795 10437 -16759
rect 10661 -16655 10695 -16619
rect 10661 -16725 10695 -16689
rect 10661 -16795 10695 -16759
rect 10919 -16655 10953 -16619
rect 10919 -16725 10953 -16689
rect 10919 -16795 10953 -16759
rect 11177 -16655 11211 -16619
rect 11177 -16725 11211 -16689
rect 11177 -16795 11211 -16759
rect 11783 -16655 11817 -16619
rect 11783 -16725 11817 -16689
rect 11783 -16795 11817 -16759
rect 12041 -16655 12075 -16619
rect 12041 -16725 12075 -16689
rect 12041 -16795 12075 -16759
rect 12299 -16655 12333 -16619
rect 12299 -16725 12333 -16689
rect 12299 -16796 12333 -16760
rect 12557 -16655 12591 -16619
rect 12557 -16725 12591 -16689
rect 12557 -16795 12591 -16759
rect 12815 -16655 12849 -16619
rect 12815 -16725 12849 -16689
rect 12815 -16795 12849 -16759
rect 13073 -16655 13107 -16619
rect 13073 -16725 13107 -16689
rect 13073 -16795 13107 -16759
rect 13331 -16655 13365 -16619
rect 13331 -16725 13365 -16689
rect 13331 -16795 13365 -16759
rect 13589 -16655 13623 -16619
rect 13589 -16725 13623 -16689
rect 13589 -16795 13623 -16759
rect 13847 -16655 13881 -16619
rect 13847 -16725 13881 -16689
rect 13847 -16795 13881 -16759
rect 14446 -16654 14480 -16618
rect 14446 -16724 14480 -16688
rect 14446 -16794 14480 -16758
rect 14704 -16654 14738 -16618
rect 14704 -16724 14738 -16688
rect 14704 -16794 14738 -16758
rect 14962 -16654 14996 -16618
rect 14962 -16724 14996 -16688
rect 14962 -16795 14996 -16759
rect 15220 -16654 15254 -16618
rect 15220 -16724 15254 -16688
rect 15220 -16794 15254 -16758
rect 15478 -16654 15512 -16618
rect 15478 -16724 15512 -16688
rect 15478 -16794 15512 -16758
rect 15736 -16654 15770 -16618
rect 15736 -16724 15770 -16688
rect 15736 -16794 15770 -16758
rect 15994 -16654 16028 -16618
rect 15994 -16724 16028 -16688
rect 15994 -16794 16028 -16758
rect 16252 -16654 16286 -16618
rect 16252 -16724 16286 -16688
rect 16252 -16794 16286 -16758
rect 16510 -16654 16544 -16618
rect 16510 -16724 16544 -16688
rect 16510 -16794 16544 -16758
rect 9113 -17073 9147 -17037
rect 9113 -17143 9147 -17107
rect 9113 -17213 9147 -17177
rect 9371 -17073 9405 -17037
rect 9371 -17143 9405 -17107
rect 9371 -17213 9405 -17177
rect 9629 -17073 9663 -17037
rect 9629 -17143 9663 -17107
rect 9629 -17214 9663 -17178
rect 9887 -17073 9921 -17037
rect 9887 -17143 9921 -17107
rect 9887 -17213 9921 -17177
rect 10145 -17073 10179 -17037
rect 10145 -17143 10179 -17107
rect 10145 -17213 10179 -17177
rect 10403 -17073 10437 -17037
rect 10403 -17143 10437 -17107
rect 10403 -17213 10437 -17177
rect 10661 -17073 10695 -17037
rect 10661 -17143 10695 -17107
rect 10661 -17213 10695 -17177
rect 10919 -17073 10953 -17037
rect 10919 -17143 10953 -17107
rect 10919 -17213 10953 -17177
rect 11177 -17073 11211 -17037
rect 11177 -17143 11211 -17107
rect 11177 -17213 11211 -17177
rect 11783 -17073 11817 -17037
rect 11783 -17143 11817 -17107
rect 11783 -17213 11817 -17177
rect 12041 -17073 12075 -17037
rect 12041 -17143 12075 -17107
rect 12041 -17213 12075 -17177
rect 12299 -17073 12333 -17037
rect 12299 -17143 12333 -17107
rect 12299 -17214 12333 -17178
rect 12557 -17073 12591 -17037
rect 12557 -17143 12591 -17107
rect 12557 -17213 12591 -17177
rect 12815 -17073 12849 -17037
rect 12815 -17143 12849 -17107
rect 12815 -17213 12849 -17177
rect 13073 -17073 13107 -17037
rect 13073 -17143 13107 -17107
rect 13073 -17213 13107 -17177
rect 13331 -17073 13365 -17037
rect 13331 -17143 13365 -17107
rect 13331 -17213 13365 -17177
rect 13589 -17073 13623 -17037
rect 13589 -17143 13623 -17107
rect 13589 -17213 13623 -17177
rect 13847 -17073 13881 -17037
rect 13847 -17143 13881 -17107
rect 13847 -17213 13881 -17177
rect 14446 -17072 14480 -17036
rect 14446 -17142 14480 -17106
rect 14446 -17212 14480 -17176
rect 14704 -17072 14738 -17036
rect 14704 -17142 14738 -17106
rect 14704 -17212 14738 -17176
rect 14962 -17072 14996 -17036
rect 14962 -17142 14996 -17106
rect 14962 -17213 14996 -17177
rect 15220 -17072 15254 -17036
rect 15220 -17142 15254 -17106
rect 15220 -17212 15254 -17176
rect 15478 -17072 15512 -17036
rect 15478 -17142 15512 -17106
rect 15478 -17212 15512 -17176
rect 15736 -17072 15770 -17036
rect 15736 -17142 15770 -17106
rect 15736 -17212 15770 -17176
rect 15994 -17072 16028 -17036
rect 15994 -17142 16028 -17106
rect 15994 -17212 16028 -17176
rect 16252 -17072 16286 -17036
rect 16252 -17142 16286 -17106
rect 16252 -17212 16286 -17176
rect 16510 -17072 16544 -17036
rect 16510 -17142 16544 -17106
rect 16510 -17212 16544 -17176
rect 9113 -17491 9147 -17455
rect 9113 -17561 9147 -17525
rect 9113 -17631 9147 -17595
rect 9371 -17491 9405 -17455
rect 9371 -17561 9405 -17525
rect 9371 -17631 9405 -17595
rect 9629 -17491 9663 -17455
rect 9629 -17561 9663 -17525
rect 9629 -17632 9663 -17596
rect 9887 -17491 9921 -17455
rect 9887 -17561 9921 -17525
rect 9887 -17631 9921 -17595
rect 10145 -17491 10179 -17455
rect 10145 -17561 10179 -17525
rect 10145 -17631 10179 -17595
rect 10403 -17491 10437 -17455
rect 10403 -17561 10437 -17525
rect 10403 -17631 10437 -17595
rect 10661 -17491 10695 -17455
rect 10661 -17561 10695 -17525
rect 10661 -17631 10695 -17595
rect 10919 -17491 10953 -17455
rect 10919 -17561 10953 -17525
rect 10919 -17631 10953 -17595
rect 11177 -17491 11211 -17455
rect 11177 -17561 11211 -17525
rect 11177 -17631 11211 -17595
rect 11783 -17491 11817 -17455
rect 11783 -17561 11817 -17525
rect 11783 -17631 11817 -17595
rect 12041 -17491 12075 -17455
rect 12041 -17561 12075 -17525
rect 12041 -17631 12075 -17595
rect 12299 -17491 12333 -17455
rect 12299 -17561 12333 -17525
rect 12299 -17632 12333 -17596
rect 12557 -17491 12591 -17455
rect 12557 -17561 12591 -17525
rect 12557 -17631 12591 -17595
rect 12815 -17491 12849 -17455
rect 12815 -17561 12849 -17525
rect 12815 -17631 12849 -17595
rect 13073 -17491 13107 -17455
rect 13073 -17561 13107 -17525
rect 13073 -17631 13107 -17595
rect 13331 -17491 13365 -17455
rect 13331 -17561 13365 -17525
rect 13331 -17631 13365 -17595
rect 13589 -17491 13623 -17455
rect 13589 -17561 13623 -17525
rect 13589 -17631 13623 -17595
rect 13847 -17491 13881 -17455
rect 13847 -17561 13881 -17525
rect 13847 -17631 13881 -17595
rect 14446 -17490 14480 -17454
rect 14446 -17560 14480 -17524
rect 14446 -17630 14480 -17594
rect 14704 -17490 14738 -17454
rect 14704 -17560 14738 -17524
rect 14704 -17630 14738 -17594
rect 14962 -17490 14996 -17454
rect 14962 -17560 14996 -17524
rect 14962 -17631 14996 -17595
rect 15220 -17490 15254 -17454
rect 15220 -17560 15254 -17524
rect 15220 -17630 15254 -17594
rect 15478 -17490 15512 -17454
rect 15478 -17560 15512 -17524
rect 15478 -17630 15512 -17594
rect 15736 -17490 15770 -17454
rect 15736 -17560 15770 -17524
rect 15736 -17630 15770 -17594
rect 15994 -17490 16028 -17454
rect 15994 -17560 16028 -17524
rect 15994 -17630 16028 -17594
rect 16252 -17490 16286 -17454
rect 16252 -17560 16286 -17524
rect 16252 -17630 16286 -17594
rect 16510 -17490 16544 -17454
rect 16510 -17560 16544 -17524
rect 16510 -17630 16544 -17594
rect 9113 -17909 9147 -17873
rect 9113 -17979 9147 -17943
rect 9113 -18049 9147 -18013
rect 9371 -17909 9405 -17873
rect 9371 -17979 9405 -17943
rect 9371 -18049 9405 -18013
rect 9629 -17909 9663 -17873
rect 9629 -17979 9663 -17943
rect 9629 -18050 9663 -18014
rect 9887 -17909 9921 -17873
rect 9887 -17979 9921 -17943
rect 9887 -18049 9921 -18013
rect 10145 -17909 10179 -17873
rect 10145 -17979 10179 -17943
rect 10145 -18049 10179 -18013
rect 10403 -17909 10437 -17873
rect 10403 -17979 10437 -17943
rect 10403 -18049 10437 -18013
rect 10661 -17909 10695 -17873
rect 10661 -17979 10695 -17943
rect 10661 -18049 10695 -18013
rect 10919 -17909 10953 -17873
rect 10919 -17979 10953 -17943
rect 10919 -18049 10953 -18013
rect 11177 -17909 11211 -17873
rect 11177 -17979 11211 -17943
rect 11177 -18049 11211 -18013
rect 11783 -17909 11817 -17873
rect 11783 -17979 11817 -17943
rect 11783 -18049 11817 -18013
rect 12041 -17909 12075 -17873
rect 12041 -17979 12075 -17943
rect 12041 -18049 12075 -18013
rect 12299 -17909 12333 -17873
rect 12299 -17979 12333 -17943
rect 12299 -18050 12333 -18014
rect 12557 -17909 12591 -17873
rect 12557 -17979 12591 -17943
rect 12557 -18049 12591 -18013
rect 12815 -17909 12849 -17873
rect 12815 -17979 12849 -17943
rect 12815 -18049 12849 -18013
rect 13073 -17909 13107 -17873
rect 13073 -17979 13107 -17943
rect 13073 -18049 13107 -18013
rect 13331 -17909 13365 -17873
rect 13331 -17979 13365 -17943
rect 13331 -18049 13365 -18013
rect 13589 -17909 13623 -17873
rect 13589 -17979 13623 -17943
rect 13589 -18049 13623 -18013
rect 13847 -17909 13881 -17873
rect 13847 -17979 13881 -17943
rect 13847 -18049 13881 -18013
rect 14446 -17908 14480 -17872
rect 14446 -17978 14480 -17942
rect 14446 -18048 14480 -18012
rect 14704 -17908 14738 -17872
rect 14704 -17978 14738 -17942
rect 14704 -18048 14738 -18012
rect 14962 -17908 14996 -17872
rect 14962 -17978 14996 -17942
rect 14962 -18049 14996 -18013
rect 15220 -17908 15254 -17872
rect 15220 -17978 15254 -17942
rect 15220 -18048 15254 -18012
rect 15478 -17908 15512 -17872
rect 15478 -17978 15512 -17942
rect 15478 -18048 15512 -18012
rect 15736 -17908 15770 -17872
rect 15736 -17978 15770 -17942
rect 15736 -18048 15770 -18012
rect 15994 -17908 16028 -17872
rect 15994 -17978 16028 -17942
rect 15994 -18048 16028 -18012
rect 16252 -17908 16286 -17872
rect 16252 -17978 16286 -17942
rect 16252 -18048 16286 -18012
rect 16510 -17908 16544 -17872
rect 16510 -17978 16544 -17942
rect 16510 -18048 16544 -18012
rect 8993 -18561 9027 -18527
rect 8993 -18631 9027 -18595
rect 8993 -18699 9027 -18665
rect 9251 -18561 9285 -18527
rect 9251 -18631 9285 -18595
rect 9251 -18699 9285 -18665
rect 9533 -18561 9567 -18527
rect 9533 -18631 9567 -18595
rect 9533 -18699 9567 -18665
rect 9791 -18561 9825 -18527
rect 9791 -18631 9825 -18595
rect 9791 -18699 9825 -18665
rect 10013 -18561 10047 -18527
rect 10013 -18631 10047 -18595
rect 10013 -18699 10047 -18665
rect 10271 -18561 10305 -18527
rect 10271 -18631 10305 -18595
rect 10271 -18699 10305 -18665
rect 10516 -18559 10550 -18525
rect 10516 -18629 10550 -18593
rect 10516 -18697 10550 -18663
rect 10774 -18559 10808 -18525
rect 10774 -18629 10808 -18593
rect 10774 -18697 10808 -18663
rect 11026 -18549 11060 -18515
rect 11026 -18619 11060 -18583
rect 11026 -18687 11060 -18653
rect 11284 -18549 11318 -18515
rect 11284 -18619 11318 -18583
rect 11284 -18687 11318 -18653
rect 11663 -18561 11697 -18527
rect 11663 -18631 11697 -18595
rect 11663 -18699 11697 -18665
rect 11921 -18561 11955 -18527
rect 11921 -18631 11955 -18595
rect 11921 -18699 11955 -18665
rect 12203 -18561 12237 -18527
rect 12203 -18631 12237 -18595
rect 12203 -18699 12237 -18665
rect 12461 -18561 12495 -18527
rect 12461 -18631 12495 -18595
rect 12461 -18699 12495 -18665
rect 12683 -18561 12717 -18527
rect 12683 -18631 12717 -18595
rect 12683 -18699 12717 -18665
rect 12941 -18561 12975 -18527
rect 12941 -18631 12975 -18595
rect 12941 -18699 12975 -18665
rect 13186 -18559 13220 -18525
rect 13186 -18629 13220 -18593
rect 13186 -18697 13220 -18663
rect 13444 -18559 13478 -18525
rect 13444 -18629 13478 -18593
rect 13444 -18697 13478 -18663
rect 13696 -18549 13730 -18515
rect 13696 -18619 13730 -18583
rect 13696 -18687 13730 -18653
rect 13954 -18549 13988 -18515
rect 13954 -18619 13988 -18583
rect 13954 -18687 13988 -18653
rect 14326 -18560 14360 -18526
rect 14326 -18630 14360 -18594
rect 14326 -18698 14360 -18664
rect 14584 -18560 14618 -18526
rect 14584 -18630 14618 -18594
rect 14584 -18698 14618 -18664
rect 14866 -18560 14900 -18526
rect 14866 -18630 14900 -18594
rect 14866 -18698 14900 -18664
rect 15124 -18560 15158 -18526
rect 15124 -18630 15158 -18594
rect 15124 -18698 15158 -18664
rect 15346 -18560 15380 -18526
rect 15346 -18630 15380 -18594
rect 15346 -18698 15380 -18664
rect 15604 -18560 15638 -18526
rect 15604 -18630 15638 -18594
rect 15604 -18698 15638 -18664
rect 15849 -18558 15883 -18524
rect 15849 -18628 15883 -18592
rect 15849 -18696 15883 -18662
rect 16107 -18558 16141 -18524
rect 16107 -18628 16141 -18592
rect 16107 -18696 16141 -18662
rect 16359 -18548 16393 -18514
rect 16359 -18618 16393 -18582
rect 16359 -18686 16393 -18652
rect 16617 -18548 16651 -18514
rect 16617 -18618 16651 -18582
rect 16617 -18686 16651 -18652
rect 16658 -20481 16692 -20421
rect 16746 -20481 16780 -20421
rect 17048 -20481 17082 -20421
rect 17136 -20481 17170 -20421
rect 9113 -21305 9147 -21269
rect 9113 -21375 9147 -21339
rect 9113 -21445 9147 -21409
rect 9371 -21305 9405 -21269
rect 9371 -21375 9405 -21339
rect 9371 -21445 9405 -21409
rect 9629 -21305 9663 -21269
rect 9629 -21375 9663 -21339
rect 9629 -21446 9663 -21410
rect 9887 -21305 9921 -21269
rect 9887 -21375 9921 -21339
rect 9887 -21445 9921 -21409
rect 10145 -21305 10179 -21269
rect 10145 -21375 10179 -21339
rect 10145 -21445 10179 -21409
rect 10403 -21305 10437 -21269
rect 10403 -21375 10437 -21339
rect 10403 -21445 10437 -21409
rect 10661 -21305 10695 -21269
rect 10661 -21375 10695 -21339
rect 10661 -21445 10695 -21409
rect 10919 -21305 10953 -21269
rect 10919 -21375 10953 -21339
rect 10919 -21445 10953 -21409
rect 11177 -21305 11211 -21269
rect 11177 -21375 11211 -21339
rect 11177 -21445 11211 -21409
rect 11783 -21305 11817 -21269
rect 11783 -21375 11817 -21339
rect 11783 -21445 11817 -21409
rect 12041 -21305 12075 -21269
rect 12041 -21375 12075 -21339
rect 12041 -21445 12075 -21409
rect 12299 -21305 12333 -21269
rect 12299 -21375 12333 -21339
rect 12299 -21446 12333 -21410
rect 12557 -21305 12591 -21269
rect 12557 -21375 12591 -21339
rect 12557 -21445 12591 -21409
rect 12815 -21305 12849 -21269
rect 12815 -21375 12849 -21339
rect 12815 -21445 12849 -21409
rect 13073 -21305 13107 -21269
rect 13073 -21375 13107 -21339
rect 13073 -21445 13107 -21409
rect 13331 -21305 13365 -21269
rect 13331 -21375 13365 -21339
rect 13331 -21445 13365 -21409
rect 13589 -21305 13623 -21269
rect 13589 -21375 13623 -21339
rect 13589 -21445 13623 -21409
rect 13847 -21305 13881 -21269
rect 13847 -21375 13881 -21339
rect 13847 -21445 13881 -21409
rect 14446 -21304 14480 -21268
rect 14446 -21374 14480 -21338
rect 14446 -21444 14480 -21408
rect 14704 -21304 14738 -21268
rect 14704 -21374 14738 -21338
rect 14704 -21444 14738 -21408
rect 14962 -21304 14996 -21268
rect 14962 -21374 14996 -21338
rect 14962 -21445 14996 -21409
rect 15220 -21304 15254 -21268
rect 15220 -21374 15254 -21338
rect 15220 -21444 15254 -21408
rect 15478 -21304 15512 -21268
rect 15478 -21374 15512 -21338
rect 15478 -21444 15512 -21408
rect 15736 -21304 15770 -21268
rect 15736 -21374 15770 -21338
rect 15736 -21444 15770 -21408
rect 15994 -21304 16028 -21268
rect 15994 -21374 16028 -21338
rect 15994 -21444 16028 -21408
rect 16252 -21304 16286 -21268
rect 16252 -21374 16286 -21338
rect 16252 -21444 16286 -21408
rect 16510 -21304 16544 -21268
rect 16510 -21374 16544 -21338
rect 16510 -21444 16544 -21408
rect 9113 -21723 9147 -21687
rect 9113 -21793 9147 -21757
rect 9113 -21863 9147 -21827
rect 9371 -21723 9405 -21687
rect 9371 -21793 9405 -21757
rect 9371 -21863 9405 -21827
rect 9629 -21723 9663 -21687
rect 9629 -21793 9663 -21757
rect 9629 -21864 9663 -21828
rect 9887 -21723 9921 -21687
rect 9887 -21793 9921 -21757
rect 9887 -21863 9921 -21827
rect 10145 -21723 10179 -21687
rect 10145 -21793 10179 -21757
rect 10145 -21863 10179 -21827
rect 10403 -21723 10437 -21687
rect 10403 -21793 10437 -21757
rect 10403 -21863 10437 -21827
rect 10661 -21723 10695 -21687
rect 10661 -21793 10695 -21757
rect 10661 -21863 10695 -21827
rect 10919 -21723 10953 -21687
rect 10919 -21793 10953 -21757
rect 10919 -21863 10953 -21827
rect 11177 -21723 11211 -21687
rect 11177 -21793 11211 -21757
rect 11177 -21863 11211 -21827
rect 11783 -21723 11817 -21687
rect 11783 -21793 11817 -21757
rect 11783 -21863 11817 -21827
rect 12041 -21723 12075 -21687
rect 12041 -21793 12075 -21757
rect 12041 -21863 12075 -21827
rect 12299 -21723 12333 -21687
rect 12299 -21793 12333 -21757
rect 12299 -21864 12333 -21828
rect 12557 -21723 12591 -21687
rect 12557 -21793 12591 -21757
rect 12557 -21863 12591 -21827
rect 12815 -21723 12849 -21687
rect 12815 -21793 12849 -21757
rect 12815 -21863 12849 -21827
rect 13073 -21723 13107 -21687
rect 13073 -21793 13107 -21757
rect 13073 -21863 13107 -21827
rect 13331 -21723 13365 -21687
rect 13331 -21793 13365 -21757
rect 13331 -21863 13365 -21827
rect 13589 -21723 13623 -21687
rect 13589 -21793 13623 -21757
rect 13589 -21863 13623 -21827
rect 13847 -21723 13881 -21687
rect 13847 -21793 13881 -21757
rect 13847 -21863 13881 -21827
rect 14446 -21722 14480 -21686
rect 14446 -21792 14480 -21756
rect 14446 -21862 14480 -21826
rect 14704 -21722 14738 -21686
rect 14704 -21792 14738 -21756
rect 14704 -21862 14738 -21826
rect 14962 -21722 14996 -21686
rect 14962 -21792 14996 -21756
rect 14962 -21863 14996 -21827
rect 15220 -21722 15254 -21686
rect 15220 -21792 15254 -21756
rect 15220 -21862 15254 -21826
rect 15478 -21722 15512 -21686
rect 15478 -21792 15512 -21756
rect 15478 -21862 15512 -21826
rect 15736 -21722 15770 -21686
rect 15736 -21792 15770 -21756
rect 15736 -21862 15770 -21826
rect 15994 -21722 16028 -21686
rect 15994 -21792 16028 -21756
rect 15994 -21862 16028 -21826
rect 16252 -21722 16286 -21686
rect 16252 -21792 16286 -21756
rect 16252 -21862 16286 -21826
rect 16510 -21722 16544 -21686
rect 16510 -21792 16544 -21756
rect 16510 -21862 16544 -21826
rect 9113 -22141 9147 -22105
rect 9113 -22211 9147 -22175
rect 9113 -22281 9147 -22245
rect 9371 -22141 9405 -22105
rect 9371 -22211 9405 -22175
rect 9371 -22281 9405 -22245
rect 9629 -22141 9663 -22105
rect 9629 -22211 9663 -22175
rect 9629 -22282 9663 -22246
rect 9887 -22141 9921 -22105
rect 9887 -22211 9921 -22175
rect 9887 -22281 9921 -22245
rect 10145 -22141 10179 -22105
rect 10145 -22211 10179 -22175
rect 10145 -22281 10179 -22245
rect 10403 -22141 10437 -22105
rect 10403 -22211 10437 -22175
rect 10403 -22281 10437 -22245
rect 10661 -22141 10695 -22105
rect 10661 -22211 10695 -22175
rect 10661 -22281 10695 -22245
rect 10919 -22141 10953 -22105
rect 10919 -22211 10953 -22175
rect 10919 -22281 10953 -22245
rect 11177 -22141 11211 -22105
rect 11177 -22211 11211 -22175
rect 11177 -22281 11211 -22245
rect 11783 -22141 11817 -22105
rect 11783 -22211 11817 -22175
rect 11783 -22281 11817 -22245
rect 12041 -22141 12075 -22105
rect 12041 -22211 12075 -22175
rect 12041 -22281 12075 -22245
rect 12299 -22141 12333 -22105
rect 12299 -22211 12333 -22175
rect 12299 -22282 12333 -22246
rect 12557 -22141 12591 -22105
rect 12557 -22211 12591 -22175
rect 12557 -22281 12591 -22245
rect 12815 -22141 12849 -22105
rect 12815 -22211 12849 -22175
rect 12815 -22281 12849 -22245
rect 13073 -22141 13107 -22105
rect 13073 -22211 13107 -22175
rect 13073 -22281 13107 -22245
rect 13331 -22141 13365 -22105
rect 13331 -22211 13365 -22175
rect 13331 -22281 13365 -22245
rect 13589 -22141 13623 -22105
rect 13589 -22211 13623 -22175
rect 13589 -22281 13623 -22245
rect 13847 -22141 13881 -22105
rect 13847 -22211 13881 -22175
rect 13847 -22281 13881 -22245
rect 14446 -22140 14480 -22104
rect 14446 -22210 14480 -22174
rect 14446 -22280 14480 -22244
rect 14704 -22140 14738 -22104
rect 14704 -22210 14738 -22174
rect 14704 -22280 14738 -22244
rect 14962 -22140 14996 -22104
rect 14962 -22210 14996 -22174
rect 14962 -22281 14996 -22245
rect 15220 -22140 15254 -22104
rect 15220 -22210 15254 -22174
rect 15220 -22280 15254 -22244
rect 15478 -22140 15512 -22104
rect 15478 -22210 15512 -22174
rect 15478 -22280 15512 -22244
rect 15736 -22140 15770 -22104
rect 15736 -22210 15770 -22174
rect 15736 -22280 15770 -22244
rect 15994 -22140 16028 -22104
rect 15994 -22210 16028 -22174
rect 15994 -22280 16028 -22244
rect 16252 -22140 16286 -22104
rect 16252 -22210 16286 -22174
rect 16252 -22280 16286 -22244
rect 16510 -22140 16544 -22104
rect 16510 -22210 16544 -22174
rect 16510 -22280 16544 -22244
rect 9113 -22559 9147 -22523
rect 9113 -22629 9147 -22593
rect 9113 -22699 9147 -22663
rect 9371 -22559 9405 -22523
rect 9371 -22629 9405 -22593
rect 9371 -22699 9405 -22663
rect 9629 -22559 9663 -22523
rect 9629 -22629 9663 -22593
rect 9629 -22700 9663 -22664
rect 9887 -22559 9921 -22523
rect 9887 -22629 9921 -22593
rect 9887 -22699 9921 -22663
rect 10145 -22559 10179 -22523
rect 10145 -22629 10179 -22593
rect 10145 -22699 10179 -22663
rect 10403 -22559 10437 -22523
rect 10403 -22629 10437 -22593
rect 10403 -22699 10437 -22663
rect 10661 -22559 10695 -22523
rect 10661 -22629 10695 -22593
rect 10661 -22699 10695 -22663
rect 10919 -22559 10953 -22523
rect 10919 -22629 10953 -22593
rect 10919 -22699 10953 -22663
rect 11177 -22559 11211 -22523
rect 11177 -22629 11211 -22593
rect 11177 -22699 11211 -22663
rect 11783 -22559 11817 -22523
rect 11783 -22629 11817 -22593
rect 11783 -22699 11817 -22663
rect 12041 -22559 12075 -22523
rect 12041 -22629 12075 -22593
rect 12041 -22699 12075 -22663
rect 12299 -22559 12333 -22523
rect 12299 -22629 12333 -22593
rect 12299 -22700 12333 -22664
rect 12557 -22559 12591 -22523
rect 12557 -22629 12591 -22593
rect 12557 -22699 12591 -22663
rect 12815 -22559 12849 -22523
rect 12815 -22629 12849 -22593
rect 12815 -22699 12849 -22663
rect 13073 -22559 13107 -22523
rect 13073 -22629 13107 -22593
rect 13073 -22699 13107 -22663
rect 13331 -22559 13365 -22523
rect 13331 -22629 13365 -22593
rect 13331 -22699 13365 -22663
rect 13589 -22559 13623 -22523
rect 13589 -22629 13623 -22593
rect 13589 -22699 13623 -22663
rect 13847 -22559 13881 -22523
rect 13847 -22629 13881 -22593
rect 13847 -22699 13881 -22663
rect 14446 -22558 14480 -22522
rect 14446 -22628 14480 -22592
rect 14446 -22698 14480 -22662
rect 14704 -22558 14738 -22522
rect 14704 -22628 14738 -22592
rect 14704 -22698 14738 -22662
rect 14962 -22558 14996 -22522
rect 14962 -22628 14996 -22592
rect 14962 -22699 14996 -22663
rect 15220 -22558 15254 -22522
rect 15220 -22628 15254 -22592
rect 15220 -22698 15254 -22662
rect 15478 -22558 15512 -22522
rect 15478 -22628 15512 -22592
rect 15478 -22698 15512 -22662
rect 15736 -22558 15770 -22522
rect 15736 -22628 15770 -22592
rect 15736 -22698 15770 -22662
rect 15994 -22558 16028 -22522
rect 15994 -22628 16028 -22592
rect 15994 -22698 16028 -22662
rect 16252 -22558 16286 -22522
rect 16252 -22628 16286 -22592
rect 16252 -22698 16286 -22662
rect 16510 -22558 16544 -22522
rect 16510 -22628 16544 -22592
rect 16510 -22698 16544 -22662
rect 9113 -22977 9147 -22941
rect 9113 -23047 9147 -23011
rect 9113 -23117 9147 -23081
rect 9371 -22977 9405 -22941
rect 9371 -23047 9405 -23011
rect 9371 -23117 9405 -23081
rect 9629 -22977 9663 -22941
rect 9629 -23047 9663 -23011
rect 9629 -23118 9663 -23082
rect 9887 -22977 9921 -22941
rect 9887 -23047 9921 -23011
rect 9887 -23117 9921 -23081
rect 10145 -22977 10179 -22941
rect 10145 -23047 10179 -23011
rect 10145 -23117 10179 -23081
rect 10403 -22977 10437 -22941
rect 10403 -23047 10437 -23011
rect 10403 -23117 10437 -23081
rect 10661 -22977 10695 -22941
rect 10661 -23047 10695 -23011
rect 10661 -23117 10695 -23081
rect 10919 -22977 10953 -22941
rect 10919 -23047 10953 -23011
rect 10919 -23117 10953 -23081
rect 11177 -22977 11211 -22941
rect 11177 -23047 11211 -23011
rect 11177 -23117 11211 -23081
rect 11783 -22977 11817 -22941
rect 11783 -23047 11817 -23011
rect 11783 -23117 11817 -23081
rect 12041 -22977 12075 -22941
rect 12041 -23047 12075 -23011
rect 12041 -23117 12075 -23081
rect 12299 -22977 12333 -22941
rect 12299 -23047 12333 -23011
rect 12299 -23118 12333 -23082
rect 12557 -22977 12591 -22941
rect 12557 -23047 12591 -23011
rect 12557 -23117 12591 -23081
rect 12815 -22977 12849 -22941
rect 12815 -23047 12849 -23011
rect 12815 -23117 12849 -23081
rect 13073 -22977 13107 -22941
rect 13073 -23047 13107 -23011
rect 13073 -23117 13107 -23081
rect 13331 -22977 13365 -22941
rect 13331 -23047 13365 -23011
rect 13331 -23117 13365 -23081
rect 13589 -22977 13623 -22941
rect 13589 -23047 13623 -23011
rect 13589 -23117 13623 -23081
rect 13847 -22977 13881 -22941
rect 13847 -23047 13881 -23011
rect 13847 -23117 13881 -23081
rect 14446 -22976 14480 -22940
rect 14446 -23046 14480 -23010
rect 14446 -23116 14480 -23080
rect 14704 -22976 14738 -22940
rect 14704 -23046 14738 -23010
rect 14704 -23116 14738 -23080
rect 14962 -22976 14996 -22940
rect 14962 -23046 14996 -23010
rect 14962 -23117 14996 -23081
rect 15220 -22976 15254 -22940
rect 15220 -23046 15254 -23010
rect 15220 -23116 15254 -23080
rect 15478 -22976 15512 -22940
rect 15478 -23046 15512 -23010
rect 15478 -23116 15512 -23080
rect 15736 -22976 15770 -22940
rect 15736 -23046 15770 -23010
rect 15736 -23116 15770 -23080
rect 15994 -22976 16028 -22940
rect 15994 -23046 16028 -23010
rect 15994 -23116 16028 -23080
rect 16252 -22976 16286 -22940
rect 16252 -23046 16286 -23010
rect 16252 -23116 16286 -23080
rect 16510 -22976 16544 -22940
rect 16510 -23046 16544 -23010
rect 16510 -23116 16544 -23080
rect 9113 -23395 9147 -23359
rect 9113 -23465 9147 -23429
rect 9113 -23535 9147 -23499
rect 9371 -23395 9405 -23359
rect 9371 -23465 9405 -23429
rect 9371 -23535 9405 -23499
rect 9629 -23395 9663 -23359
rect 9629 -23465 9663 -23429
rect 9629 -23536 9663 -23500
rect 9887 -23395 9921 -23359
rect 9887 -23465 9921 -23429
rect 9887 -23535 9921 -23499
rect 10145 -23395 10179 -23359
rect 10145 -23465 10179 -23429
rect 10145 -23535 10179 -23499
rect 10403 -23395 10437 -23359
rect 10403 -23465 10437 -23429
rect 10403 -23535 10437 -23499
rect 10661 -23395 10695 -23359
rect 10661 -23465 10695 -23429
rect 10661 -23535 10695 -23499
rect 10919 -23395 10953 -23359
rect 10919 -23465 10953 -23429
rect 10919 -23535 10953 -23499
rect 11177 -23395 11211 -23359
rect 11177 -23465 11211 -23429
rect 11177 -23535 11211 -23499
rect 11783 -23395 11817 -23359
rect 11783 -23465 11817 -23429
rect 11783 -23535 11817 -23499
rect 12041 -23395 12075 -23359
rect 12041 -23465 12075 -23429
rect 12041 -23535 12075 -23499
rect 12299 -23395 12333 -23359
rect 12299 -23465 12333 -23429
rect 12299 -23536 12333 -23500
rect 12557 -23395 12591 -23359
rect 12557 -23465 12591 -23429
rect 12557 -23535 12591 -23499
rect 12815 -23395 12849 -23359
rect 12815 -23465 12849 -23429
rect 12815 -23535 12849 -23499
rect 13073 -23395 13107 -23359
rect 13073 -23465 13107 -23429
rect 13073 -23535 13107 -23499
rect 13331 -23395 13365 -23359
rect 13331 -23465 13365 -23429
rect 13331 -23535 13365 -23499
rect 13589 -23395 13623 -23359
rect 13589 -23465 13623 -23429
rect 13589 -23535 13623 -23499
rect 13847 -23395 13881 -23359
rect 13847 -23465 13881 -23429
rect 13847 -23535 13881 -23499
rect 14446 -23394 14480 -23358
rect 14446 -23464 14480 -23428
rect 14446 -23534 14480 -23498
rect 14704 -23394 14738 -23358
rect 14704 -23464 14738 -23428
rect 14704 -23534 14738 -23498
rect 14962 -23394 14996 -23358
rect 14962 -23464 14996 -23428
rect 14962 -23535 14996 -23499
rect 15220 -23394 15254 -23358
rect 15220 -23464 15254 -23428
rect 15220 -23534 15254 -23498
rect 15478 -23394 15512 -23358
rect 15478 -23464 15512 -23428
rect 15478 -23534 15512 -23498
rect 15736 -23394 15770 -23358
rect 15736 -23464 15770 -23428
rect 15736 -23534 15770 -23498
rect 15994 -23394 16028 -23358
rect 15994 -23464 16028 -23428
rect 15994 -23534 16028 -23498
rect 16252 -23394 16286 -23358
rect 16252 -23464 16286 -23428
rect 16252 -23534 16286 -23498
rect 16510 -23394 16544 -23358
rect 16510 -23464 16544 -23428
rect 16510 -23534 16544 -23498
rect 9113 -23813 9147 -23777
rect 9113 -23883 9147 -23847
rect 9113 -23953 9147 -23917
rect 9371 -23813 9405 -23777
rect 9371 -23883 9405 -23847
rect 9371 -23953 9405 -23917
rect 9629 -23813 9663 -23777
rect 9629 -23883 9663 -23847
rect 9629 -23954 9663 -23918
rect 9887 -23813 9921 -23777
rect 9887 -23883 9921 -23847
rect 9887 -23953 9921 -23917
rect 10145 -23813 10179 -23777
rect 10145 -23883 10179 -23847
rect 10145 -23953 10179 -23917
rect 10403 -23813 10437 -23777
rect 10403 -23883 10437 -23847
rect 10403 -23953 10437 -23917
rect 10661 -23813 10695 -23777
rect 10661 -23883 10695 -23847
rect 10661 -23953 10695 -23917
rect 10919 -23813 10953 -23777
rect 10919 -23883 10953 -23847
rect 10919 -23953 10953 -23917
rect 11177 -23813 11211 -23777
rect 11177 -23883 11211 -23847
rect 11177 -23953 11211 -23917
rect 11783 -23813 11817 -23777
rect 11783 -23883 11817 -23847
rect 11783 -23953 11817 -23917
rect 12041 -23813 12075 -23777
rect 12041 -23883 12075 -23847
rect 12041 -23953 12075 -23917
rect 12299 -23813 12333 -23777
rect 12299 -23883 12333 -23847
rect 12299 -23954 12333 -23918
rect 12557 -23813 12591 -23777
rect 12557 -23883 12591 -23847
rect 12557 -23953 12591 -23917
rect 12815 -23813 12849 -23777
rect 12815 -23883 12849 -23847
rect 12815 -23953 12849 -23917
rect 13073 -23813 13107 -23777
rect 13073 -23883 13107 -23847
rect 13073 -23953 13107 -23917
rect 13331 -23813 13365 -23777
rect 13331 -23883 13365 -23847
rect 13331 -23953 13365 -23917
rect 13589 -23813 13623 -23777
rect 13589 -23883 13623 -23847
rect 13589 -23953 13623 -23917
rect 13847 -23813 13881 -23777
rect 13847 -23883 13881 -23847
rect 13847 -23953 13881 -23917
rect 14446 -23812 14480 -23776
rect 14446 -23882 14480 -23846
rect 14446 -23952 14480 -23916
rect 14704 -23812 14738 -23776
rect 14704 -23882 14738 -23846
rect 14704 -23952 14738 -23916
rect 14962 -23812 14996 -23776
rect 14962 -23882 14996 -23846
rect 14962 -23953 14996 -23917
rect 15220 -23812 15254 -23776
rect 15220 -23882 15254 -23846
rect 15220 -23952 15254 -23916
rect 15478 -23812 15512 -23776
rect 15478 -23882 15512 -23846
rect 15478 -23952 15512 -23916
rect 15736 -23812 15770 -23776
rect 15736 -23882 15770 -23846
rect 15736 -23952 15770 -23916
rect 15994 -23812 16028 -23776
rect 15994 -23882 16028 -23846
rect 15994 -23952 16028 -23916
rect 16252 -23812 16286 -23776
rect 16252 -23882 16286 -23846
rect 16252 -23952 16286 -23916
rect 16510 -23812 16544 -23776
rect 16510 -23882 16544 -23846
rect 16510 -23952 16544 -23916
rect 8993 -24465 9027 -24431
rect 8993 -24535 9027 -24499
rect 8993 -24603 9027 -24569
rect 9251 -24465 9285 -24431
rect 9251 -24535 9285 -24499
rect 9251 -24603 9285 -24569
rect 9533 -24465 9567 -24431
rect 9533 -24535 9567 -24499
rect 9533 -24603 9567 -24569
rect 9791 -24465 9825 -24431
rect 9791 -24535 9825 -24499
rect 9791 -24603 9825 -24569
rect 10013 -24465 10047 -24431
rect 10013 -24535 10047 -24499
rect 10013 -24603 10047 -24569
rect 10271 -24465 10305 -24431
rect 10271 -24535 10305 -24499
rect 10271 -24603 10305 -24569
rect 10516 -24463 10550 -24429
rect 10516 -24533 10550 -24497
rect 10516 -24601 10550 -24567
rect 10774 -24463 10808 -24429
rect 10774 -24533 10808 -24497
rect 10774 -24601 10808 -24567
rect 11026 -24453 11060 -24419
rect 11026 -24523 11060 -24487
rect 11026 -24591 11060 -24557
rect 11284 -24453 11318 -24419
rect 11284 -24523 11318 -24487
rect 11284 -24591 11318 -24557
rect 11663 -24465 11697 -24431
rect 11663 -24535 11697 -24499
rect 11663 -24603 11697 -24569
rect 11921 -24465 11955 -24431
rect 11921 -24535 11955 -24499
rect 11921 -24603 11955 -24569
rect 12203 -24465 12237 -24431
rect 12203 -24535 12237 -24499
rect 12203 -24603 12237 -24569
rect 12461 -24465 12495 -24431
rect 12461 -24535 12495 -24499
rect 12461 -24603 12495 -24569
rect 12683 -24465 12717 -24431
rect 12683 -24535 12717 -24499
rect 12683 -24603 12717 -24569
rect 12941 -24465 12975 -24431
rect 12941 -24535 12975 -24499
rect 12941 -24603 12975 -24569
rect 13186 -24463 13220 -24429
rect 13186 -24533 13220 -24497
rect 13186 -24601 13220 -24567
rect 13444 -24463 13478 -24429
rect 13444 -24533 13478 -24497
rect 13444 -24601 13478 -24567
rect 13696 -24453 13730 -24419
rect 13696 -24523 13730 -24487
rect 13696 -24591 13730 -24557
rect 13954 -24453 13988 -24419
rect 13954 -24523 13988 -24487
rect 13954 -24591 13988 -24557
rect 14326 -24464 14360 -24430
rect 14326 -24534 14360 -24498
rect 14326 -24602 14360 -24568
rect 14584 -24464 14618 -24430
rect 14584 -24534 14618 -24498
rect 14584 -24602 14618 -24568
rect 14866 -24464 14900 -24430
rect 14866 -24534 14900 -24498
rect 14866 -24602 14900 -24568
rect 15124 -24464 15158 -24430
rect 15124 -24534 15158 -24498
rect 15124 -24602 15158 -24568
rect 15346 -24464 15380 -24430
rect 15346 -24534 15380 -24498
rect 15346 -24602 15380 -24568
rect 15604 -24464 15638 -24430
rect 15604 -24534 15638 -24498
rect 15604 -24602 15638 -24568
rect 15849 -24462 15883 -24428
rect 15849 -24532 15883 -24496
rect 15849 -24600 15883 -24566
rect 16107 -24462 16141 -24428
rect 16107 -24532 16141 -24496
rect 16107 -24600 16141 -24566
rect 16359 -24452 16393 -24418
rect 16359 -24522 16393 -24486
rect 16359 -24590 16393 -24556
rect 16617 -24452 16651 -24418
rect 16617 -24522 16651 -24486
rect 16617 -24590 16651 -24556
rect 17990 -9010 18024 -7634
rect 19648 -9010 19682 -7634
rect 21306 -9010 21340 -7634
rect 17990 -10520 18024 -9144
rect 19648 -10520 19682 -9144
rect 21306 -10520 21340 -9144
rect 17990 -12030 18024 -10654
rect 19648 -12030 19682 -10654
rect 21306 -12030 21340 -10654
rect 17990 -13540 18024 -12164
rect 19648 -13540 19682 -12164
rect 21306 -13540 21340 -12164
rect 17990 -15050 18024 -13674
rect 19648 -15050 19682 -13674
rect 21306 -15050 21340 -13674
rect 17990 -16560 18024 -15184
rect 19648 -16560 19682 -15184
rect 21306 -16560 21340 -15184
rect 17990 -18070 18024 -16694
rect 19648 -18070 19682 -16694
rect 21306 -18070 21340 -16694
rect 17990 -19580 18024 -18204
rect 19648 -19580 19682 -18204
rect 21306 -19580 21340 -18204
rect 17990 -21090 18024 -19714
rect 19648 -21090 19682 -19714
rect 21306 -21090 21340 -19714
rect 17990 -22600 18024 -21224
rect 19648 -22600 19682 -21224
rect 21306 -22600 21340 -21224
rect 17990 -24110 18024 -22734
rect 19648 -24110 19682 -22734
rect 21306 -24110 21340 -22734
rect 17990 -25620 18024 -24244
rect 19648 -25620 19682 -24244
rect 21306 -25620 21340 -24244
<< pdiffc >>
rect -94610 19524 -94576 20212
rect -92952 19524 -92918 20212
rect -91294 19524 -91260 20212
rect -89636 19524 -89602 20212
rect -87978 19524 -87944 20212
rect -86320 19524 -86286 20212
rect -84662 19524 -84628 20212
rect -83004 19524 -82970 20212
rect -81346 19524 -81312 20212
rect -79688 19524 -79654 20212
rect -78030 19524 -77996 20212
rect -76372 19524 -76338 20212
rect -74714 19524 -74680 20212
rect -73056 19524 -73022 20212
rect -71398 19524 -71364 20212
rect -69740 19524 -69706 20212
rect -68082 19524 -68048 20212
rect -66424 19524 -66390 20212
rect -64766 19524 -64732 20212
rect -63108 19524 -63074 20212
rect -61450 19524 -61416 20212
rect -59792 19524 -59758 20212
rect -58134 19524 -58100 20212
rect -56476 19524 -56442 20212
rect -54818 19524 -54784 20212
rect -53160 19524 -53126 20212
rect -51502 19524 -51468 20212
rect -49844 19524 -49810 20212
rect -48186 19524 -48152 20212
rect -46528 19524 -46494 20212
rect -44870 19524 -44836 20212
rect -43212 19524 -43178 20212
rect -41554 19524 -41520 20212
rect -39896 19524 -39862 20212
rect -38238 19524 -38204 20212
rect -36580 19524 -36546 20212
rect -34922 19524 -34888 20212
rect -33264 19524 -33230 20212
rect -31606 19524 -31572 20212
rect -29948 19524 -29914 20212
rect -28290 19524 -28256 20212
rect -94610 17888 -94576 18576
rect -92952 17888 -92918 18576
rect -91294 17888 -91260 18576
rect -89636 17888 -89602 18576
rect -87978 17888 -87944 18576
rect -86320 17888 -86286 18576
rect -84662 17888 -84628 18576
rect -83004 17888 -82970 18576
rect -81346 17888 -81312 18576
rect -79688 17888 -79654 18576
rect -78030 17888 -77996 18576
rect -76372 17888 -76338 18576
rect -74714 17888 -74680 18576
rect -73056 17888 -73022 18576
rect -71398 17888 -71364 18576
rect -69740 17888 -69706 18576
rect -68082 17888 -68048 18576
rect -66424 17888 -66390 18576
rect -64766 17888 -64732 18576
rect -63108 17888 -63074 18576
rect -61450 17888 -61416 18576
rect -59792 17888 -59758 18576
rect -58134 17888 -58100 18576
rect -56476 17888 -56442 18576
rect -54818 17888 -54784 18576
rect -53160 17888 -53126 18576
rect -51502 17888 -51468 18576
rect -49844 17888 -49810 18576
rect -48186 17888 -48152 18576
rect -46528 17888 -46494 18576
rect -44870 17888 -44836 18576
rect -43212 17888 -43178 18576
rect -41554 17888 -41520 18576
rect -39896 17888 -39862 18576
rect -38238 17888 -38204 18576
rect -36580 17888 -36546 18576
rect -34922 17888 -34888 18576
rect -33264 17888 -33230 18576
rect -31606 17888 -31572 18576
rect -29948 17888 -29914 18576
rect -28290 17888 -28256 18576
rect -94608 16142 -94574 16830
rect -92950 16142 -92916 16830
rect -91292 16142 -91258 16830
rect -89634 16142 -89600 16830
rect -87976 16142 -87942 16830
rect -86318 16142 -86284 16830
rect -84660 16142 -84626 16830
rect -83002 16142 -82968 16830
rect -81344 16142 -81310 16830
rect -79686 16142 -79652 16830
rect -78028 16142 -77994 16830
rect -76370 16142 -76336 16830
rect -74712 16142 -74678 16830
rect -73054 16142 -73020 16830
rect -71396 16142 -71362 16830
rect -69738 16142 -69704 16830
rect -68080 16142 -68046 16830
rect -66422 16142 -66388 16830
rect -64764 16142 -64730 16830
rect -63106 16142 -63072 16830
rect -61448 16142 -61414 16830
rect -59790 16142 -59756 16830
rect -58132 16142 -58098 16830
rect -56474 16142 -56440 16830
rect -54816 16142 -54782 16830
rect -53158 16142 -53124 16830
rect -51500 16142 -51466 16830
rect -49842 16142 -49808 16830
rect -48184 16142 -48150 16830
rect -46526 16142 -46492 16830
rect -44868 16142 -44834 16830
rect -43210 16142 -43176 16830
rect -41552 16142 -41518 16830
rect -39894 16142 -39860 16830
rect -38236 16142 -38202 16830
rect -36578 16142 -36544 16830
rect -34920 16142 -34886 16830
rect -33262 16142 -33228 16830
rect -31604 16142 -31570 16830
rect -29946 16142 -29912 16830
rect -28288 16142 -28254 16830
rect -94608 14506 -94574 15194
rect -92950 14506 -92916 15194
rect -91292 14506 -91258 15194
rect -89634 14506 -89600 15194
rect -87976 14506 -87942 15194
rect -86318 14506 -86284 15194
rect -84660 14506 -84626 15194
rect -83002 14506 -82968 15194
rect -81344 14506 -81310 15194
rect -79686 14506 -79652 15194
rect -78028 14506 -77994 15194
rect -76370 14506 -76336 15194
rect -74712 14506 -74678 15194
rect -73054 14506 -73020 15194
rect -71396 14506 -71362 15194
rect -69738 14506 -69704 15194
rect -68080 14506 -68046 15194
rect -66422 14506 -66388 15194
rect -64764 14506 -64730 15194
rect -63106 14506 -63072 15194
rect -61448 14506 -61414 15194
rect -59790 14506 -59756 15194
rect -58132 14506 -58098 15194
rect -56474 14506 -56440 15194
rect -54816 14506 -54782 15194
rect -53158 14506 -53124 15194
rect -51500 14506 -51466 15194
rect -49842 14506 -49808 15194
rect -48184 14506 -48150 15194
rect -46526 14506 -46492 15194
rect -44868 14506 -44834 15194
rect -43210 14506 -43176 15194
rect -41552 14506 -41518 15194
rect -39894 14506 -39860 15194
rect -38236 14506 -38202 15194
rect -36578 14506 -36544 15194
rect -34920 14506 -34886 15194
rect -33262 14506 -33228 15194
rect -31604 14506 -31570 15194
rect -29946 14506 -29912 15194
rect -28288 14506 -28254 15194
rect -94608 12870 -94574 13558
rect -92950 12870 -92916 13558
rect -91292 12870 -91258 13558
rect -89634 12870 -89600 13558
rect -87976 12870 -87942 13558
rect -86318 12870 -86284 13558
rect -84660 12870 -84626 13558
rect -83002 12870 -82968 13558
rect -81344 12870 -81310 13558
rect -79686 12870 -79652 13558
rect -78028 12870 -77994 13558
rect -76370 12870 -76336 13558
rect -74712 12870 -74678 13558
rect -73054 12870 -73020 13558
rect -71396 12870 -71362 13558
rect -69738 12870 -69704 13558
rect -68080 12870 -68046 13558
rect -66422 12870 -66388 13558
rect -64764 12870 -64730 13558
rect -63106 12870 -63072 13558
rect -61448 12870 -61414 13558
rect -59790 12870 -59756 13558
rect -58132 12870 -58098 13558
rect -56474 12870 -56440 13558
rect -54816 12870 -54782 13558
rect -53158 12870 -53124 13558
rect -51500 12870 -51466 13558
rect -49842 12870 -49808 13558
rect -48184 12870 -48150 13558
rect -46526 12870 -46492 13558
rect -44868 12870 -44834 13558
rect -43210 12870 -43176 13558
rect -41552 12870 -41518 13558
rect -39894 12870 -39860 13558
rect -38236 12870 -38202 13558
rect -36578 12870 -36544 13558
rect -34920 12870 -34886 13558
rect -33262 12870 -33228 13558
rect -31604 12870 -31570 13558
rect -29946 12870 -29912 13558
rect -28288 12870 -28254 13558
rect -94608 11234 -94574 11922
rect -92950 11234 -92916 11922
rect -91292 11234 -91258 11922
rect -89634 11234 -89600 11922
rect -87976 11234 -87942 11922
rect -86318 11234 -86284 11922
rect -84660 11234 -84626 11922
rect -83002 11234 -82968 11922
rect -81344 11234 -81310 11922
rect -79686 11234 -79652 11922
rect -78028 11234 -77994 11922
rect -76370 11234 -76336 11922
rect -74712 11234 -74678 11922
rect -73054 11234 -73020 11922
rect -71396 11234 -71362 11922
rect -69738 11234 -69704 11922
rect -68080 11234 -68046 11922
rect -66422 11234 -66388 11922
rect -64764 11234 -64730 11922
rect -63106 11234 -63072 11922
rect -61448 11234 -61414 11922
rect -59790 11234 -59756 11922
rect -58132 11234 -58098 11922
rect -56474 11234 -56440 11922
rect -54816 11234 -54782 11922
rect -53158 11234 -53124 11922
rect -51500 11234 -51466 11922
rect -49842 11234 -49808 11922
rect -48184 11234 -48150 11922
rect -46526 11234 -46492 11922
rect -44868 11234 -44834 11922
rect -43210 11234 -43176 11922
rect -41552 11234 -41518 11922
rect -39894 11234 -39860 11922
rect -38236 11234 -38202 11922
rect -36578 11234 -36544 11922
rect -34920 11234 -34886 11922
rect -33262 11234 -33228 11922
rect -31604 11234 -31570 11922
rect -29946 11234 -29912 11922
rect -28288 11234 -28254 11922
rect -94608 9596 -94574 10284
rect -92950 9596 -92916 10284
rect -91292 9596 -91258 10284
rect -89634 9596 -89600 10284
rect -87976 9596 -87942 10284
rect -86318 9596 -86284 10284
rect -84660 9596 -84626 10284
rect -83002 9596 -82968 10284
rect -81344 9596 -81310 10284
rect -79686 9596 -79652 10284
rect -78028 9596 -77994 10284
rect -76370 9596 -76336 10284
rect -74712 9596 -74678 10284
rect -73054 9596 -73020 10284
rect -71396 9596 -71362 10284
rect -69738 9596 -69704 10284
rect -68080 9596 -68046 10284
rect -66422 9596 -66388 10284
rect -64764 9596 -64730 10284
rect -63106 9596 -63072 10284
rect -61448 9596 -61414 10284
rect -59790 9596 -59756 10284
rect -58132 9596 -58098 10284
rect -56474 9596 -56440 10284
rect -54816 9596 -54782 10284
rect -53158 9596 -53124 10284
rect -51500 9596 -51466 10284
rect -49842 9596 -49808 10284
rect -48184 9596 -48150 10284
rect -46526 9596 -46492 10284
rect -44868 9596 -44834 10284
rect -43210 9596 -43176 10284
rect -41552 9596 -41518 10284
rect -39894 9596 -39860 10284
rect -38236 9596 -38202 10284
rect -36578 9596 -36544 10284
rect -34920 9596 -34886 10284
rect -33262 9596 -33228 10284
rect -31604 9596 -31570 10284
rect -29946 9596 -29912 10284
rect -28288 9596 -28254 10284
rect -94608 7960 -94574 8648
rect -92950 7960 -92916 8648
rect -91292 7960 -91258 8648
rect -89634 7960 -89600 8648
rect -87976 7960 -87942 8648
rect -86318 7960 -86284 8648
rect -84660 7960 -84626 8648
rect -83002 7960 -82968 8648
rect -81344 7960 -81310 8648
rect -79686 7960 -79652 8648
rect -78028 7960 -77994 8648
rect -76370 7960 -76336 8648
rect -74712 7960 -74678 8648
rect -73054 7960 -73020 8648
rect -71396 7960 -71362 8648
rect -69738 7960 -69704 8648
rect -68080 7960 -68046 8648
rect -66422 7960 -66388 8648
rect -64764 7960 -64730 8648
rect -63106 7960 -63072 8648
rect -61448 7960 -61414 8648
rect -59790 7960 -59756 8648
rect -58132 7960 -58098 8648
rect -56474 7960 -56440 8648
rect -54816 7960 -54782 8648
rect -53158 7960 -53124 8648
rect -51500 7960 -51466 8648
rect -49842 7960 -49808 8648
rect -48184 7960 -48150 8648
rect -46526 7960 -46492 8648
rect -44868 7960 -44834 8648
rect -43210 7960 -43176 8648
rect -41552 7960 -41518 8648
rect -39894 7960 -39860 8648
rect -38236 7960 -38202 8648
rect -36578 7960 -36544 8648
rect -34920 7960 -34886 8648
rect -33262 7960 -33228 8648
rect -31604 7960 -31570 8648
rect -29946 7960 -29912 8648
rect -28288 7960 -28254 8648
rect -94608 6324 -94574 7012
rect -92950 6324 -92916 7012
rect -91292 6324 -91258 7012
rect -89634 6324 -89600 7012
rect -87976 6324 -87942 7012
rect -86318 6324 -86284 7012
rect -84660 6324 -84626 7012
rect -83002 6324 -82968 7012
rect -81344 6324 -81310 7012
rect -79686 6324 -79652 7012
rect -78028 6324 -77994 7012
rect -76370 6324 -76336 7012
rect -74712 6324 -74678 7012
rect -73054 6324 -73020 7012
rect -71396 6324 -71362 7012
rect -69738 6324 -69704 7012
rect -68080 6324 -68046 7012
rect -66422 6324 -66388 7012
rect -64764 6324 -64730 7012
rect -63106 6324 -63072 7012
rect -61448 6324 -61414 7012
rect -59790 6324 -59756 7012
rect -58132 6324 -58098 7012
rect -56474 6324 -56440 7012
rect -54816 6324 -54782 7012
rect -53158 6324 -53124 7012
rect -51500 6324 -51466 7012
rect -49842 6324 -49808 7012
rect -48184 6324 -48150 7012
rect -46526 6324 -46492 7012
rect -44868 6324 -44834 7012
rect -43210 6324 -43176 7012
rect -41552 6324 -41518 7012
rect -39894 6324 -39860 7012
rect -38236 6324 -38202 7012
rect -36578 6324 -36544 7012
rect -34920 6324 -34886 7012
rect -33262 6324 -33228 7012
rect -31604 6324 -31570 7012
rect -29946 6324 -29912 7012
rect -28288 6324 -28254 7012
rect -94608 4688 -94574 5376
rect -92950 4688 -92916 5376
rect -91292 4688 -91258 5376
rect -89634 4688 -89600 5376
rect -87976 4688 -87942 5376
rect -86318 4688 -86284 5376
rect -84660 4688 -84626 5376
rect -83002 4688 -82968 5376
rect -81344 4688 -81310 5376
rect -79686 4688 -79652 5376
rect -78028 4688 -77994 5376
rect -76370 4688 -76336 5376
rect -74712 4688 -74678 5376
rect -73054 4688 -73020 5376
rect -71396 4688 -71362 5376
rect -69738 4688 -69704 5376
rect -68080 4688 -68046 5376
rect -66422 4688 -66388 5376
rect -64764 4688 -64730 5376
rect -63106 4688 -63072 5376
rect -61448 4688 -61414 5376
rect -59790 4688 -59756 5376
rect -58132 4688 -58098 5376
rect -56474 4688 -56440 5376
rect -54816 4688 -54782 5376
rect -53158 4688 -53124 5376
rect -51500 4688 -51466 5376
rect -49842 4688 -49808 5376
rect -48184 4688 -48150 5376
rect -46526 4688 -46492 5376
rect -44868 4688 -44834 5376
rect -43210 4688 -43176 5376
rect -41552 4688 -41518 5376
rect -39894 4688 -39860 5376
rect -38236 4688 -38202 5376
rect -36578 4688 -36544 5376
rect -34920 4688 -34886 5376
rect -33262 4688 -33228 5376
rect -31604 4688 -31570 5376
rect -29946 4688 -29912 5376
rect -28288 4688 -28254 5376
rect -61770 3596 -61736 3784
rect -61674 3596 -61640 3784
rect -61578 3596 -61544 3784
rect -61482 3596 -61448 3784
rect 2620 5172 2654 5660
rect 1074 4744 1108 4932
rect 1162 4744 1196 4932
rect 1306 4742 1340 4930
rect 1394 4742 1428 4930
rect 1534 4740 1568 4928
rect 1622 4740 1656 4928
rect 1752 4742 1786 4930
rect 1840 4742 1874 4930
rect 2878 5172 2912 5660
rect 3276 5180 3310 5668
rect 3534 5180 3568 5668
rect 3792 5180 3826 5668
rect 4276 5180 4310 5668
rect 4534 5180 4568 5668
rect 4792 5180 4826 5668
rect 5182 5184 5216 5672
rect 5440 5184 5474 5672
rect 6260 4762 6294 4950
rect 6348 4762 6382 4950
rect 6492 4760 6526 4948
rect 6580 4760 6614 4948
rect 6720 4758 6754 4946
rect 6808 4758 6842 4946
rect 6938 4760 6972 4948
rect 7026 4760 7060 4948
rect 8556 4912 8590 5400
rect 8814 4912 8848 5400
rect 9035 4904 9069 5392
rect 9293 4904 9327 5392
rect 9551 4904 9585 5392
rect 9693 4906 9727 5394
rect 9951 5040 9985 5394
rect 10209 4906 10243 5394
rect 10350 4886 10384 5374
rect 10608 4886 10642 5374
rect 11436 4774 11470 4962
rect 11524 4774 11558 4962
rect 11668 4772 11702 4960
rect 11756 4772 11790 4960
rect 11896 4770 11930 4958
rect 11984 4770 12018 4958
rect 12114 4772 12148 4960
rect 12202 4772 12236 4960
rect 13830 4784 13864 5272
rect 14088 4784 14122 5272
rect 14224 4766 14258 5254
rect 14682 4766 14716 5254
rect 14796 4766 14830 5254
rect 15254 4766 15288 5254
rect 15418 4796 15452 5284
rect 15676 4796 15710 5284
rect 17092 4566 17126 4754
rect 17180 4566 17214 4754
rect 17324 4564 17358 4752
rect 17412 4564 17446 4752
rect 17552 4562 17586 4750
rect 17640 4562 17674 4750
rect 17770 4564 17804 4752
rect 17858 4564 17892 4752
rect -61386 3596 -61352 3784
rect 26886 2482 26920 2794
rect 26974 2482 27008 2794
rect 27090 2520 27124 2832
rect 27178 2520 27212 2832
rect 27498 2490 27532 2802
rect 27586 2490 27620 2802
rect 27702 2528 27736 2840
rect 27790 2528 27824 2840
rect 28076 2486 28110 2798
rect 28164 2486 28198 2798
rect 28280 2524 28314 2836
rect 28368 2524 28402 2836
rect 28650 2494 28684 2806
rect 28738 2494 28772 2806
rect 28854 2532 28888 2844
rect 28942 2532 28976 2844
rect 29228 2494 29262 2806
rect 29316 2494 29350 2806
rect 29432 2532 29466 2844
rect 29520 2532 29554 2844
rect 29806 2494 29840 2806
rect 29894 2494 29928 2806
rect 30010 2532 30044 2844
rect 30098 2532 30132 2844
rect 30388 2498 30422 2810
rect 30476 2498 30510 2810
rect 30592 2536 30626 2848
rect 30680 2536 30714 2848
rect 30964 2494 30998 2806
rect 31052 2494 31086 2806
rect 31168 2532 31202 2844
rect 31256 2532 31290 2844
rect 31534 2490 31568 2802
rect 31622 2490 31656 2802
rect 31738 2528 31772 2840
rect 31826 2528 31860 2840
rect 28280 428 28314 740
rect 28368 428 28402 740
rect 28480 466 28514 778
rect 28568 466 28602 778
rect 28682 426 28716 738
rect 28770 426 28804 738
rect 28280 -78 28314 234
rect 28368 -78 28402 234
rect 28480 -40 28514 272
rect 28568 -40 28602 272
rect 28680 -78 28714 234
rect 28768 -78 28802 234
rect 28280 -586 28314 -274
rect 28368 -586 28402 -274
rect 28480 -548 28514 -236
rect 28568 -548 28602 -236
rect 28680 -586 28714 -274
rect 28768 -586 28802 -274
rect 8769 -1076 8803 -1042
rect 8769 -1144 8803 -1110
rect 8853 -1092 8887 -1058
rect 8937 -1076 8971 -1042
rect 9120 -1068 9154 -1034
rect 9204 -1076 9238 -1042
rect 9297 -1070 9331 -1036
rect 9451 -1094 9485 -1060
rect 9548 -1078 9582 -1044
rect 9632 -1094 9666 -1060
rect 9745 -1068 9779 -1034
rect 8937 -1144 8971 -1110
rect 9833 -1076 9867 -1042
rect 9930 -1069 9964 -1035
rect 10122 -1068 10156 -1034
rect 10206 -1094 10240 -1060
rect 10292 -1068 10326 -1034
rect 10370 -1068 10404 -1034
rect 10454 -1076 10488 -1042
rect 10454 -1144 10488 -1110
rect 10589 -1068 10623 -1034
rect 10589 -1136 10623 -1102
rect 10686 -1068 10720 -1034
rect 10686 -1136 10720 -1102
rect 10454 -1212 10488 -1178
rect 10686 -1204 10720 -1170
rect 10770 -1104 10804 -1070
rect 10770 -1172 10804 -1138
rect 11235 -1076 11269 -1042
rect 11235 -1144 11269 -1110
rect 11319 -1092 11353 -1058
rect 11403 -1076 11437 -1042
rect 11586 -1068 11620 -1034
rect 11670 -1076 11704 -1042
rect 11763 -1070 11797 -1036
rect 11917 -1094 11951 -1060
rect 12014 -1078 12048 -1044
rect 12098 -1094 12132 -1060
rect 12211 -1068 12245 -1034
rect 11403 -1144 11437 -1110
rect 12299 -1076 12333 -1042
rect 12396 -1069 12430 -1035
rect 12588 -1068 12622 -1034
rect 12672 -1094 12706 -1060
rect 12758 -1068 12792 -1034
rect 12836 -1068 12870 -1034
rect 12920 -1076 12954 -1042
rect 12920 -1144 12954 -1110
rect 13055 -1068 13089 -1034
rect 13055 -1136 13089 -1102
rect 13152 -1068 13186 -1034
rect 13152 -1136 13186 -1102
rect 12920 -1212 12954 -1178
rect 13152 -1204 13186 -1170
rect 13236 -1104 13270 -1070
rect 13236 -1172 13270 -1138
rect 10189 -1870 10223 -1836
rect 10189 -1938 10223 -1904
rect 10189 -2006 10223 -1972
rect 10273 -1870 10307 -1836
rect 10273 -1938 10307 -1904
rect 10273 -2006 10307 -1972
rect 10357 -1870 10391 -1836
rect 10357 -1938 10391 -1904
rect 11235 -1878 11269 -1844
rect 11235 -1946 11269 -1912
rect 11319 -1894 11353 -1860
rect 11403 -1878 11437 -1844
rect 11586 -1870 11620 -1836
rect 11670 -1878 11704 -1844
rect 11763 -1872 11797 -1838
rect 11917 -1896 11951 -1862
rect 12014 -1880 12048 -1846
rect 12098 -1896 12132 -1862
rect 12211 -1870 12245 -1836
rect 11403 -1946 11437 -1912
rect 10357 -2006 10391 -1972
rect 12299 -1878 12333 -1844
rect 12396 -1871 12430 -1837
rect 12588 -1870 12622 -1836
rect 12672 -1896 12706 -1862
rect 12758 -1870 12792 -1836
rect 12836 -1870 12870 -1836
rect 12920 -1878 12954 -1844
rect 12920 -1946 12954 -1912
rect 13055 -1870 13089 -1836
rect 13055 -1938 13089 -1904
rect 13152 -1870 13186 -1836
rect 13152 -1938 13186 -1904
rect 12920 -2014 12954 -1980
rect 13152 -2006 13186 -1972
rect 13236 -1906 13270 -1872
rect 13236 -1974 13270 -1940
rect -9123 -4346 -9089 -4312
rect -9123 -4414 -9089 -4380
rect -9039 -4362 -9005 -4328
rect -8955 -4346 -8921 -4312
rect -8772 -4338 -8738 -4304
rect -8688 -4346 -8654 -4312
rect -8595 -4340 -8561 -4306
rect -8441 -4364 -8407 -4330
rect -8344 -4348 -8310 -4314
rect -8260 -4364 -8226 -4330
rect -8147 -4338 -8113 -4304
rect -8955 -4414 -8921 -4380
rect -8059 -4346 -8025 -4312
rect -7962 -4339 -7928 -4305
rect -7770 -4338 -7736 -4304
rect -7686 -4364 -7652 -4330
rect -7600 -4338 -7566 -4304
rect -7522 -4338 -7488 -4304
rect -7438 -4346 -7404 -4312
rect -7438 -4414 -7404 -4380
rect -7303 -4338 -7269 -4304
rect -7303 -4406 -7269 -4372
rect -7206 -4338 -7172 -4304
rect -7206 -4406 -7172 -4372
rect -7438 -4482 -7404 -4448
rect -7206 -4474 -7172 -4440
rect -7122 -4374 -7088 -4340
rect -7122 -4442 -7088 -4408
rect -7007 -4346 -6973 -4312
rect -7007 -4414 -6973 -4380
rect -6923 -4362 -6889 -4328
rect -6839 -4346 -6805 -4312
rect -6656 -4338 -6622 -4304
rect -6572 -4346 -6538 -4312
rect -6479 -4340 -6445 -4306
rect -6325 -4364 -6291 -4330
rect -6228 -4348 -6194 -4314
rect -6144 -4364 -6110 -4330
rect -6031 -4338 -5997 -4304
rect -6839 -4414 -6805 -4380
rect -5943 -4346 -5909 -4312
rect -5846 -4339 -5812 -4305
rect -5654 -4338 -5620 -4304
rect -5570 -4364 -5536 -4330
rect -5484 -4338 -5450 -4304
rect -5406 -4338 -5372 -4304
rect -5322 -4346 -5288 -4312
rect -5322 -4414 -5288 -4380
rect -5187 -4338 -5153 -4304
rect -5187 -4406 -5153 -4372
rect -5090 -4338 -5056 -4304
rect -5090 -4406 -5056 -4372
rect -5322 -4482 -5288 -4448
rect -5090 -4474 -5056 -4440
rect -5006 -4374 -4972 -4340
rect -5006 -4442 -4972 -4408
rect -4891 -4346 -4857 -4312
rect -4891 -4414 -4857 -4380
rect -4807 -4362 -4773 -4328
rect -4723 -4346 -4689 -4312
rect -4540 -4338 -4506 -4304
rect -4456 -4346 -4422 -4312
rect -4363 -4340 -4329 -4306
rect -4209 -4364 -4175 -4330
rect -4112 -4348 -4078 -4314
rect -4028 -4364 -3994 -4330
rect -3915 -4338 -3881 -4304
rect -4723 -4414 -4689 -4380
rect -3827 -4346 -3793 -4312
rect -3730 -4339 -3696 -4305
rect -3538 -4338 -3504 -4304
rect -3454 -4364 -3420 -4330
rect -3368 -4338 -3334 -4304
rect -3290 -4338 -3256 -4304
rect -3206 -4346 -3172 -4312
rect -3206 -4414 -3172 -4380
rect -3071 -4338 -3037 -4304
rect -3071 -4406 -3037 -4372
rect -2974 -4338 -2940 -4304
rect -2974 -4406 -2940 -4372
rect -3206 -4482 -3172 -4448
rect -2974 -4474 -2940 -4440
rect -2890 -4374 -2856 -4340
rect -2890 -4442 -2856 -4408
rect -2775 -4346 -2741 -4312
rect -2775 -4414 -2741 -4380
rect -2691 -4362 -2657 -4328
rect -2607 -4346 -2573 -4312
rect -2424 -4338 -2390 -4304
rect -2340 -4346 -2306 -4312
rect -2247 -4340 -2213 -4306
rect -2093 -4364 -2059 -4330
rect -1996 -4348 -1962 -4314
rect -1912 -4364 -1878 -4330
rect -1799 -4338 -1765 -4304
rect -2607 -4414 -2573 -4380
rect -1711 -4346 -1677 -4312
rect -1614 -4339 -1580 -4305
rect -1422 -4338 -1388 -4304
rect -1338 -4364 -1304 -4330
rect -1252 -4338 -1218 -4304
rect -1174 -4338 -1140 -4304
rect -1090 -4346 -1056 -4312
rect -1090 -4414 -1056 -4380
rect -955 -4338 -921 -4304
rect -955 -4406 -921 -4372
rect -858 -4338 -824 -4304
rect -858 -4406 -824 -4372
rect -1090 -4482 -1056 -4448
rect -858 -4474 -824 -4440
rect -774 -4374 -740 -4340
rect -774 -4442 -740 -4408
rect -659 -4346 -625 -4312
rect -659 -4414 -625 -4380
rect -575 -4362 -541 -4328
rect -491 -4346 -457 -4312
rect -308 -4338 -274 -4304
rect -224 -4346 -190 -4312
rect -131 -4340 -97 -4306
rect 23 -4364 57 -4330
rect 120 -4348 154 -4314
rect 204 -4364 238 -4330
rect 317 -4338 351 -4304
rect -491 -4414 -457 -4380
rect 405 -4346 439 -4312
rect 502 -4339 536 -4305
rect 694 -4338 728 -4304
rect 778 -4364 812 -4330
rect 864 -4338 898 -4304
rect 942 -4338 976 -4304
rect 1026 -4346 1060 -4312
rect 1026 -4414 1060 -4380
rect 1161 -4338 1195 -4304
rect 1161 -4406 1195 -4372
rect 1258 -4338 1292 -4304
rect 1258 -4406 1292 -4372
rect 1026 -4482 1060 -4448
rect 1258 -4474 1292 -4440
rect 1342 -4374 1376 -4340
rect 1342 -4442 1376 -4408
rect 1457 -4346 1491 -4312
rect 1457 -4414 1491 -4380
rect 1541 -4362 1575 -4328
rect 1625 -4346 1659 -4312
rect 1808 -4338 1842 -4304
rect 1892 -4346 1926 -4312
rect 1985 -4340 2019 -4306
rect 2139 -4364 2173 -4330
rect 2236 -4348 2270 -4314
rect 2320 -4364 2354 -4330
rect 2433 -4338 2467 -4304
rect 1625 -4414 1659 -4380
rect 2521 -4346 2555 -4312
rect 2618 -4339 2652 -4305
rect 2810 -4338 2844 -4304
rect 2894 -4364 2928 -4330
rect 2980 -4338 3014 -4304
rect 3058 -4338 3092 -4304
rect 3142 -4346 3176 -4312
rect 3142 -4414 3176 -4380
rect 3277 -4338 3311 -4304
rect 3277 -4406 3311 -4372
rect 3374 -4338 3408 -4304
rect 3374 -4406 3408 -4372
rect 3142 -4482 3176 -4448
rect 3374 -4474 3408 -4440
rect 3458 -4374 3492 -4340
rect 3458 -4442 3492 -4408
rect 3573 -4346 3607 -4312
rect 3573 -4414 3607 -4380
rect 3657 -4362 3691 -4328
rect 3741 -4346 3775 -4312
rect 3924 -4338 3958 -4304
rect 4008 -4346 4042 -4312
rect 4101 -4340 4135 -4306
rect 4255 -4364 4289 -4330
rect 4352 -4348 4386 -4314
rect 4436 -4364 4470 -4330
rect 4549 -4338 4583 -4304
rect 3741 -4414 3775 -4380
rect 4637 -4346 4671 -4312
rect 4734 -4339 4768 -4305
rect 4926 -4338 4960 -4304
rect 5010 -4364 5044 -4330
rect 5096 -4338 5130 -4304
rect 5174 -4338 5208 -4304
rect 5258 -4346 5292 -4312
rect 5258 -4414 5292 -4380
rect 5393 -4338 5427 -4304
rect 5393 -4406 5427 -4372
rect 5490 -4338 5524 -4304
rect 5490 -4406 5524 -4372
rect 5258 -4482 5292 -4448
rect 5490 -4474 5524 -4440
rect 5574 -4374 5608 -4340
rect 5574 -4442 5608 -4408
rect 5689 -4346 5723 -4312
rect 5689 -4414 5723 -4380
rect 5773 -4362 5807 -4328
rect 5857 -4346 5891 -4312
rect 6040 -4338 6074 -4304
rect 6124 -4346 6158 -4312
rect 6217 -4340 6251 -4306
rect 6371 -4364 6405 -4330
rect 6468 -4348 6502 -4314
rect 6552 -4364 6586 -4330
rect 6665 -4338 6699 -4304
rect 5857 -4414 5891 -4380
rect 6753 -4346 6787 -4312
rect 6850 -4339 6884 -4305
rect 7042 -4338 7076 -4304
rect 7126 -4364 7160 -4330
rect 7212 -4338 7246 -4304
rect 7290 -4338 7324 -4304
rect 7374 -4346 7408 -4312
rect 7374 -4414 7408 -4380
rect 7509 -4338 7543 -4304
rect 7509 -4406 7543 -4372
rect 7606 -4338 7640 -4304
rect 7606 -4406 7640 -4372
rect 7374 -4482 7408 -4448
rect 7606 -4474 7640 -4440
rect 7690 -4374 7724 -4340
rect 7690 -4442 7724 -4408
rect 7805 -4346 7839 -4312
rect 7805 -4414 7839 -4380
rect 7889 -4362 7923 -4328
rect 7973 -4346 8007 -4312
rect 8156 -4338 8190 -4304
rect 8240 -4346 8274 -4312
rect 8333 -4340 8367 -4306
rect 8487 -4364 8521 -4330
rect 8584 -4348 8618 -4314
rect 8668 -4364 8702 -4330
rect 8781 -4338 8815 -4304
rect 7973 -4414 8007 -4380
rect 8869 -4346 8903 -4312
rect 8966 -4339 9000 -4305
rect 9158 -4338 9192 -4304
rect 9242 -4364 9276 -4330
rect 9328 -4338 9362 -4304
rect 9406 -4338 9440 -4304
rect 9490 -4346 9524 -4312
rect 9490 -4414 9524 -4380
rect 9625 -4338 9659 -4304
rect 9625 -4406 9659 -4372
rect 9722 -4338 9756 -4304
rect 9722 -4406 9756 -4372
rect 9490 -4482 9524 -4448
rect 9722 -4474 9756 -4440
rect 9806 -4374 9840 -4340
rect 9806 -4442 9840 -4408
rect 9921 -4346 9955 -4312
rect 9921 -4414 9955 -4380
rect 10005 -4362 10039 -4328
rect 10089 -4346 10123 -4312
rect 10272 -4338 10306 -4304
rect 10356 -4346 10390 -4312
rect 10449 -4340 10483 -4306
rect 10603 -4364 10637 -4330
rect 10700 -4348 10734 -4314
rect 10784 -4364 10818 -4330
rect 10897 -4338 10931 -4304
rect 10089 -4414 10123 -4380
rect 10985 -4346 11019 -4312
rect 11082 -4339 11116 -4305
rect 11274 -4338 11308 -4304
rect 11358 -4364 11392 -4330
rect 11444 -4338 11478 -4304
rect 11522 -4338 11556 -4304
rect 11606 -4346 11640 -4312
rect 11606 -4414 11640 -4380
rect 11741 -4338 11775 -4304
rect 11741 -4406 11775 -4372
rect 11838 -4338 11872 -4304
rect 11838 -4406 11872 -4372
rect 11606 -4482 11640 -4448
rect 11838 -4474 11872 -4440
rect 11922 -4374 11956 -4340
rect 11922 -4442 11956 -4408
rect 12037 -4346 12071 -4312
rect 12037 -4414 12071 -4380
rect 12121 -4362 12155 -4328
rect 12205 -4346 12239 -4312
rect 12388 -4338 12422 -4304
rect 12472 -4346 12506 -4312
rect 12565 -4340 12599 -4306
rect 12719 -4364 12753 -4330
rect 12816 -4348 12850 -4314
rect 12900 -4364 12934 -4330
rect 13013 -4338 13047 -4304
rect 12205 -4414 12239 -4380
rect 13101 -4346 13135 -4312
rect 13198 -4339 13232 -4305
rect 13390 -4338 13424 -4304
rect 13474 -4364 13508 -4330
rect 13560 -4338 13594 -4304
rect 13638 -4338 13672 -4304
rect 13722 -4346 13756 -4312
rect 13722 -4414 13756 -4380
rect 13857 -4338 13891 -4304
rect 13857 -4406 13891 -4372
rect 13954 -4338 13988 -4304
rect 13954 -4406 13988 -4372
rect 13722 -4482 13756 -4448
rect 13954 -4474 13988 -4440
rect 14038 -4374 14072 -4340
rect 14038 -4442 14072 -4408
rect 14153 -4346 14187 -4312
rect 14153 -4414 14187 -4380
rect 14237 -4362 14271 -4328
rect 14321 -4346 14355 -4312
rect 14504 -4338 14538 -4304
rect 14588 -4346 14622 -4312
rect 14681 -4340 14715 -4306
rect 14835 -4364 14869 -4330
rect 14932 -4348 14966 -4314
rect 15016 -4364 15050 -4330
rect 15129 -4338 15163 -4304
rect 14321 -4414 14355 -4380
rect 15217 -4346 15251 -4312
rect 15314 -4339 15348 -4305
rect 15506 -4338 15540 -4304
rect 15590 -4364 15624 -4330
rect 15676 -4338 15710 -4304
rect 15754 -4338 15788 -4304
rect 15838 -4346 15872 -4312
rect 15838 -4414 15872 -4380
rect 15973 -4338 16007 -4304
rect 15973 -4406 16007 -4372
rect 16070 -4338 16104 -4304
rect 16070 -4406 16104 -4372
rect 15838 -4482 15872 -4448
rect 16070 -4474 16104 -4440
rect 16154 -4374 16188 -4340
rect 16154 -4442 16188 -4408
rect 16269 -4346 16303 -4312
rect 16269 -4414 16303 -4380
rect 16353 -4362 16387 -4328
rect 16437 -4346 16471 -4312
rect 16620 -4338 16654 -4304
rect 16704 -4346 16738 -4312
rect 16797 -4340 16831 -4306
rect 16951 -4364 16985 -4330
rect 17048 -4348 17082 -4314
rect 17132 -4364 17166 -4330
rect 17245 -4338 17279 -4304
rect 16437 -4414 16471 -4380
rect 17333 -4346 17367 -4312
rect 17430 -4339 17464 -4305
rect 17622 -4338 17656 -4304
rect 17706 -4364 17740 -4330
rect 17792 -4338 17826 -4304
rect 17870 -4338 17904 -4304
rect 17954 -4346 17988 -4312
rect 17954 -4414 17988 -4380
rect 18089 -4338 18123 -4304
rect 18089 -4406 18123 -4372
rect 18186 -4338 18220 -4304
rect 18186 -4406 18220 -4372
rect 17954 -4482 17988 -4448
rect 18186 -4474 18220 -4440
rect 18270 -4374 18304 -4340
rect 18270 -4442 18304 -4408
rect 18385 -4346 18419 -4312
rect 18385 -4414 18419 -4380
rect 18469 -4362 18503 -4328
rect 18553 -4346 18587 -4312
rect 18736 -4338 18770 -4304
rect 18820 -4346 18854 -4312
rect 18913 -4340 18947 -4306
rect 19067 -4364 19101 -4330
rect 19164 -4348 19198 -4314
rect 19248 -4364 19282 -4330
rect 19361 -4338 19395 -4304
rect 18553 -4414 18587 -4380
rect 19449 -4346 19483 -4312
rect 19546 -4339 19580 -4305
rect 19738 -4338 19772 -4304
rect 19822 -4364 19856 -4330
rect 19908 -4338 19942 -4304
rect 19986 -4338 20020 -4304
rect 20070 -4346 20104 -4312
rect 20070 -4414 20104 -4380
rect 20205 -4338 20239 -4304
rect 20205 -4406 20239 -4372
rect 20302 -4338 20336 -4304
rect 20302 -4406 20336 -4372
rect 20070 -4482 20104 -4448
rect 20302 -4474 20336 -4440
rect 20386 -4374 20420 -4340
rect 20386 -4442 20420 -4408
rect 20501 -4346 20535 -4312
rect 20501 -4414 20535 -4380
rect 20585 -4362 20619 -4328
rect 20669 -4346 20703 -4312
rect 20852 -4338 20886 -4304
rect 20936 -4346 20970 -4312
rect 21029 -4340 21063 -4306
rect 21183 -4364 21217 -4330
rect 21280 -4348 21314 -4314
rect 21364 -4364 21398 -4330
rect 21477 -4338 21511 -4304
rect 20669 -4414 20703 -4380
rect 21565 -4346 21599 -4312
rect 21662 -4339 21696 -4305
rect 21854 -4338 21888 -4304
rect 21938 -4364 21972 -4330
rect 22024 -4338 22058 -4304
rect 22102 -4338 22136 -4304
rect 22186 -4346 22220 -4312
rect 22186 -4414 22220 -4380
rect 22321 -4338 22355 -4304
rect 22321 -4406 22355 -4372
rect 22418 -4338 22452 -4304
rect 22418 -4406 22452 -4372
rect 22186 -4482 22220 -4448
rect 22418 -4474 22452 -4440
rect 22502 -4374 22536 -4340
rect 22502 -4442 22536 -4408
rect 22617 -4346 22651 -4312
rect 22617 -4414 22651 -4380
rect 22701 -4362 22735 -4328
rect 22785 -4346 22819 -4312
rect 22968 -4338 23002 -4304
rect 23052 -4346 23086 -4312
rect 23145 -4340 23179 -4306
rect 23299 -4364 23333 -4330
rect 23396 -4348 23430 -4314
rect 23480 -4364 23514 -4330
rect 23593 -4338 23627 -4304
rect 22785 -4414 22819 -4380
rect 23681 -4346 23715 -4312
rect 23778 -4339 23812 -4305
rect 23970 -4338 24004 -4304
rect 24054 -4364 24088 -4330
rect 24140 -4338 24174 -4304
rect 24218 -4338 24252 -4304
rect 24302 -4346 24336 -4312
rect 24302 -4414 24336 -4380
rect 24437 -4338 24471 -4304
rect 24437 -4406 24471 -4372
rect 24534 -4338 24568 -4304
rect 24534 -4406 24568 -4372
rect 24302 -4482 24336 -4448
rect 24534 -4474 24568 -4440
rect 24618 -4374 24652 -4340
rect 24618 -4442 24652 -4408
rect 24733 -4346 24767 -4312
rect 24733 -4414 24767 -4380
rect 24817 -4362 24851 -4328
rect 24901 -4346 24935 -4312
rect 25084 -4338 25118 -4304
rect 25168 -4346 25202 -4312
rect 25261 -4340 25295 -4306
rect 25415 -4364 25449 -4330
rect 25512 -4348 25546 -4314
rect 25596 -4364 25630 -4330
rect 25709 -4338 25743 -4304
rect 24901 -4414 24935 -4380
rect 25797 -4346 25831 -4312
rect 25894 -4339 25928 -4305
rect 26086 -4338 26120 -4304
rect 26170 -4364 26204 -4330
rect 26256 -4338 26290 -4304
rect 26334 -4338 26368 -4304
rect 26418 -4346 26452 -4312
rect 26418 -4414 26452 -4380
rect 26553 -4338 26587 -4304
rect 26553 -4406 26587 -4372
rect 26650 -4338 26684 -4304
rect 26650 -4406 26684 -4372
rect 26418 -4482 26452 -4448
rect 26650 -4474 26684 -4440
rect 26734 -4374 26768 -4340
rect 26734 -4442 26768 -4408
rect 26849 -4346 26883 -4312
rect 26849 -4414 26883 -4380
rect 26933 -4362 26967 -4328
rect 27017 -4346 27051 -4312
rect 27200 -4338 27234 -4304
rect 27284 -4346 27318 -4312
rect 27377 -4340 27411 -4306
rect 27531 -4364 27565 -4330
rect 27628 -4348 27662 -4314
rect 27712 -4364 27746 -4330
rect 27825 -4338 27859 -4304
rect 27017 -4414 27051 -4380
rect 27913 -4346 27947 -4312
rect 28010 -4339 28044 -4305
rect 28202 -4338 28236 -4304
rect 28286 -4364 28320 -4330
rect 28372 -4338 28406 -4304
rect 28450 -4338 28484 -4304
rect 28534 -4346 28568 -4312
rect 28534 -4414 28568 -4380
rect 28669 -4338 28703 -4304
rect 28669 -4406 28703 -4372
rect 28766 -4338 28800 -4304
rect 28766 -4406 28800 -4372
rect 28534 -4482 28568 -4448
rect 28766 -4474 28800 -4440
rect 28850 -4374 28884 -4340
rect 28850 -4442 28884 -4408
rect 28965 -4346 28999 -4312
rect 28965 -4414 28999 -4380
rect 29049 -4362 29083 -4328
rect 29133 -4346 29167 -4312
rect 29316 -4338 29350 -4304
rect 29400 -4346 29434 -4312
rect 29493 -4340 29527 -4306
rect 29647 -4364 29681 -4330
rect 29744 -4348 29778 -4314
rect 29828 -4364 29862 -4330
rect 29941 -4338 29975 -4304
rect 29133 -4414 29167 -4380
rect 30029 -4346 30063 -4312
rect 30126 -4339 30160 -4305
rect 30318 -4338 30352 -4304
rect 30402 -4364 30436 -4330
rect 30488 -4338 30522 -4304
rect 30566 -4338 30600 -4304
rect 30650 -4346 30684 -4312
rect 30650 -4414 30684 -4380
rect 30785 -4338 30819 -4304
rect 30785 -4406 30819 -4372
rect 30882 -4338 30916 -4304
rect 30882 -4406 30916 -4372
rect 30650 -4482 30684 -4448
rect 30882 -4474 30916 -4440
rect 30966 -4374 31000 -4340
rect 30966 -4442 31000 -4408
rect 31081 -4346 31115 -4312
rect 31081 -4414 31115 -4380
rect 31165 -4362 31199 -4328
rect 31249 -4346 31283 -4312
rect 31432 -4338 31466 -4304
rect 31516 -4346 31550 -4312
rect 31609 -4340 31643 -4306
rect 31763 -4364 31797 -4330
rect 31860 -4348 31894 -4314
rect 31944 -4364 31978 -4330
rect 32057 -4338 32091 -4304
rect 31249 -4414 31283 -4380
rect 32145 -4346 32179 -4312
rect 32242 -4339 32276 -4305
rect 32434 -4338 32468 -4304
rect 32518 -4364 32552 -4330
rect 32604 -4338 32638 -4304
rect 32682 -4338 32716 -4304
rect 32766 -4346 32800 -4312
rect 32766 -4414 32800 -4380
rect 32901 -4338 32935 -4304
rect 32901 -4406 32935 -4372
rect 32998 -4338 33032 -4304
rect 32998 -4406 33032 -4372
rect 32766 -4482 32800 -4448
rect 32998 -4474 33032 -4440
rect 33082 -4374 33116 -4340
rect 33082 -4442 33116 -4408
rect 9388 -7719 9422 -7683
rect 9387 -7793 9421 -7757
rect 9387 -7866 9421 -7830
rect 9645 -7723 9679 -7687
rect 9645 -7793 9679 -7757
rect 9644 -7866 9678 -7830
rect 10048 -7719 10082 -7683
rect 10047 -7793 10081 -7757
rect 10047 -7866 10081 -7830
rect 10305 -7723 10339 -7687
rect 10305 -7793 10339 -7757
rect 10304 -7866 10338 -7830
rect 10518 -7719 10552 -7683
rect 10517 -7793 10551 -7757
rect 10517 -7866 10551 -7830
rect 10775 -7723 10809 -7687
rect 10775 -7793 10809 -7757
rect 10774 -7866 10808 -7830
rect 11120 -7723 11154 -7687
rect 11120 -7794 11154 -7758
rect 11120 -7865 11154 -7829
rect 11378 -7723 11412 -7687
rect 11378 -7794 11412 -7758
rect 11378 -7865 11412 -7829
rect 11636 -7723 11670 -7687
rect 11636 -7794 11670 -7758
rect 11636 -7865 11670 -7829
rect 11894 -7723 11928 -7687
rect 11894 -7794 11928 -7758
rect 11894 -7865 11928 -7829
rect 12152 -7723 12186 -7687
rect 12152 -7794 12186 -7758
rect 12152 -7865 12186 -7829
rect 12410 -7723 12444 -7687
rect 12410 -7794 12444 -7758
rect 12410 -7865 12444 -7829
rect 12935 -7723 12969 -7687
rect 12935 -7794 12969 -7758
rect 12935 -7865 12969 -7829
rect 13193 -7723 13227 -7687
rect 13193 -7794 13227 -7758
rect 13193 -7865 13227 -7829
rect 13451 -7723 13485 -7687
rect 13451 -7794 13485 -7758
rect 13451 -7865 13485 -7829
rect 13709 -7723 13743 -7687
rect 13709 -7794 13743 -7758
rect 13709 -7865 13743 -7829
rect 13967 -7723 14001 -7687
rect 13967 -7794 14001 -7758
rect 13967 -7865 14001 -7829
rect 14225 -7723 14259 -7687
rect 14225 -7794 14259 -7758
rect 14225 -7865 14259 -7829
rect 14741 -7723 14775 -7687
rect 14741 -7794 14775 -7758
rect 14741 -7865 14775 -7829
rect 14999 -7723 15033 -7687
rect 14999 -7794 15033 -7758
rect 14999 -7865 15033 -7829
rect 15257 -7723 15291 -7687
rect 15257 -7794 15291 -7758
rect 15257 -7865 15291 -7829
rect 15515 -7723 15549 -7687
rect 15515 -7794 15549 -7758
rect 15515 -7865 15549 -7829
rect 15773 -7723 15807 -7687
rect 15773 -7794 15807 -7758
rect 15773 -7865 15807 -7829
rect 16031 -7723 16065 -7687
rect 16031 -7794 16065 -7758
rect 16031 -7865 16065 -7829
rect 9330 -8723 9368 -8687
rect 9516 -8721 9554 -8685
rect 9691 -8721 9725 -8687
rect 10549 -8721 10583 -8687
rect 10716 -8723 10754 -8687
rect 10902 -8721 10940 -8685
rect 11086 -8723 11124 -8687
rect 11272 -8721 11310 -8685
rect 11508 -8723 11546 -8687
rect 11694 -8721 11732 -8685
rect 11930 -8723 11968 -8687
rect 12116 -8721 12154 -8685
rect 12361 -8721 12395 -8687
rect 13219 -8721 13253 -8687
rect 13430 -8723 13468 -8687
rect 13616 -8721 13654 -8685
rect 13800 -8723 13838 -8687
rect 13986 -8721 14024 -8685
rect 14222 -8723 14260 -8687
rect 14408 -8721 14446 -8685
rect 14644 -8723 14682 -8687
rect 14830 -8721 14868 -8685
rect 15024 -8720 15058 -8686
rect 15882 -8720 15916 -8686
rect 16084 -8723 16122 -8687
rect 16270 -8721 16308 -8685
rect 9330 -14405 9368 -14369
rect 9516 -14403 9554 -14367
rect 9683 -14403 9717 -14369
rect 10541 -14403 10575 -14369
rect 10716 -14406 10754 -14370
rect 10902 -14404 10940 -14368
rect 11086 -14406 11124 -14370
rect 11272 -14404 11310 -14368
rect 11508 -14406 11546 -14370
rect 11694 -14404 11732 -14368
rect 11930 -14406 11968 -14370
rect 12116 -14404 12154 -14368
rect 12360 -14403 12394 -14369
rect 13218 -14403 13252 -14369
rect 13430 -14402 13468 -14366
rect 13616 -14400 13654 -14364
rect 13800 -14402 13838 -14366
rect 13986 -14400 14024 -14364
rect 14222 -14402 14260 -14366
rect 14408 -14400 14446 -14364
rect 14644 -14402 14682 -14366
rect 14830 -14400 14868 -14364
rect 15024 -14402 15058 -14368
rect 15882 -14402 15916 -14368
rect 16028 -14405 16066 -14369
rect 16214 -14403 16252 -14367
rect 9375 -20329 9413 -20293
rect 9561 -20327 9599 -20291
rect 9691 -20328 9725 -20294
rect 10549 -20328 10583 -20294
rect 10716 -20331 10754 -20295
rect 10902 -20329 10940 -20293
rect 11086 -20331 11124 -20295
rect 11272 -20329 11310 -20293
rect 11508 -20331 11546 -20295
rect 11694 -20329 11732 -20293
rect 11930 -20331 11968 -20295
rect 12116 -20329 12154 -20293
rect 12361 -20328 12395 -20294
rect 13219 -20328 13253 -20294
rect 13417 -20331 13455 -20295
rect 13603 -20329 13641 -20293
rect 13787 -20331 13825 -20295
rect 13973 -20329 14011 -20293
rect 14209 -20331 14247 -20295
rect 14395 -20329 14433 -20293
rect 14631 -20331 14669 -20295
rect 14817 -20329 14855 -20293
rect 15024 -20327 15058 -20293
rect 15882 -20327 15916 -20293
rect 16654 -19946 16688 -19634
rect 16742 -19946 16776 -19634
rect 17044 -19948 17078 -19636
rect 17132 -19948 17166 -19636
<< psubdiff >>
rect -20494 56772 -18660 56858
rect -21182 56736 -18660 56772
rect -21182 56190 38928 56736
rect -21182 55462 -18978 56190
rect -17592 55462 -14978 56190
rect -13592 55462 -10978 56190
rect -9592 55462 -6978 56190
rect -5592 55462 -2978 56190
rect -1592 55462 1022 56190
rect 2408 55462 5022 56190
rect 6408 55462 9022 56190
rect 10408 55462 13022 56190
rect 14408 55462 17022 56190
rect 18408 55462 21022 56190
rect 22408 55462 25022 56190
rect 26408 55462 29022 56190
rect 30408 55462 33022 56190
rect 34408 55462 37022 56190
rect 38408 55462 38928 56190
rect -21182 54840 38928 55462
rect -21182 54026 -18660 54840
rect -21182 53298 -20714 54026
rect -19328 53298 -18660 54026
rect -21182 50026 -18660 53298
rect -21182 49298 -20714 50026
rect -19328 49298 -18660 50026
rect 36666 52988 38866 54840
rect 36666 52260 37064 52988
rect 38450 52260 38866 52988
rect -21182 46026 -18660 49298
rect -21182 45298 -20714 46026
rect -19328 45298 -18660 46026
rect -21182 42026 -18660 45298
rect 36666 48988 38866 52260
rect 36666 48260 37064 48988
rect 38450 48260 38866 48988
rect 36666 44988 38866 48260
rect 36666 44260 37064 44988
rect 38450 44260 38866 44988
rect -21182 41298 -20714 42026
rect -19328 41298 -18660 42026
rect -21182 38026 -18660 41298
rect -21182 37298 -20714 38026
rect -19328 37298 -18660 38026
rect -21182 34026 -18660 37298
rect 36666 40988 38866 44260
rect 36666 40260 37064 40988
rect 38450 40260 38866 40988
rect 36666 36988 38866 40260
rect 36666 36260 37064 36988
rect 38450 36260 38866 36988
rect -21182 33298 -20714 34026
rect -19328 33298 -18660 34026
rect -21182 30026 -18660 33298
rect 36666 32988 38866 36260
rect 36666 32260 37064 32988
rect 38450 32260 38866 32988
rect -21182 29298 -20714 30026
rect -19328 29298 -18660 30026
rect -21182 26026 -18660 29298
rect -21182 25298 -20714 26026
rect -19328 25298 -18660 26026
rect -21182 22026 -18660 25298
rect 36666 28988 38866 32260
rect 36666 28260 37064 28988
rect 38450 28260 38866 28988
rect 36666 24988 38866 28260
rect 36666 24260 37064 24988
rect 38450 24260 38866 24988
rect -21182 21298 -20714 22026
rect -19328 21298 -18660 22026
rect -21182 18026 -18660 21298
rect -21182 17298 -20714 18026
rect -19328 17298 -18660 18026
rect -21182 15410 -18660 17298
rect 36666 20988 38866 24260
rect 36666 20260 37064 20988
rect 38450 20260 38866 20988
rect 36666 16988 38866 20260
rect 36666 16260 37064 16988
rect 38450 16260 38866 16988
rect 36666 15410 38866 16260
rect -21182 14908 38866 15410
rect -21182 14180 -18052 14908
rect -16666 14180 -14052 14908
rect -12666 14180 -10052 14908
rect -8666 14180 -6052 14908
rect -4666 14180 -2052 14908
rect -666 14180 1948 14908
rect 3334 14180 5948 14908
rect 7334 14180 9948 14908
rect 11334 14180 13948 14908
rect 15334 14180 17948 14908
rect 19334 14180 21948 14908
rect 23334 14180 25948 14908
rect 27334 14180 29948 14908
rect 31334 14180 33948 14908
rect 35334 14180 38866 14908
rect -21182 13758 38866 14180
rect -21182 13666 -18660 13758
rect 36666 13698 38866 13758
rect -20494 13576 -18660 13666
rect 17792 12068 19104 12262
rect 17792 11574 18000 12068
rect 18960 11574 19104 12068
rect 17792 11354 19104 11574
rect -61896 2878 -61292 2894
rect -61896 2826 -61864 2878
rect -61806 2826 -61464 2878
rect -61406 2826 -61292 2878
rect -61896 2812 -61292 2826
rect 3316 1698 4628 1892
rect 3316 1204 3524 1698
rect 4484 1204 4628 1698
rect 3316 984 4628 1204
rect 10738 1514 12050 1708
rect 10738 1020 10946 1514
rect 11906 1020 12050 1514
rect 10738 800 12050 1020
rect 26104 2352 26418 2396
rect 26104 2182 26176 2352
rect 26352 2182 26418 2352
rect 31960 2340 32274 2384
rect 26104 2132 26418 2182
rect 17370 1832 18682 2026
rect 17370 1338 17578 1832
rect 18538 1338 18682 1832
rect 26104 1884 26416 2132
rect 31960 2170 32120 2340
rect 32204 2170 32274 2340
rect 31960 2132 32274 2170
rect 31956 2130 32274 2132
rect 32364 2206 32976 2274
rect 31956 1884 32276 2130
rect 26104 1866 32276 1884
rect 26104 1840 32274 1866
rect 26104 1670 26168 1840
rect 26344 1670 26628 1840
rect 26804 1670 27228 1840
rect 27404 1670 27828 1840
rect 28004 1670 28428 1840
rect 28604 1670 29028 1840
rect 29204 1670 29628 1840
rect 29804 1670 30228 1840
rect 30404 1670 30828 1840
rect 31004 1670 31428 1840
rect 31604 1670 32028 1840
rect 32204 1670 32274 1840
rect 32364 1746 32424 2206
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 26104 1666 32274 1670
rect 26104 1620 28472 1666
rect 28936 1620 32274 1666
rect 17370 1118 18682 1338
rect 28942 1014 30164 1066
rect 28942 1012 29330 1014
rect 28942 1010 29106 1012
rect 29030 862 29106 1010
rect 29256 864 29330 1012
rect 29480 864 29546 1014
rect 29696 1012 29946 1014
rect 29696 864 29738 1012
rect 29256 862 29738 864
rect 29888 864 29946 1012
rect 30096 864 30164 1014
rect 29888 862 30164 864
rect 29030 860 30164 862
rect 28942 818 30164 860
rect 28984 816 29014 818
rect 29910 790 30160 818
rect 29910 640 29956 790
rect 30106 640 30160 790
rect 29910 598 30160 640
rect 29910 448 29962 598
rect 30112 448 30160 598
rect 29910 404 30160 448
rect 29910 294 29966 404
rect 29912 254 29966 294
rect 30116 254 30160 404
rect 29912 218 30160 254
rect 29912 68 29968 218
rect 30118 68 30160 218
rect 29912 32 30160 68
rect 29912 -88 29974 32
rect 29910 -118 29974 -88
rect 30124 -118 30160 32
rect 29910 -176 30160 -118
rect 29910 -326 29970 -176
rect 30120 -324 30160 -176
rect 30120 -326 30162 -324
rect 29910 -382 30162 -326
rect 29910 -412 30160 -382
rect 29910 -446 29964 -412
rect 29868 -450 29964 -446
rect 29808 -452 29964 -450
rect 28880 -488 29964 -452
rect 28880 -636 28912 -488
rect 29062 -490 29964 -488
rect 29062 -636 29124 -490
rect 28880 -640 29124 -636
rect 29274 -496 29964 -490
rect 29274 -640 29332 -496
rect 28880 -646 29332 -640
rect 29482 -498 29964 -496
rect 29482 -500 29752 -498
rect 29482 -646 29540 -500
rect 28880 -650 29540 -646
rect 29690 -648 29752 -500
rect 29902 -562 29964 -498
rect 30114 -456 30160 -412
rect 30114 -562 30162 -456
rect 29902 -648 30162 -562
rect 29690 -650 30162 -648
rect 28880 -670 30162 -650
rect 28880 -680 30160 -670
rect 28908 -684 30160 -680
rect 29806 -692 30160 -684
rect 8734 -1564 8763 -1530
rect 8797 -1564 8855 -1530
rect 8889 -1564 8947 -1530
rect 8981 -1564 9039 -1530
rect 9073 -1564 9131 -1530
rect 9165 -1564 9223 -1530
rect 9257 -1564 9315 -1530
rect 9349 -1564 9407 -1530
rect 9441 -1564 9499 -1530
rect 9533 -1564 9591 -1530
rect 9625 -1564 9683 -1530
rect 9717 -1564 9775 -1530
rect 9809 -1564 9867 -1530
rect 9901 -1564 9959 -1530
rect 9993 -1564 10051 -1530
rect 10085 -1564 10143 -1530
rect 10177 -1564 10235 -1530
rect 10269 -1564 10327 -1530
rect 10361 -1564 10419 -1530
rect 10453 -1564 10511 -1530
rect 10545 -1564 10603 -1530
rect 10637 -1564 10695 -1530
rect 10729 -1564 10787 -1530
rect 10821 -1564 10850 -1530
rect 11200 -1563 11229 -1529
rect 11263 -1563 11321 -1529
rect 11355 -1563 11413 -1529
rect 11447 -1563 11505 -1529
rect 11539 -1563 11597 -1529
rect 11631 -1563 11689 -1529
rect 11723 -1563 11781 -1529
rect 11815 -1563 11873 -1529
rect 11907 -1563 11965 -1529
rect 11999 -1563 12057 -1529
rect 12091 -1563 12149 -1529
rect 12183 -1563 12241 -1529
rect 12275 -1563 12333 -1529
rect 12367 -1563 12425 -1529
rect 12459 -1563 12517 -1529
rect 12551 -1563 12609 -1529
rect 12643 -1563 12701 -1529
rect 12735 -1563 12793 -1529
rect 12827 -1563 12885 -1529
rect 12919 -1563 12977 -1529
rect 13011 -1563 13069 -1529
rect 13103 -1563 13161 -1529
rect 13195 -1563 13253 -1529
rect 13287 -1563 13316 -1529
rect 10152 -2364 10181 -2330
rect 10215 -2364 10273 -2330
rect 10307 -2364 10365 -2330
rect 10399 -2364 10428 -2330
rect 11199 -2366 11229 -2332
rect 11263 -2366 11321 -2332
rect 11355 -2366 11413 -2332
rect 11447 -2366 11505 -2332
rect 11539 -2366 11597 -2332
rect 11631 -2366 11689 -2332
rect 11723 -2366 11781 -2332
rect 11815 -2366 11873 -2332
rect 11907 -2366 11965 -2332
rect 11999 -2366 12057 -2332
rect 12091 -2366 12149 -2332
rect 12183 -2366 12241 -2332
rect 12275 -2366 12333 -2332
rect 12367 -2366 12425 -2332
rect 12459 -2366 12517 -2332
rect 12551 -2366 12609 -2332
rect 12643 -2366 12701 -2332
rect 12735 -2366 12793 -2332
rect 12827 -2366 12885 -2332
rect 12919 -2366 12977 -2332
rect 13011 -2366 13069 -2332
rect 13103 -2366 13161 -2332
rect 13195 -2366 13253 -2332
rect 13287 -2366 13316 -2332
rect -9158 -4830 -9129 -4796
rect -9095 -4830 -9037 -4796
rect -9003 -4830 -8945 -4796
rect -8911 -4830 -8853 -4796
rect -8819 -4830 -8761 -4796
rect -8727 -4830 -8669 -4796
rect -8635 -4830 -8577 -4796
rect -8543 -4830 -8485 -4796
rect -8451 -4830 -8393 -4796
rect -8359 -4830 -8301 -4796
rect -8267 -4830 -8209 -4796
rect -8175 -4830 -8117 -4796
rect -8083 -4830 -8025 -4796
rect -7991 -4830 -7933 -4796
rect -7899 -4830 -7841 -4796
rect -7807 -4830 -7749 -4796
rect -7715 -4830 -7657 -4796
rect -7623 -4830 -7565 -4796
rect -7531 -4830 -7473 -4796
rect -7439 -4830 -7381 -4796
rect -7347 -4830 -7289 -4796
rect -7255 -4830 -7197 -4796
rect -7163 -4830 -7105 -4796
rect -7071 -4830 -7013 -4796
rect -6979 -4830 -6921 -4796
rect -6887 -4830 -6829 -4796
rect -6795 -4830 -6737 -4796
rect -6703 -4830 -6645 -4796
rect -6611 -4830 -6553 -4796
rect -6519 -4830 -6461 -4796
rect -6427 -4830 -6369 -4796
rect -6335 -4830 -6277 -4796
rect -6243 -4830 -6185 -4796
rect -6151 -4830 -6093 -4796
rect -6059 -4830 -6001 -4796
rect -5967 -4830 -5909 -4796
rect -5875 -4830 -5817 -4796
rect -5783 -4830 -5725 -4796
rect -5691 -4830 -5633 -4796
rect -5599 -4830 -5541 -4796
rect -5507 -4830 -5449 -4796
rect -5415 -4830 -5357 -4796
rect -5323 -4830 -5265 -4796
rect -5231 -4830 -5173 -4796
rect -5139 -4830 -5081 -4796
rect -5047 -4830 -4989 -4796
rect -4955 -4830 -4897 -4796
rect -4863 -4830 -4805 -4796
rect -4771 -4830 -4713 -4796
rect -4679 -4830 -4621 -4796
rect -4587 -4830 -4529 -4796
rect -4495 -4830 -4437 -4796
rect -4403 -4830 -4345 -4796
rect -4311 -4830 -4253 -4796
rect -4219 -4830 -4161 -4796
rect -4127 -4830 -4069 -4796
rect -4035 -4830 -3977 -4796
rect -3943 -4830 -3885 -4796
rect -3851 -4830 -3793 -4796
rect -3759 -4830 -3701 -4796
rect -3667 -4830 -3609 -4796
rect -3575 -4830 -3517 -4796
rect -3483 -4830 -3425 -4796
rect -3391 -4830 -3333 -4796
rect -3299 -4830 -3241 -4796
rect -3207 -4830 -3149 -4796
rect -3115 -4830 -3057 -4796
rect -3023 -4830 -2965 -4796
rect -2931 -4830 -2873 -4796
rect -2839 -4830 -2781 -4796
rect -2747 -4830 -2689 -4796
rect -2655 -4830 -2597 -4796
rect -2563 -4830 -2505 -4796
rect -2471 -4830 -2413 -4796
rect -2379 -4830 -2321 -4796
rect -2287 -4830 -2229 -4796
rect -2195 -4830 -2137 -4796
rect -2103 -4830 -2045 -4796
rect -2011 -4830 -1953 -4796
rect -1919 -4830 -1861 -4796
rect -1827 -4830 -1769 -4796
rect -1735 -4830 -1677 -4796
rect -1643 -4830 -1585 -4796
rect -1551 -4830 -1493 -4796
rect -1459 -4830 -1401 -4796
rect -1367 -4830 -1309 -4796
rect -1275 -4830 -1217 -4796
rect -1183 -4830 -1125 -4796
rect -1091 -4830 -1033 -4796
rect -999 -4830 -941 -4796
rect -907 -4830 -849 -4796
rect -815 -4830 -757 -4796
rect -723 -4830 -665 -4796
rect -631 -4830 -573 -4796
rect -539 -4830 -481 -4796
rect -447 -4830 -389 -4796
rect -355 -4830 -297 -4796
rect -263 -4830 -205 -4796
rect -171 -4830 -113 -4796
rect -79 -4830 -21 -4796
rect 13 -4830 71 -4796
rect 105 -4830 163 -4796
rect 197 -4830 255 -4796
rect 289 -4830 347 -4796
rect 381 -4830 439 -4796
rect 473 -4830 531 -4796
rect 565 -4830 623 -4796
rect 657 -4830 715 -4796
rect 749 -4830 807 -4796
rect 841 -4830 899 -4796
rect 933 -4830 991 -4796
rect 1025 -4830 1083 -4796
rect 1117 -4830 1175 -4796
rect 1209 -4830 1267 -4796
rect 1301 -4830 1359 -4796
rect 1393 -4830 1451 -4796
rect 1485 -4830 1543 -4796
rect 1577 -4830 1635 -4796
rect 1669 -4830 1727 -4796
rect 1761 -4830 1819 -4796
rect 1853 -4830 1911 -4796
rect 1945 -4830 2003 -4796
rect 2037 -4830 2095 -4796
rect 2129 -4830 2187 -4796
rect 2221 -4830 2279 -4796
rect 2313 -4830 2371 -4796
rect 2405 -4830 2463 -4796
rect 2497 -4830 2555 -4796
rect 2589 -4830 2647 -4796
rect 2681 -4830 2739 -4796
rect 2773 -4830 2831 -4796
rect 2865 -4830 2923 -4796
rect 2957 -4830 3015 -4796
rect 3049 -4830 3107 -4796
rect 3141 -4830 3199 -4796
rect 3233 -4830 3291 -4796
rect 3325 -4830 3383 -4796
rect 3417 -4830 3475 -4796
rect 3509 -4830 3567 -4796
rect 3601 -4830 3659 -4796
rect 3693 -4830 3751 -4796
rect 3785 -4830 3843 -4796
rect 3877 -4830 3935 -4796
rect 3969 -4830 4027 -4796
rect 4061 -4830 4119 -4796
rect 4153 -4830 4211 -4796
rect 4245 -4830 4303 -4796
rect 4337 -4830 4395 -4796
rect 4429 -4830 4487 -4796
rect 4521 -4830 4579 -4796
rect 4613 -4830 4671 -4796
rect 4705 -4830 4763 -4796
rect 4797 -4830 4855 -4796
rect 4889 -4830 4947 -4796
rect 4981 -4830 5039 -4796
rect 5073 -4830 5131 -4796
rect 5165 -4830 5223 -4796
rect 5257 -4830 5315 -4796
rect 5349 -4830 5407 -4796
rect 5441 -4830 5499 -4796
rect 5533 -4830 5591 -4796
rect 5625 -4830 5683 -4796
rect 5717 -4830 5775 -4796
rect 5809 -4830 5867 -4796
rect 5901 -4830 5959 -4796
rect 5993 -4830 6051 -4796
rect 6085 -4830 6143 -4796
rect 6177 -4830 6235 -4796
rect 6269 -4830 6327 -4796
rect 6361 -4830 6419 -4796
rect 6453 -4830 6511 -4796
rect 6545 -4830 6603 -4796
rect 6637 -4830 6695 -4796
rect 6729 -4830 6787 -4796
rect 6821 -4830 6879 -4796
rect 6913 -4830 6971 -4796
rect 7005 -4830 7063 -4796
rect 7097 -4830 7155 -4796
rect 7189 -4830 7247 -4796
rect 7281 -4830 7339 -4796
rect 7373 -4830 7431 -4796
rect 7465 -4830 7523 -4796
rect 7557 -4830 7615 -4796
rect 7649 -4830 7707 -4796
rect 7741 -4830 7799 -4796
rect 7833 -4830 7891 -4796
rect 7925 -4830 7983 -4796
rect 8017 -4830 8075 -4796
rect 8109 -4830 8167 -4796
rect 8201 -4830 8259 -4796
rect 8293 -4830 8351 -4796
rect 8385 -4830 8443 -4796
rect 8477 -4830 8535 -4796
rect 8569 -4830 8627 -4796
rect 8661 -4830 8719 -4796
rect 8753 -4830 8811 -4796
rect 8845 -4830 8903 -4796
rect 8937 -4830 8995 -4796
rect 9029 -4830 9087 -4796
rect 9121 -4830 9179 -4796
rect 9213 -4830 9271 -4796
rect 9305 -4830 9363 -4796
rect 9397 -4830 9455 -4796
rect 9489 -4830 9547 -4796
rect 9581 -4830 9639 -4796
rect 9673 -4830 9731 -4796
rect 9765 -4830 9823 -4796
rect 9857 -4830 9915 -4796
rect 9949 -4830 10007 -4796
rect 10041 -4830 10099 -4796
rect 10133 -4830 10191 -4796
rect 10225 -4830 10283 -4796
rect 10317 -4830 10375 -4796
rect 10409 -4830 10467 -4796
rect 10501 -4830 10559 -4796
rect 10593 -4830 10651 -4796
rect 10685 -4830 10743 -4796
rect 10777 -4830 10835 -4796
rect 10869 -4830 10927 -4796
rect 10961 -4830 11019 -4796
rect 11053 -4830 11111 -4796
rect 11145 -4830 11203 -4796
rect 11237 -4830 11295 -4796
rect 11329 -4830 11387 -4796
rect 11421 -4830 11479 -4796
rect 11513 -4830 11571 -4796
rect 11605 -4830 11663 -4796
rect 11697 -4830 11755 -4796
rect 11789 -4830 11847 -4796
rect 11881 -4830 11939 -4796
rect 11973 -4830 12031 -4796
rect 12065 -4830 12123 -4796
rect 12157 -4830 12215 -4796
rect 12249 -4830 12307 -4796
rect 12341 -4830 12399 -4796
rect 12433 -4830 12491 -4796
rect 12525 -4830 12583 -4796
rect 12617 -4830 12675 -4796
rect 12709 -4830 12767 -4796
rect 12801 -4830 12859 -4796
rect 12893 -4830 12951 -4796
rect 12985 -4830 13043 -4796
rect 13077 -4830 13135 -4796
rect 13169 -4830 13227 -4796
rect 13261 -4830 13319 -4796
rect 13353 -4830 13411 -4796
rect 13445 -4830 13503 -4796
rect 13537 -4830 13595 -4796
rect 13629 -4830 13687 -4796
rect 13721 -4830 13779 -4796
rect 13813 -4830 13871 -4796
rect 13905 -4830 13963 -4796
rect 13997 -4830 14055 -4796
rect 14089 -4830 14147 -4796
rect 14181 -4830 14239 -4796
rect 14273 -4830 14331 -4796
rect 14365 -4830 14423 -4796
rect 14457 -4830 14515 -4796
rect 14549 -4830 14607 -4796
rect 14641 -4830 14699 -4796
rect 14733 -4830 14791 -4796
rect 14825 -4830 14883 -4796
rect 14917 -4830 14975 -4796
rect 15009 -4830 15067 -4796
rect 15101 -4830 15159 -4796
rect 15193 -4830 15251 -4796
rect 15285 -4830 15343 -4796
rect 15377 -4830 15435 -4796
rect 15469 -4830 15527 -4796
rect 15561 -4830 15619 -4796
rect 15653 -4830 15711 -4796
rect 15745 -4830 15803 -4796
rect 15837 -4830 15895 -4796
rect 15929 -4830 15987 -4796
rect 16021 -4830 16079 -4796
rect 16113 -4830 16171 -4796
rect 16205 -4830 16263 -4796
rect 16297 -4830 16355 -4796
rect 16389 -4830 16447 -4796
rect 16481 -4830 16539 -4796
rect 16573 -4830 16631 -4796
rect 16665 -4830 16723 -4796
rect 16757 -4830 16815 -4796
rect 16849 -4830 16907 -4796
rect 16941 -4830 16999 -4796
rect 17033 -4830 17091 -4796
rect 17125 -4830 17183 -4796
rect 17217 -4830 17275 -4796
rect 17309 -4830 17367 -4796
rect 17401 -4830 17459 -4796
rect 17493 -4830 17551 -4796
rect 17585 -4830 17643 -4796
rect 17677 -4830 17735 -4796
rect 17769 -4830 17827 -4796
rect 17861 -4830 17919 -4796
rect 17953 -4830 18011 -4796
rect 18045 -4830 18103 -4796
rect 18137 -4830 18195 -4796
rect 18229 -4830 18287 -4796
rect 18321 -4830 18379 -4796
rect 18413 -4830 18471 -4796
rect 18505 -4830 18563 -4796
rect 18597 -4830 18655 -4796
rect 18689 -4830 18747 -4796
rect 18781 -4830 18839 -4796
rect 18873 -4830 18931 -4796
rect 18965 -4830 19023 -4796
rect 19057 -4830 19115 -4796
rect 19149 -4830 19207 -4796
rect 19241 -4830 19299 -4796
rect 19333 -4830 19391 -4796
rect 19425 -4830 19483 -4796
rect 19517 -4830 19575 -4796
rect 19609 -4830 19667 -4796
rect 19701 -4830 19759 -4796
rect 19793 -4830 19851 -4796
rect 19885 -4830 19943 -4796
rect 19977 -4830 20035 -4796
rect 20069 -4830 20127 -4796
rect 20161 -4830 20219 -4796
rect 20253 -4830 20311 -4796
rect 20345 -4830 20403 -4796
rect 20437 -4830 20495 -4796
rect 20529 -4830 20587 -4796
rect 20621 -4830 20679 -4796
rect 20713 -4830 20771 -4796
rect 20805 -4830 20863 -4796
rect 20897 -4830 20955 -4796
rect 20989 -4830 21047 -4796
rect 21081 -4830 21139 -4796
rect 21173 -4830 21231 -4796
rect 21265 -4830 21323 -4796
rect 21357 -4830 21415 -4796
rect 21449 -4830 21507 -4796
rect 21541 -4830 21599 -4796
rect 21633 -4830 21691 -4796
rect 21725 -4830 21783 -4796
rect 21817 -4830 21875 -4796
rect 21909 -4830 21967 -4796
rect 22001 -4830 22059 -4796
rect 22093 -4830 22151 -4796
rect 22185 -4830 22243 -4796
rect 22277 -4830 22335 -4796
rect 22369 -4830 22427 -4796
rect 22461 -4830 22519 -4796
rect 22553 -4830 22611 -4796
rect 22645 -4830 22703 -4796
rect 22737 -4830 22795 -4796
rect 22829 -4830 22887 -4796
rect 22921 -4830 22979 -4796
rect 23013 -4830 23071 -4796
rect 23105 -4830 23163 -4796
rect 23197 -4830 23255 -4796
rect 23289 -4830 23347 -4796
rect 23381 -4830 23439 -4796
rect 23473 -4830 23531 -4796
rect 23565 -4830 23623 -4796
rect 23657 -4830 23715 -4796
rect 23749 -4830 23807 -4796
rect 23841 -4830 23899 -4796
rect 23933 -4830 23991 -4796
rect 24025 -4830 24083 -4796
rect 24117 -4830 24175 -4796
rect 24209 -4830 24267 -4796
rect 24301 -4830 24359 -4796
rect 24393 -4830 24451 -4796
rect 24485 -4830 24543 -4796
rect 24577 -4830 24635 -4796
rect 24669 -4830 24727 -4796
rect 24761 -4830 24819 -4796
rect 24853 -4830 24911 -4796
rect 24945 -4830 25003 -4796
rect 25037 -4830 25095 -4796
rect 25129 -4830 25187 -4796
rect 25221 -4830 25279 -4796
rect 25313 -4830 25371 -4796
rect 25405 -4830 25463 -4796
rect 25497 -4830 25555 -4796
rect 25589 -4830 25647 -4796
rect 25681 -4830 25739 -4796
rect 25773 -4830 25831 -4796
rect 25865 -4830 25923 -4796
rect 25957 -4830 26015 -4796
rect 26049 -4830 26107 -4796
rect 26141 -4830 26199 -4796
rect 26233 -4830 26291 -4796
rect 26325 -4830 26383 -4796
rect 26417 -4830 26475 -4796
rect 26509 -4830 26567 -4796
rect 26601 -4830 26659 -4796
rect 26693 -4830 26751 -4796
rect 26785 -4830 26843 -4796
rect 26877 -4830 26935 -4796
rect 26969 -4830 27027 -4796
rect 27061 -4830 27119 -4796
rect 27153 -4830 27211 -4796
rect 27245 -4830 27303 -4796
rect 27337 -4830 27395 -4796
rect 27429 -4830 27487 -4796
rect 27521 -4830 27579 -4796
rect 27613 -4830 27671 -4796
rect 27705 -4830 27763 -4796
rect 27797 -4830 27855 -4796
rect 27889 -4830 27947 -4796
rect 27981 -4830 28039 -4796
rect 28073 -4830 28131 -4796
rect 28165 -4830 28223 -4796
rect 28257 -4830 28315 -4796
rect 28349 -4830 28407 -4796
rect 28441 -4830 28499 -4796
rect 28533 -4830 28591 -4796
rect 28625 -4830 28683 -4796
rect 28717 -4830 28775 -4796
rect 28809 -4830 28867 -4796
rect 28901 -4830 28959 -4796
rect 28993 -4830 29051 -4796
rect 29085 -4830 29143 -4796
rect 29177 -4830 29235 -4796
rect 29269 -4830 29327 -4796
rect 29361 -4830 29419 -4796
rect 29453 -4830 29511 -4796
rect 29545 -4830 29603 -4796
rect 29637 -4830 29695 -4796
rect 29729 -4830 29787 -4796
rect 29821 -4830 29879 -4796
rect 29913 -4830 29971 -4796
rect 30005 -4830 30063 -4796
rect 30097 -4830 30155 -4796
rect 30189 -4830 30247 -4796
rect 30281 -4830 30339 -4796
rect 30373 -4830 30431 -4796
rect 30465 -4830 30523 -4796
rect 30557 -4830 30615 -4796
rect 30649 -4830 30707 -4796
rect 30741 -4830 30799 -4796
rect 30833 -4830 30891 -4796
rect 30925 -4830 30983 -4796
rect 31017 -4830 31075 -4796
rect 31109 -4830 31167 -4796
rect 31201 -4830 31259 -4796
rect 31293 -4830 31351 -4796
rect 31385 -4830 31443 -4796
rect 31477 -4830 31535 -4796
rect 31569 -4830 31627 -4796
rect 31661 -4830 31719 -4796
rect 31753 -4830 31811 -4796
rect 31845 -4830 31903 -4796
rect 31937 -4830 31995 -4796
rect 32029 -4830 32087 -4796
rect 32121 -4830 32179 -4796
rect 32213 -4830 32271 -4796
rect 32305 -4830 32363 -4796
rect 32397 -4830 32455 -4796
rect 32489 -4830 32547 -4796
rect 32581 -4830 32639 -4796
rect 32673 -4830 32731 -4796
rect 32765 -4830 32823 -4796
rect 32857 -4830 32915 -4796
rect 32949 -4830 33007 -4796
rect 33041 -4830 33099 -4796
rect 33133 -4830 33162 -4796
rect 4255 -7545 4289 -7520
rect 7799 -7545 7833 -7520
rect 4255 -25773 4289 -25711
rect 17876 -7544 17910 -7519
rect 8716 -9507 16880 -9377
rect 8716 -13149 8926 -9507
rect 16728 -13149 16878 -9507
rect 8716 -13161 16878 -13149
rect 8716 -13267 9970 -13161
rect 10076 -13267 12634 -13161
rect 12740 -13267 15296 -13161
rect 15402 -13267 16878 -13161
rect 8716 -13303 16878 -13267
rect 8716 -13307 8926 -13303
rect 8670 -15035 16930 -15029
rect 8670 -15217 16936 -15035
rect 8670 -18865 8862 -15217
rect 16758 -18865 16936 -15217
rect 8670 -18885 16936 -18865
rect 8670 -18979 9972 -18885
rect 10064 -18979 12640 -18885
rect 12732 -18979 15306 -18885
rect 15398 -18979 16936 -18885
rect 8670 -19013 16936 -18979
rect 16520 -20269 17312 -20235
rect 16520 -20415 16578 -20269
rect 16520 -20487 16526 -20415
rect 16570 -20487 16578 -20415
rect 16520 -20633 16578 -20487
rect 16846 -20415 16968 -20269
rect 16846 -20487 16916 -20415
rect 16960 -20487 16968 -20415
rect 16846 -20633 16968 -20487
rect 17236 -20633 17312 -20269
rect 16520 -20667 17312 -20633
rect 8514 -20915 17052 -20913
rect 8514 -21113 17054 -20915
rect 8514 -24747 8818 -21113
rect 16786 -24747 17054 -21113
rect 8514 -24781 17056 -24747
rect 8514 -24875 9972 -24781
rect 10064 -24875 12642 -24781
rect 12734 -24875 15308 -24781
rect 15400 -24875 17056 -24781
rect 8514 -25041 17056 -24875
rect 7799 -25773 7833 -25711
rect 4255 -25807 4351 -25773
rect 7737 -25807 7833 -25773
rect 21420 -7544 21454 -7519
rect 17876 -25772 17910 -25710
rect 21420 -25772 21454 -25710
rect 17876 -25806 17972 -25772
rect 21358 -25806 21454 -25772
<< nsubdiff >>
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -27834 19740 -26806 21200
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -27834 17740 -26806 19274
rect -96266 15740 -95320 17274
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -27834 15740 -26806 17274
rect -96266 13740 -95320 15274
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -27834 13740 -26806 15274
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -27834 11740 -26806 13274
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -27834 9740 -26806 11274
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -27834 7740 -26806 9274
rect -96266 5740 -95320 7274
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -27834 5740 -26806 7274
rect -96266 4182 -95320 5274
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 6168 6094 6682 6190
rect 1280 5776 1374 6016
rect 1700 5776 1794 6016
rect 1280 5678 1794 5776
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -96396 3740 -62544 3910
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -27834 3846 -26806 5274
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 6168 5756 6682 5854
rect 11480 5882 11994 5978
rect 11480 5642 11574 5882
rect 11900 5642 11994 5882
rect 11480 5544 11994 5642
rect 16916 5824 17430 5920
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect -60278 3740 -26756 3846
rect -96396 2966 -62544 3274
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect 29198 3698 29398 3700
rect 29198 3696 30464 3698
rect 30724 3696 32708 3698
rect 27402 3694 32708 3696
rect 26112 3574 32708 3694
rect 26112 3550 32242 3574
rect 26112 3304 26988 3550
rect 27236 3304 27988 3550
rect 28236 3304 28988 3550
rect 29236 3304 29988 3550
rect 30236 3304 30988 3550
rect 31236 3326 32242 3550
rect 32484 3326 32708 3574
rect 31236 3304 32708 3326
rect -60278 3224 -26756 3274
rect 26112 3138 32708 3304
rect 26112 3136 31508 3138
rect 31928 3136 32708 3138
rect 26112 3132 26874 3136
rect 27398 3134 27886 3136
rect 28412 3134 30242 3136
rect 31932 3058 32708 3136
rect 31932 2904 32714 3058
rect 31932 2660 32212 2904
rect 32460 2660 32714 2904
rect 31932 2500 32714 2660
rect 27894 1150 28162 1152
rect 28822 1150 28872 1156
rect 27894 1130 28872 1150
rect 27894 1128 28422 1130
rect 27894 934 27926 1128
rect 27892 930 27926 934
rect 28126 930 28182 1128
rect 27892 928 28182 930
rect 28382 930 28422 1128
rect 28622 1128 28872 1130
rect 28622 930 28656 1128
rect 28382 928 28656 930
rect 28830 928 28872 1128
rect 27892 906 28872 928
rect 27892 904 28410 906
rect 28822 904 28872 906
rect 27892 886 28148 904
rect 27894 876 28148 886
rect 27896 856 28148 876
rect 27896 844 27926 856
rect 27902 656 27926 844
rect 28126 834 28148 856
rect 28126 656 28146 834
rect 27902 622 28146 656
rect 27902 422 27926 622
rect 28126 422 28146 622
rect 27902 382 28146 422
rect 27902 182 27926 382
rect 28126 182 28146 382
rect 27902 144 28146 182
rect 27902 -48 27924 144
rect 28124 -48 28146 144
rect 27902 -88 28146 -48
rect 27902 -288 27926 -88
rect 28126 -288 28146 -88
rect 27902 -324 28146 -288
rect 27902 -504 27924 -324
rect 27892 -524 27924 -504
rect 28124 -458 28146 -324
rect 28124 -524 28148 -458
rect 27892 -708 28148 -524
rect 28766 -708 28804 -706
rect 27892 -736 28810 -708
rect 27892 -748 28042 -736
rect 8734 -968 8763 -934
rect 8797 -968 8855 -934
rect 8889 -968 8947 -934
rect 8981 -968 9039 -934
rect 9073 -968 9131 -934
rect 9165 -968 9223 -934
rect 9257 -968 9315 -934
rect 9349 -968 9407 -934
rect 9441 -968 9499 -934
rect 9533 -968 9591 -934
rect 9625 -968 9683 -934
rect 9717 -968 9775 -934
rect 9809 -968 9867 -934
rect 9901 -968 9959 -934
rect 9993 -968 10051 -934
rect 10085 -968 10143 -934
rect 10177 -968 10235 -934
rect 10269 -968 10327 -934
rect 10361 -968 10419 -934
rect 10453 -968 10511 -934
rect 10545 -968 10603 -934
rect 10637 -968 10695 -934
rect 10729 -968 10787 -934
rect 10821 -968 10851 -934
rect 11200 -968 11229 -934
rect 11263 -968 11321 -934
rect 11355 -968 11413 -934
rect 11447 -968 11505 -934
rect 11539 -968 11597 -934
rect 11631 -968 11689 -934
rect 11723 -968 11781 -934
rect 11815 -968 11873 -934
rect 11907 -968 11965 -934
rect 11999 -968 12057 -934
rect 12091 -968 12149 -934
rect 12183 -968 12241 -934
rect 12275 -968 12333 -934
rect 12367 -968 12425 -934
rect 12459 -968 12517 -934
rect 12551 -968 12609 -934
rect 12643 -968 12701 -934
rect 12735 -968 12793 -934
rect 12827 -968 12885 -934
rect 12919 -968 12977 -934
rect 13011 -968 13069 -934
rect 13103 -968 13161 -934
rect 13195 -968 13253 -934
rect 13287 -968 13317 -934
rect 27902 -936 28042 -748
rect 28242 -738 28810 -736
rect 28242 -936 28348 -738
rect 27902 -938 28348 -936
rect 28548 -938 28628 -738
rect 28790 -938 28810 -738
rect 27902 -960 28810 -938
rect 28762 -962 28810 -960
rect 10152 -1770 10181 -1736
rect 10215 -1770 10273 -1736
rect 10307 -1770 10365 -1736
rect 10399 -1770 10428 -1736
rect 11200 -1769 11229 -1735
rect 11263 -1769 11321 -1735
rect 11355 -1769 11413 -1735
rect 11447 -1769 11505 -1735
rect 11539 -1769 11597 -1735
rect 11631 -1769 11689 -1735
rect 11723 -1769 11781 -1735
rect 11815 -1769 11873 -1735
rect 11907 -1769 11965 -1735
rect 11999 -1769 12057 -1735
rect 12091 -1769 12149 -1735
rect 12183 -1769 12241 -1735
rect 12275 -1769 12333 -1735
rect 12367 -1769 12425 -1735
rect 12459 -1769 12517 -1735
rect 12551 -1769 12609 -1735
rect 12643 -1769 12701 -1735
rect 12735 -1769 12793 -1735
rect 12827 -1769 12885 -1735
rect 12919 -1769 12977 -1735
rect 13011 -1769 13069 -1735
rect 13103 -1769 13161 -1735
rect 13195 -1769 13253 -1735
rect 13287 -1769 13316 -1735
rect -9158 -4238 -9129 -4204
rect -9095 -4238 -9037 -4204
rect -9003 -4238 -8945 -4204
rect -8911 -4238 -8853 -4204
rect -8819 -4238 -8761 -4204
rect -8727 -4238 -8669 -4204
rect -8635 -4238 -8577 -4204
rect -8543 -4238 -8485 -4204
rect -8451 -4238 -8393 -4204
rect -8359 -4238 -8301 -4204
rect -8267 -4238 -8209 -4204
rect -8175 -4238 -8117 -4204
rect -8083 -4238 -8025 -4204
rect -7991 -4238 -7933 -4204
rect -7899 -4238 -7841 -4204
rect -7807 -4238 -7749 -4204
rect -7715 -4238 -7657 -4204
rect -7623 -4238 -7565 -4204
rect -7531 -4238 -7473 -4204
rect -7439 -4238 -7381 -4204
rect -7347 -4238 -7289 -4204
rect -7255 -4238 -7197 -4204
rect -7163 -4238 -7105 -4204
rect -7071 -4238 -7013 -4204
rect -6979 -4238 -6921 -4204
rect -6887 -4238 -6829 -4204
rect -6795 -4238 -6737 -4204
rect -6703 -4238 -6645 -4204
rect -6611 -4238 -6553 -4204
rect -6519 -4238 -6461 -4204
rect -6427 -4238 -6369 -4204
rect -6335 -4238 -6277 -4204
rect -6243 -4238 -6185 -4204
rect -6151 -4238 -6093 -4204
rect -6059 -4238 -6001 -4204
rect -5967 -4238 -5909 -4204
rect -5875 -4238 -5817 -4204
rect -5783 -4238 -5725 -4204
rect -5691 -4238 -5633 -4204
rect -5599 -4238 -5541 -4204
rect -5507 -4238 -5449 -4204
rect -5415 -4238 -5357 -4204
rect -5323 -4238 -5265 -4204
rect -5231 -4238 -5173 -4204
rect -5139 -4238 -5081 -4204
rect -5047 -4238 -4989 -4204
rect -4955 -4238 -4897 -4204
rect -4863 -4238 -4805 -4204
rect -4771 -4238 -4713 -4204
rect -4679 -4238 -4621 -4204
rect -4587 -4238 -4529 -4204
rect -4495 -4238 -4437 -4204
rect -4403 -4238 -4345 -4204
rect -4311 -4238 -4253 -4204
rect -4219 -4238 -4161 -4204
rect -4127 -4238 -4069 -4204
rect -4035 -4238 -3977 -4204
rect -3943 -4238 -3885 -4204
rect -3851 -4238 -3793 -4204
rect -3759 -4238 -3701 -4204
rect -3667 -4238 -3609 -4204
rect -3575 -4238 -3517 -4204
rect -3483 -4238 -3425 -4204
rect -3391 -4238 -3333 -4204
rect -3299 -4238 -3241 -4204
rect -3207 -4238 -3149 -4204
rect -3115 -4238 -3057 -4204
rect -3023 -4238 -2965 -4204
rect -2931 -4238 -2873 -4204
rect -2839 -4238 -2781 -4204
rect -2747 -4238 -2689 -4204
rect -2655 -4238 -2597 -4204
rect -2563 -4238 -2505 -4204
rect -2471 -4238 -2413 -4204
rect -2379 -4238 -2321 -4204
rect -2287 -4238 -2229 -4204
rect -2195 -4238 -2137 -4204
rect -2103 -4238 -2045 -4204
rect -2011 -4238 -1953 -4204
rect -1919 -4238 -1861 -4204
rect -1827 -4238 -1769 -4204
rect -1735 -4238 -1677 -4204
rect -1643 -4238 -1585 -4204
rect -1551 -4238 -1493 -4204
rect -1459 -4238 -1401 -4204
rect -1367 -4238 -1309 -4204
rect -1275 -4238 -1217 -4204
rect -1183 -4238 -1125 -4204
rect -1091 -4238 -1033 -4204
rect -999 -4238 -941 -4204
rect -907 -4238 -849 -4204
rect -815 -4238 -757 -4204
rect -723 -4238 -665 -4204
rect -631 -4238 -573 -4204
rect -539 -4238 -481 -4204
rect -447 -4238 -389 -4204
rect -355 -4238 -297 -4204
rect -263 -4238 -205 -4204
rect -171 -4238 -113 -4204
rect -79 -4238 -21 -4204
rect 13 -4238 71 -4204
rect 105 -4238 163 -4204
rect 197 -4238 255 -4204
rect 289 -4238 347 -4204
rect 381 -4238 439 -4204
rect 473 -4238 531 -4204
rect 565 -4238 623 -4204
rect 657 -4238 715 -4204
rect 749 -4238 807 -4204
rect 841 -4238 899 -4204
rect 933 -4238 991 -4204
rect 1025 -4238 1083 -4204
rect 1117 -4238 1175 -4204
rect 1209 -4238 1267 -4204
rect 1301 -4238 1359 -4204
rect 1393 -4238 1451 -4204
rect 1485 -4238 1543 -4204
rect 1577 -4238 1635 -4204
rect 1669 -4238 1727 -4204
rect 1761 -4238 1819 -4204
rect 1853 -4238 1911 -4204
rect 1945 -4238 2003 -4204
rect 2037 -4238 2095 -4204
rect 2129 -4238 2187 -4204
rect 2221 -4238 2279 -4204
rect 2313 -4238 2371 -4204
rect 2405 -4238 2463 -4204
rect 2497 -4238 2555 -4204
rect 2589 -4238 2647 -4204
rect 2681 -4238 2739 -4204
rect 2773 -4238 2831 -4204
rect 2865 -4238 2923 -4204
rect 2957 -4238 3015 -4204
rect 3049 -4238 3107 -4204
rect 3141 -4238 3199 -4204
rect 3233 -4238 3291 -4204
rect 3325 -4238 3383 -4204
rect 3417 -4238 3475 -4204
rect 3509 -4238 3567 -4204
rect 3601 -4238 3659 -4204
rect 3693 -4238 3751 -4204
rect 3785 -4238 3843 -4204
rect 3877 -4238 3935 -4204
rect 3969 -4238 4027 -4204
rect 4061 -4238 4119 -4204
rect 4153 -4238 4211 -4204
rect 4245 -4238 4303 -4204
rect 4337 -4238 4395 -4204
rect 4429 -4238 4487 -4204
rect 4521 -4238 4579 -4204
rect 4613 -4238 4671 -4204
rect 4705 -4238 4763 -4204
rect 4797 -4238 4855 -4204
rect 4889 -4238 4947 -4204
rect 4981 -4238 5039 -4204
rect 5073 -4238 5131 -4204
rect 5165 -4238 5223 -4204
rect 5257 -4238 5315 -4204
rect 5349 -4238 5407 -4204
rect 5441 -4238 5499 -4204
rect 5533 -4238 5591 -4204
rect 5625 -4238 5683 -4204
rect 5717 -4238 5775 -4204
rect 5809 -4238 5867 -4204
rect 5901 -4238 5959 -4204
rect 5993 -4238 6051 -4204
rect 6085 -4238 6143 -4204
rect 6177 -4238 6235 -4204
rect 6269 -4238 6327 -4204
rect 6361 -4238 6419 -4204
rect 6453 -4238 6511 -4204
rect 6545 -4238 6603 -4204
rect 6637 -4238 6695 -4204
rect 6729 -4238 6787 -4204
rect 6821 -4238 6879 -4204
rect 6913 -4238 6971 -4204
rect 7005 -4238 7063 -4204
rect 7097 -4238 7155 -4204
rect 7189 -4238 7247 -4204
rect 7281 -4238 7339 -4204
rect 7373 -4238 7431 -4204
rect 7465 -4238 7523 -4204
rect 7557 -4238 7615 -4204
rect 7649 -4238 7707 -4204
rect 7741 -4238 7799 -4204
rect 7833 -4238 7891 -4204
rect 7925 -4238 7983 -4204
rect 8017 -4238 8075 -4204
rect 8109 -4238 8167 -4204
rect 8201 -4238 8259 -4204
rect 8293 -4238 8351 -4204
rect 8385 -4238 8443 -4204
rect 8477 -4238 8535 -4204
rect 8569 -4238 8627 -4204
rect 8661 -4238 8719 -4204
rect 8753 -4238 8811 -4204
rect 8845 -4238 8903 -4204
rect 8937 -4238 8995 -4204
rect 9029 -4238 9087 -4204
rect 9121 -4238 9179 -4204
rect 9213 -4238 9271 -4204
rect 9305 -4238 9363 -4204
rect 9397 -4238 9455 -4204
rect 9489 -4238 9547 -4204
rect 9581 -4238 9639 -4204
rect 9673 -4238 9731 -4204
rect 9765 -4238 9823 -4204
rect 9857 -4238 9915 -4204
rect 9949 -4238 10007 -4204
rect 10041 -4238 10099 -4204
rect 10133 -4238 10191 -4204
rect 10225 -4238 10283 -4204
rect 10317 -4238 10375 -4204
rect 10409 -4238 10467 -4204
rect 10501 -4238 10559 -4204
rect 10593 -4238 10651 -4204
rect 10685 -4238 10743 -4204
rect 10777 -4238 10835 -4204
rect 10869 -4238 10927 -4204
rect 10961 -4238 11019 -4204
rect 11053 -4238 11111 -4204
rect 11145 -4238 11203 -4204
rect 11237 -4238 11295 -4204
rect 11329 -4238 11387 -4204
rect 11421 -4238 11479 -4204
rect 11513 -4238 11571 -4204
rect 11605 -4238 11663 -4204
rect 11697 -4238 11755 -4204
rect 11789 -4238 11847 -4204
rect 11881 -4238 11939 -4204
rect 11973 -4238 12031 -4204
rect 12065 -4238 12123 -4204
rect 12157 -4238 12215 -4204
rect 12249 -4238 12307 -4204
rect 12341 -4238 12399 -4204
rect 12433 -4238 12491 -4204
rect 12525 -4238 12583 -4204
rect 12617 -4238 12675 -4204
rect 12709 -4238 12767 -4204
rect 12801 -4238 12859 -4204
rect 12893 -4238 12951 -4204
rect 12985 -4238 13043 -4204
rect 13077 -4238 13135 -4204
rect 13169 -4238 13227 -4204
rect 13261 -4238 13319 -4204
rect 13353 -4238 13411 -4204
rect 13445 -4238 13503 -4204
rect 13537 -4238 13595 -4204
rect 13629 -4238 13687 -4204
rect 13721 -4238 13779 -4204
rect 13813 -4238 13871 -4204
rect 13905 -4238 13963 -4204
rect 13997 -4238 14055 -4204
rect 14089 -4238 14147 -4204
rect 14181 -4238 14239 -4204
rect 14273 -4238 14331 -4204
rect 14365 -4238 14423 -4204
rect 14457 -4238 14515 -4204
rect 14549 -4238 14607 -4204
rect 14641 -4238 14699 -4204
rect 14733 -4238 14791 -4204
rect 14825 -4238 14883 -4204
rect 14917 -4238 14975 -4204
rect 15009 -4238 15067 -4204
rect 15101 -4238 15159 -4204
rect 15193 -4238 15251 -4204
rect 15285 -4238 15343 -4204
rect 15377 -4238 15435 -4204
rect 15469 -4238 15527 -4204
rect 15561 -4238 15619 -4204
rect 15653 -4238 15711 -4204
rect 15745 -4238 15803 -4204
rect 15837 -4238 15895 -4204
rect 15929 -4238 15987 -4204
rect 16021 -4238 16079 -4204
rect 16113 -4238 16171 -4204
rect 16205 -4238 16263 -4204
rect 16297 -4238 16355 -4204
rect 16389 -4238 16447 -4204
rect 16481 -4238 16539 -4204
rect 16573 -4238 16631 -4204
rect 16665 -4238 16723 -4204
rect 16757 -4238 16815 -4204
rect 16849 -4238 16907 -4204
rect 16941 -4238 16999 -4204
rect 17033 -4238 17091 -4204
rect 17125 -4238 17183 -4204
rect 17217 -4238 17275 -4204
rect 17309 -4238 17367 -4204
rect 17401 -4238 17459 -4204
rect 17493 -4238 17551 -4204
rect 17585 -4238 17643 -4204
rect 17677 -4238 17735 -4204
rect 17769 -4238 17827 -4204
rect 17861 -4238 17919 -4204
rect 17953 -4238 18011 -4204
rect 18045 -4238 18103 -4204
rect 18137 -4238 18195 -4204
rect 18229 -4238 18287 -4204
rect 18321 -4238 18379 -4204
rect 18413 -4238 18471 -4204
rect 18505 -4238 18563 -4204
rect 18597 -4238 18655 -4204
rect 18689 -4238 18747 -4204
rect 18781 -4238 18839 -4204
rect 18873 -4238 18931 -4204
rect 18965 -4238 19023 -4204
rect 19057 -4238 19115 -4204
rect 19149 -4238 19207 -4204
rect 19241 -4238 19299 -4204
rect 19333 -4238 19391 -4204
rect 19425 -4238 19483 -4204
rect 19517 -4238 19575 -4204
rect 19609 -4238 19667 -4204
rect 19701 -4238 19759 -4204
rect 19793 -4238 19851 -4204
rect 19885 -4238 19943 -4204
rect 19977 -4238 20035 -4204
rect 20069 -4238 20127 -4204
rect 20161 -4238 20219 -4204
rect 20253 -4238 20311 -4204
rect 20345 -4238 20403 -4204
rect 20437 -4238 20495 -4204
rect 20529 -4238 20587 -4204
rect 20621 -4238 20679 -4204
rect 20713 -4238 20771 -4204
rect 20805 -4238 20863 -4204
rect 20897 -4238 20955 -4204
rect 20989 -4238 21047 -4204
rect 21081 -4238 21139 -4204
rect 21173 -4238 21231 -4204
rect 21265 -4238 21323 -4204
rect 21357 -4238 21415 -4204
rect 21449 -4238 21507 -4204
rect 21541 -4238 21599 -4204
rect 21633 -4238 21691 -4204
rect 21725 -4238 21783 -4204
rect 21817 -4238 21875 -4204
rect 21909 -4238 21967 -4204
rect 22001 -4238 22059 -4204
rect 22093 -4238 22151 -4204
rect 22185 -4238 22243 -4204
rect 22277 -4238 22335 -4204
rect 22369 -4238 22427 -4204
rect 22461 -4238 22519 -4204
rect 22553 -4238 22611 -4204
rect 22645 -4238 22703 -4204
rect 22737 -4238 22795 -4204
rect 22829 -4238 22887 -4204
rect 22921 -4238 22979 -4204
rect 23013 -4238 23071 -4204
rect 23105 -4238 23163 -4204
rect 23197 -4238 23255 -4204
rect 23289 -4238 23347 -4204
rect 23381 -4238 23439 -4204
rect 23473 -4238 23531 -4204
rect 23565 -4238 23623 -4204
rect 23657 -4238 23715 -4204
rect 23749 -4238 23807 -4204
rect 23841 -4238 23899 -4204
rect 23933 -4238 23991 -4204
rect 24025 -4238 24083 -4204
rect 24117 -4238 24175 -4204
rect 24209 -4238 24267 -4204
rect 24301 -4238 24359 -4204
rect 24393 -4238 24451 -4204
rect 24485 -4238 24543 -4204
rect 24577 -4238 24635 -4204
rect 24669 -4238 24727 -4204
rect 24761 -4238 24819 -4204
rect 24853 -4238 24911 -4204
rect 24945 -4238 25003 -4204
rect 25037 -4238 25095 -4204
rect 25129 -4238 25187 -4204
rect 25221 -4238 25279 -4204
rect 25313 -4238 25371 -4204
rect 25405 -4238 25463 -4204
rect 25497 -4238 25555 -4204
rect 25589 -4238 25647 -4204
rect 25681 -4238 25739 -4204
rect 25773 -4238 25831 -4204
rect 25865 -4238 25923 -4204
rect 25957 -4238 26015 -4204
rect 26049 -4238 26107 -4204
rect 26141 -4238 26199 -4204
rect 26233 -4238 26291 -4204
rect 26325 -4238 26383 -4204
rect 26417 -4238 26475 -4204
rect 26509 -4238 26567 -4204
rect 26601 -4238 26659 -4204
rect 26693 -4238 26751 -4204
rect 26785 -4238 26843 -4204
rect 26877 -4238 26935 -4204
rect 26969 -4238 27027 -4204
rect 27061 -4238 27119 -4204
rect 27153 -4238 27211 -4204
rect 27245 -4238 27303 -4204
rect 27337 -4238 27395 -4204
rect 27429 -4238 27487 -4204
rect 27521 -4238 27579 -4204
rect 27613 -4238 27671 -4204
rect 27705 -4238 27763 -4204
rect 27797 -4238 27855 -4204
rect 27889 -4238 27947 -4204
rect 27981 -4238 28039 -4204
rect 28073 -4238 28131 -4204
rect 28165 -4238 28223 -4204
rect 28257 -4238 28315 -4204
rect 28349 -4238 28407 -4204
rect 28441 -4238 28499 -4204
rect 28533 -4238 28591 -4204
rect 28625 -4238 28683 -4204
rect 28717 -4238 28775 -4204
rect 28809 -4238 28867 -4204
rect 28901 -4238 28959 -4204
rect 28993 -4238 29051 -4204
rect 29085 -4238 29143 -4204
rect 29177 -4238 29235 -4204
rect 29269 -4238 29327 -4204
rect 29361 -4238 29419 -4204
rect 29453 -4238 29511 -4204
rect 29545 -4238 29603 -4204
rect 29637 -4238 29695 -4204
rect 29729 -4238 29787 -4204
rect 29821 -4238 29879 -4204
rect 29913 -4238 29971 -4204
rect 30005 -4238 30063 -4204
rect 30097 -4238 30155 -4204
rect 30189 -4238 30247 -4204
rect 30281 -4238 30339 -4204
rect 30373 -4238 30431 -4204
rect 30465 -4238 30523 -4204
rect 30557 -4238 30615 -4204
rect 30649 -4238 30707 -4204
rect 30741 -4238 30799 -4204
rect 30833 -4238 30891 -4204
rect 30925 -4238 30983 -4204
rect 31017 -4238 31075 -4204
rect 31109 -4238 31167 -4204
rect 31201 -4238 31259 -4204
rect 31293 -4238 31351 -4204
rect 31385 -4238 31443 -4204
rect 31477 -4238 31535 -4204
rect 31569 -4238 31627 -4204
rect 31661 -4238 31719 -4204
rect 31753 -4238 31811 -4204
rect 31845 -4238 31903 -4204
rect 31937 -4238 31995 -4204
rect 32029 -4238 32087 -4204
rect 32121 -4238 32179 -4204
rect 32213 -4238 32271 -4204
rect 32305 -4238 32363 -4204
rect 32397 -4238 32455 -4204
rect 32489 -4238 32547 -4204
rect 32581 -4238 32639 -4204
rect 32673 -4238 32731 -4204
rect 32765 -4238 32823 -4204
rect 32857 -4238 32915 -4204
rect 32949 -4238 33007 -4204
rect 33041 -4238 33099 -4204
rect 33133 -4238 33162 -4204
rect 9006 -7313 9238 -7309
rect 8996 -7379 16690 -7313
rect 8996 -7474 10166 -7379
rect 10794 -7383 16690 -7379
rect 10794 -7474 12946 -7383
rect 8996 -7478 12946 -7474
rect 13574 -7478 16690 -7383
rect 8996 -7493 16690 -7478
rect 9006 -8675 9238 -7493
rect 16062 -7495 16690 -7493
rect 16406 -8135 16690 -7495
rect 9006 -8937 9055 -8675
rect 9192 -8937 9238 -8675
rect 16404 -8694 16690 -8135
rect 9006 -9033 9238 -8937
rect 16404 -8956 16474 -8694
rect 16611 -8956 16690 -8694
rect 16404 -9033 16690 -8956
rect 9004 -9269 16690 -9033
rect 9004 -9273 16558 -9269
rect 16062 -9275 16558 -9273
rect 8996 -13829 16608 -13825
rect 8990 -13835 16608 -13829
rect 8990 -13977 16658 -13835
rect 8990 -14241 9206 -13977
rect 8990 -14503 9014 -14241
rect 9151 -14503 9206 -14241
rect 8990 -14709 9206 -14503
rect 16358 -14248 16658 -13977
rect 16358 -14510 16428 -14248
rect 16565 -14510 16658 -14248
rect 16358 -14709 16658 -14510
rect 8990 -14849 16658 -14709
rect 8996 -14855 16658 -14849
rect 16500 -19441 16890 -19439
rect 16500 -19473 17280 -19441
rect 8689 -19537 9166 -19527
rect 8689 -19543 9310 -19537
rect 8689 -19545 16374 -19543
rect 16500 -19545 16574 -19473
rect 16844 -19475 17280 -19473
rect 8689 -19579 16574 -19545
rect 8689 -19723 16248 -19579
rect 8689 -20124 9273 -19723
rect 8689 -20385 8973 -20124
rect 9109 -20385 9273 -20124
rect 16104 -19893 16248 -19723
rect 16450 -19581 16574 -19579
rect 16450 -19749 16588 -19581
rect 16450 -19811 16510 -19749
rect 16566 -19811 16588 -19749
rect 16450 -19893 16588 -19811
rect 16104 -19895 16588 -19893
rect 16104 -19933 16574 -19895
rect 8689 -20565 9273 -20385
rect 16104 -20565 16374 -19933
rect 16500 -20103 16574 -19933
rect 16844 -19751 16964 -19475
rect 16844 -19813 16900 -19751
rect 16956 -19813 16964 -19751
rect 16844 -20103 16964 -19813
rect 17234 -20103 17280 -19475
rect 16500 -20133 17280 -20103
rect 16500 -20141 16800 -20133
rect 16500 -20143 16572 -20141
rect 16968 -20143 17280 -20133
rect 8689 -20744 16374 -20565
rect 9056 -20745 16374 -20744
<< psubdiffcont >>
rect -18978 55462 -17592 56190
rect -14978 55462 -13592 56190
rect -10978 55462 -9592 56190
rect -6978 55462 -5592 56190
rect -2978 55462 -1592 56190
rect 1022 55462 2408 56190
rect 5022 55462 6408 56190
rect 9022 55462 10408 56190
rect 13022 55462 14408 56190
rect 17022 55462 18408 56190
rect 21022 55462 22408 56190
rect 25022 55462 26408 56190
rect 29022 55462 30408 56190
rect 33022 55462 34408 56190
rect 37022 55462 38408 56190
rect -20714 53298 -19328 54026
rect -20714 49298 -19328 50026
rect 37064 52260 38450 52988
rect -20714 45298 -19328 46026
rect 37064 48260 38450 48988
rect 37064 44260 38450 44988
rect -20714 41298 -19328 42026
rect -20714 37298 -19328 38026
rect 37064 40260 38450 40988
rect 37064 36260 38450 36988
rect -20714 33298 -19328 34026
rect 37064 32260 38450 32988
rect -20714 29298 -19328 30026
rect -20714 25298 -19328 26026
rect 37064 28260 38450 28988
rect 37064 24260 38450 24988
rect -20714 21298 -19328 22026
rect -20714 17298 -19328 18026
rect 37064 20260 38450 20988
rect 37064 16260 38450 16988
rect -18052 14180 -16666 14908
rect -14052 14180 -12666 14908
rect -10052 14180 -8666 14908
rect -6052 14180 -4666 14908
rect -2052 14180 -666 14908
rect 1948 14180 3334 14908
rect 5948 14180 7334 14908
rect 9948 14180 11334 14908
rect 13948 14180 15334 14908
rect 17948 14180 19334 14908
rect 21948 14180 23334 14908
rect 25948 14180 27334 14908
rect 29948 14180 31334 14908
rect 33948 14180 35334 14908
rect 18000 11574 18960 12068
rect -61864 2826 -61806 2878
rect -61464 2826 -61406 2878
rect 3524 1204 4484 1698
rect 10946 1020 11906 1514
rect 26176 2182 26352 2352
rect 17578 1338 18538 1832
rect 32120 2170 32204 2340
rect 26168 1670 26344 1840
rect 26628 1670 26804 1840
rect 27228 1670 27404 1840
rect 27828 1670 28004 1840
rect 28428 1670 28604 1840
rect 29028 1670 29204 1840
rect 29628 1670 29804 1840
rect 30228 1670 30404 1840
rect 30828 1670 31004 1840
rect 31428 1670 31604 1840
rect 32028 1670 32204 1840
rect 32424 1746 32904 2206
rect 28942 860 29030 1010
rect 29106 862 29256 1012
rect 29330 864 29480 1014
rect 29546 864 29696 1014
rect 29738 862 29888 1012
rect 29946 864 30096 1014
rect 29956 640 30106 790
rect 29962 448 30112 598
rect 29966 254 30116 404
rect 29968 68 30118 218
rect 29974 -118 30124 32
rect 29970 -326 30120 -176
rect 28912 -636 29062 -488
rect 29124 -640 29274 -490
rect 29332 -646 29482 -496
rect 29540 -650 29690 -500
rect 29752 -648 29902 -498
rect 29964 -562 30114 -412
rect 8763 -1564 8797 -1530
rect 8855 -1564 8889 -1530
rect 8947 -1564 8981 -1530
rect 9039 -1564 9073 -1530
rect 9131 -1564 9165 -1530
rect 9223 -1564 9257 -1530
rect 9315 -1564 9349 -1530
rect 9407 -1564 9441 -1530
rect 9499 -1564 9533 -1530
rect 9591 -1564 9625 -1530
rect 9683 -1564 9717 -1530
rect 9775 -1564 9809 -1530
rect 9867 -1564 9901 -1530
rect 9959 -1564 9993 -1530
rect 10051 -1564 10085 -1530
rect 10143 -1564 10177 -1530
rect 10235 -1564 10269 -1530
rect 10327 -1564 10361 -1530
rect 10419 -1564 10453 -1530
rect 10511 -1564 10545 -1530
rect 10603 -1564 10637 -1530
rect 10695 -1564 10729 -1530
rect 10787 -1564 10821 -1530
rect 11229 -1563 11263 -1529
rect 11321 -1563 11355 -1529
rect 11413 -1563 11447 -1529
rect 11505 -1563 11539 -1529
rect 11597 -1563 11631 -1529
rect 11689 -1563 11723 -1529
rect 11781 -1563 11815 -1529
rect 11873 -1563 11907 -1529
rect 11965 -1563 11999 -1529
rect 12057 -1563 12091 -1529
rect 12149 -1563 12183 -1529
rect 12241 -1563 12275 -1529
rect 12333 -1563 12367 -1529
rect 12425 -1563 12459 -1529
rect 12517 -1563 12551 -1529
rect 12609 -1563 12643 -1529
rect 12701 -1563 12735 -1529
rect 12793 -1563 12827 -1529
rect 12885 -1563 12919 -1529
rect 12977 -1563 13011 -1529
rect 13069 -1563 13103 -1529
rect 13161 -1563 13195 -1529
rect 13253 -1563 13287 -1529
rect 10181 -2364 10215 -2330
rect 10273 -2364 10307 -2330
rect 10365 -2364 10399 -2330
rect 11229 -2366 11263 -2332
rect 11321 -2366 11355 -2332
rect 11413 -2366 11447 -2332
rect 11505 -2366 11539 -2332
rect 11597 -2366 11631 -2332
rect 11689 -2366 11723 -2332
rect 11781 -2366 11815 -2332
rect 11873 -2366 11907 -2332
rect 11965 -2366 11999 -2332
rect 12057 -2366 12091 -2332
rect 12149 -2366 12183 -2332
rect 12241 -2366 12275 -2332
rect 12333 -2366 12367 -2332
rect 12425 -2366 12459 -2332
rect 12517 -2366 12551 -2332
rect 12609 -2366 12643 -2332
rect 12701 -2366 12735 -2332
rect 12793 -2366 12827 -2332
rect 12885 -2366 12919 -2332
rect 12977 -2366 13011 -2332
rect 13069 -2366 13103 -2332
rect 13161 -2366 13195 -2332
rect 13253 -2366 13287 -2332
rect -9129 -4830 -9095 -4796
rect -9037 -4830 -9003 -4796
rect -8945 -4830 -8911 -4796
rect -8853 -4830 -8819 -4796
rect -8761 -4830 -8727 -4796
rect -8669 -4830 -8635 -4796
rect -8577 -4830 -8543 -4796
rect -8485 -4830 -8451 -4796
rect -8393 -4830 -8359 -4796
rect -8301 -4830 -8267 -4796
rect -8209 -4830 -8175 -4796
rect -8117 -4830 -8083 -4796
rect -8025 -4830 -7991 -4796
rect -7933 -4830 -7899 -4796
rect -7841 -4830 -7807 -4796
rect -7749 -4830 -7715 -4796
rect -7657 -4830 -7623 -4796
rect -7565 -4830 -7531 -4796
rect -7473 -4830 -7439 -4796
rect -7381 -4830 -7347 -4796
rect -7289 -4830 -7255 -4796
rect -7197 -4830 -7163 -4796
rect -7105 -4830 -7071 -4796
rect -7013 -4830 -6979 -4796
rect -6921 -4830 -6887 -4796
rect -6829 -4830 -6795 -4796
rect -6737 -4830 -6703 -4796
rect -6645 -4830 -6611 -4796
rect -6553 -4830 -6519 -4796
rect -6461 -4830 -6427 -4796
rect -6369 -4830 -6335 -4796
rect -6277 -4830 -6243 -4796
rect -6185 -4830 -6151 -4796
rect -6093 -4830 -6059 -4796
rect -6001 -4830 -5967 -4796
rect -5909 -4830 -5875 -4796
rect -5817 -4830 -5783 -4796
rect -5725 -4830 -5691 -4796
rect -5633 -4830 -5599 -4796
rect -5541 -4830 -5507 -4796
rect -5449 -4830 -5415 -4796
rect -5357 -4830 -5323 -4796
rect -5265 -4830 -5231 -4796
rect -5173 -4830 -5139 -4796
rect -5081 -4830 -5047 -4796
rect -4989 -4830 -4955 -4796
rect -4897 -4830 -4863 -4796
rect -4805 -4830 -4771 -4796
rect -4713 -4830 -4679 -4796
rect -4621 -4830 -4587 -4796
rect -4529 -4830 -4495 -4796
rect -4437 -4830 -4403 -4796
rect -4345 -4830 -4311 -4796
rect -4253 -4830 -4219 -4796
rect -4161 -4830 -4127 -4796
rect -4069 -4830 -4035 -4796
rect -3977 -4830 -3943 -4796
rect -3885 -4830 -3851 -4796
rect -3793 -4830 -3759 -4796
rect -3701 -4830 -3667 -4796
rect -3609 -4830 -3575 -4796
rect -3517 -4830 -3483 -4796
rect -3425 -4830 -3391 -4796
rect -3333 -4830 -3299 -4796
rect -3241 -4830 -3207 -4796
rect -3149 -4830 -3115 -4796
rect -3057 -4830 -3023 -4796
rect -2965 -4830 -2931 -4796
rect -2873 -4830 -2839 -4796
rect -2781 -4830 -2747 -4796
rect -2689 -4830 -2655 -4796
rect -2597 -4830 -2563 -4796
rect -2505 -4830 -2471 -4796
rect -2413 -4830 -2379 -4796
rect -2321 -4830 -2287 -4796
rect -2229 -4830 -2195 -4796
rect -2137 -4830 -2103 -4796
rect -2045 -4830 -2011 -4796
rect -1953 -4830 -1919 -4796
rect -1861 -4830 -1827 -4796
rect -1769 -4830 -1735 -4796
rect -1677 -4830 -1643 -4796
rect -1585 -4830 -1551 -4796
rect -1493 -4830 -1459 -4796
rect -1401 -4830 -1367 -4796
rect -1309 -4830 -1275 -4796
rect -1217 -4830 -1183 -4796
rect -1125 -4830 -1091 -4796
rect -1033 -4830 -999 -4796
rect -941 -4830 -907 -4796
rect -849 -4830 -815 -4796
rect -757 -4830 -723 -4796
rect -665 -4830 -631 -4796
rect -573 -4830 -539 -4796
rect -481 -4830 -447 -4796
rect -389 -4830 -355 -4796
rect -297 -4830 -263 -4796
rect -205 -4830 -171 -4796
rect -113 -4830 -79 -4796
rect -21 -4830 13 -4796
rect 71 -4830 105 -4796
rect 163 -4830 197 -4796
rect 255 -4830 289 -4796
rect 347 -4830 381 -4796
rect 439 -4830 473 -4796
rect 531 -4830 565 -4796
rect 623 -4830 657 -4796
rect 715 -4830 749 -4796
rect 807 -4830 841 -4796
rect 899 -4830 933 -4796
rect 991 -4830 1025 -4796
rect 1083 -4830 1117 -4796
rect 1175 -4830 1209 -4796
rect 1267 -4830 1301 -4796
rect 1359 -4830 1393 -4796
rect 1451 -4830 1485 -4796
rect 1543 -4830 1577 -4796
rect 1635 -4830 1669 -4796
rect 1727 -4830 1761 -4796
rect 1819 -4830 1853 -4796
rect 1911 -4830 1945 -4796
rect 2003 -4830 2037 -4796
rect 2095 -4830 2129 -4796
rect 2187 -4830 2221 -4796
rect 2279 -4830 2313 -4796
rect 2371 -4830 2405 -4796
rect 2463 -4830 2497 -4796
rect 2555 -4830 2589 -4796
rect 2647 -4830 2681 -4796
rect 2739 -4830 2773 -4796
rect 2831 -4830 2865 -4796
rect 2923 -4830 2957 -4796
rect 3015 -4830 3049 -4796
rect 3107 -4830 3141 -4796
rect 3199 -4830 3233 -4796
rect 3291 -4830 3325 -4796
rect 3383 -4830 3417 -4796
rect 3475 -4830 3509 -4796
rect 3567 -4830 3601 -4796
rect 3659 -4830 3693 -4796
rect 3751 -4830 3785 -4796
rect 3843 -4830 3877 -4796
rect 3935 -4830 3969 -4796
rect 4027 -4830 4061 -4796
rect 4119 -4830 4153 -4796
rect 4211 -4830 4245 -4796
rect 4303 -4830 4337 -4796
rect 4395 -4830 4429 -4796
rect 4487 -4830 4521 -4796
rect 4579 -4830 4613 -4796
rect 4671 -4830 4705 -4796
rect 4763 -4830 4797 -4796
rect 4855 -4830 4889 -4796
rect 4947 -4830 4981 -4796
rect 5039 -4830 5073 -4796
rect 5131 -4830 5165 -4796
rect 5223 -4830 5257 -4796
rect 5315 -4830 5349 -4796
rect 5407 -4830 5441 -4796
rect 5499 -4830 5533 -4796
rect 5591 -4830 5625 -4796
rect 5683 -4830 5717 -4796
rect 5775 -4830 5809 -4796
rect 5867 -4830 5901 -4796
rect 5959 -4830 5993 -4796
rect 6051 -4830 6085 -4796
rect 6143 -4830 6177 -4796
rect 6235 -4830 6269 -4796
rect 6327 -4830 6361 -4796
rect 6419 -4830 6453 -4796
rect 6511 -4830 6545 -4796
rect 6603 -4830 6637 -4796
rect 6695 -4830 6729 -4796
rect 6787 -4830 6821 -4796
rect 6879 -4830 6913 -4796
rect 6971 -4830 7005 -4796
rect 7063 -4830 7097 -4796
rect 7155 -4830 7189 -4796
rect 7247 -4830 7281 -4796
rect 7339 -4830 7373 -4796
rect 7431 -4830 7465 -4796
rect 7523 -4830 7557 -4796
rect 7615 -4830 7649 -4796
rect 7707 -4830 7741 -4796
rect 7799 -4830 7833 -4796
rect 7891 -4830 7925 -4796
rect 7983 -4830 8017 -4796
rect 8075 -4830 8109 -4796
rect 8167 -4830 8201 -4796
rect 8259 -4830 8293 -4796
rect 8351 -4830 8385 -4796
rect 8443 -4830 8477 -4796
rect 8535 -4830 8569 -4796
rect 8627 -4830 8661 -4796
rect 8719 -4830 8753 -4796
rect 8811 -4830 8845 -4796
rect 8903 -4830 8937 -4796
rect 8995 -4830 9029 -4796
rect 9087 -4830 9121 -4796
rect 9179 -4830 9213 -4796
rect 9271 -4830 9305 -4796
rect 9363 -4830 9397 -4796
rect 9455 -4830 9489 -4796
rect 9547 -4830 9581 -4796
rect 9639 -4830 9673 -4796
rect 9731 -4830 9765 -4796
rect 9823 -4830 9857 -4796
rect 9915 -4830 9949 -4796
rect 10007 -4830 10041 -4796
rect 10099 -4830 10133 -4796
rect 10191 -4830 10225 -4796
rect 10283 -4830 10317 -4796
rect 10375 -4830 10409 -4796
rect 10467 -4830 10501 -4796
rect 10559 -4830 10593 -4796
rect 10651 -4830 10685 -4796
rect 10743 -4830 10777 -4796
rect 10835 -4830 10869 -4796
rect 10927 -4830 10961 -4796
rect 11019 -4830 11053 -4796
rect 11111 -4830 11145 -4796
rect 11203 -4830 11237 -4796
rect 11295 -4830 11329 -4796
rect 11387 -4830 11421 -4796
rect 11479 -4830 11513 -4796
rect 11571 -4830 11605 -4796
rect 11663 -4830 11697 -4796
rect 11755 -4830 11789 -4796
rect 11847 -4830 11881 -4796
rect 11939 -4830 11973 -4796
rect 12031 -4830 12065 -4796
rect 12123 -4830 12157 -4796
rect 12215 -4830 12249 -4796
rect 12307 -4830 12341 -4796
rect 12399 -4830 12433 -4796
rect 12491 -4830 12525 -4796
rect 12583 -4830 12617 -4796
rect 12675 -4830 12709 -4796
rect 12767 -4830 12801 -4796
rect 12859 -4830 12893 -4796
rect 12951 -4830 12985 -4796
rect 13043 -4830 13077 -4796
rect 13135 -4830 13169 -4796
rect 13227 -4830 13261 -4796
rect 13319 -4830 13353 -4796
rect 13411 -4830 13445 -4796
rect 13503 -4830 13537 -4796
rect 13595 -4830 13629 -4796
rect 13687 -4830 13721 -4796
rect 13779 -4830 13813 -4796
rect 13871 -4830 13905 -4796
rect 13963 -4830 13997 -4796
rect 14055 -4830 14089 -4796
rect 14147 -4830 14181 -4796
rect 14239 -4830 14273 -4796
rect 14331 -4830 14365 -4796
rect 14423 -4830 14457 -4796
rect 14515 -4830 14549 -4796
rect 14607 -4830 14641 -4796
rect 14699 -4830 14733 -4796
rect 14791 -4830 14825 -4796
rect 14883 -4830 14917 -4796
rect 14975 -4830 15009 -4796
rect 15067 -4830 15101 -4796
rect 15159 -4830 15193 -4796
rect 15251 -4830 15285 -4796
rect 15343 -4830 15377 -4796
rect 15435 -4830 15469 -4796
rect 15527 -4830 15561 -4796
rect 15619 -4830 15653 -4796
rect 15711 -4830 15745 -4796
rect 15803 -4830 15837 -4796
rect 15895 -4830 15929 -4796
rect 15987 -4830 16021 -4796
rect 16079 -4830 16113 -4796
rect 16171 -4830 16205 -4796
rect 16263 -4830 16297 -4796
rect 16355 -4830 16389 -4796
rect 16447 -4830 16481 -4796
rect 16539 -4830 16573 -4796
rect 16631 -4830 16665 -4796
rect 16723 -4830 16757 -4796
rect 16815 -4830 16849 -4796
rect 16907 -4830 16941 -4796
rect 16999 -4830 17033 -4796
rect 17091 -4830 17125 -4796
rect 17183 -4830 17217 -4796
rect 17275 -4830 17309 -4796
rect 17367 -4830 17401 -4796
rect 17459 -4830 17493 -4796
rect 17551 -4830 17585 -4796
rect 17643 -4830 17677 -4796
rect 17735 -4830 17769 -4796
rect 17827 -4830 17861 -4796
rect 17919 -4830 17953 -4796
rect 18011 -4830 18045 -4796
rect 18103 -4830 18137 -4796
rect 18195 -4830 18229 -4796
rect 18287 -4830 18321 -4796
rect 18379 -4830 18413 -4796
rect 18471 -4830 18505 -4796
rect 18563 -4830 18597 -4796
rect 18655 -4830 18689 -4796
rect 18747 -4830 18781 -4796
rect 18839 -4830 18873 -4796
rect 18931 -4830 18965 -4796
rect 19023 -4830 19057 -4796
rect 19115 -4830 19149 -4796
rect 19207 -4830 19241 -4796
rect 19299 -4830 19333 -4796
rect 19391 -4830 19425 -4796
rect 19483 -4830 19517 -4796
rect 19575 -4830 19609 -4796
rect 19667 -4830 19701 -4796
rect 19759 -4830 19793 -4796
rect 19851 -4830 19885 -4796
rect 19943 -4830 19977 -4796
rect 20035 -4830 20069 -4796
rect 20127 -4830 20161 -4796
rect 20219 -4830 20253 -4796
rect 20311 -4830 20345 -4796
rect 20403 -4830 20437 -4796
rect 20495 -4830 20529 -4796
rect 20587 -4830 20621 -4796
rect 20679 -4830 20713 -4796
rect 20771 -4830 20805 -4796
rect 20863 -4830 20897 -4796
rect 20955 -4830 20989 -4796
rect 21047 -4830 21081 -4796
rect 21139 -4830 21173 -4796
rect 21231 -4830 21265 -4796
rect 21323 -4830 21357 -4796
rect 21415 -4830 21449 -4796
rect 21507 -4830 21541 -4796
rect 21599 -4830 21633 -4796
rect 21691 -4830 21725 -4796
rect 21783 -4830 21817 -4796
rect 21875 -4830 21909 -4796
rect 21967 -4830 22001 -4796
rect 22059 -4830 22093 -4796
rect 22151 -4830 22185 -4796
rect 22243 -4830 22277 -4796
rect 22335 -4830 22369 -4796
rect 22427 -4830 22461 -4796
rect 22519 -4830 22553 -4796
rect 22611 -4830 22645 -4796
rect 22703 -4830 22737 -4796
rect 22795 -4830 22829 -4796
rect 22887 -4830 22921 -4796
rect 22979 -4830 23013 -4796
rect 23071 -4830 23105 -4796
rect 23163 -4830 23197 -4796
rect 23255 -4830 23289 -4796
rect 23347 -4830 23381 -4796
rect 23439 -4830 23473 -4796
rect 23531 -4830 23565 -4796
rect 23623 -4830 23657 -4796
rect 23715 -4830 23749 -4796
rect 23807 -4830 23841 -4796
rect 23899 -4830 23933 -4796
rect 23991 -4830 24025 -4796
rect 24083 -4830 24117 -4796
rect 24175 -4830 24209 -4796
rect 24267 -4830 24301 -4796
rect 24359 -4830 24393 -4796
rect 24451 -4830 24485 -4796
rect 24543 -4830 24577 -4796
rect 24635 -4830 24669 -4796
rect 24727 -4830 24761 -4796
rect 24819 -4830 24853 -4796
rect 24911 -4830 24945 -4796
rect 25003 -4830 25037 -4796
rect 25095 -4830 25129 -4796
rect 25187 -4830 25221 -4796
rect 25279 -4830 25313 -4796
rect 25371 -4830 25405 -4796
rect 25463 -4830 25497 -4796
rect 25555 -4830 25589 -4796
rect 25647 -4830 25681 -4796
rect 25739 -4830 25773 -4796
rect 25831 -4830 25865 -4796
rect 25923 -4830 25957 -4796
rect 26015 -4830 26049 -4796
rect 26107 -4830 26141 -4796
rect 26199 -4830 26233 -4796
rect 26291 -4830 26325 -4796
rect 26383 -4830 26417 -4796
rect 26475 -4830 26509 -4796
rect 26567 -4830 26601 -4796
rect 26659 -4830 26693 -4796
rect 26751 -4830 26785 -4796
rect 26843 -4830 26877 -4796
rect 26935 -4830 26969 -4796
rect 27027 -4830 27061 -4796
rect 27119 -4830 27153 -4796
rect 27211 -4830 27245 -4796
rect 27303 -4830 27337 -4796
rect 27395 -4830 27429 -4796
rect 27487 -4830 27521 -4796
rect 27579 -4830 27613 -4796
rect 27671 -4830 27705 -4796
rect 27763 -4830 27797 -4796
rect 27855 -4830 27889 -4796
rect 27947 -4830 27981 -4796
rect 28039 -4830 28073 -4796
rect 28131 -4830 28165 -4796
rect 28223 -4830 28257 -4796
rect 28315 -4830 28349 -4796
rect 28407 -4830 28441 -4796
rect 28499 -4830 28533 -4796
rect 28591 -4830 28625 -4796
rect 28683 -4830 28717 -4796
rect 28775 -4830 28809 -4796
rect 28867 -4830 28901 -4796
rect 28959 -4830 28993 -4796
rect 29051 -4830 29085 -4796
rect 29143 -4830 29177 -4796
rect 29235 -4830 29269 -4796
rect 29327 -4830 29361 -4796
rect 29419 -4830 29453 -4796
rect 29511 -4830 29545 -4796
rect 29603 -4830 29637 -4796
rect 29695 -4830 29729 -4796
rect 29787 -4830 29821 -4796
rect 29879 -4830 29913 -4796
rect 29971 -4830 30005 -4796
rect 30063 -4830 30097 -4796
rect 30155 -4830 30189 -4796
rect 30247 -4830 30281 -4796
rect 30339 -4830 30373 -4796
rect 30431 -4830 30465 -4796
rect 30523 -4830 30557 -4796
rect 30615 -4830 30649 -4796
rect 30707 -4830 30741 -4796
rect 30799 -4830 30833 -4796
rect 30891 -4830 30925 -4796
rect 30983 -4830 31017 -4796
rect 31075 -4830 31109 -4796
rect 31167 -4830 31201 -4796
rect 31259 -4830 31293 -4796
rect 31351 -4830 31385 -4796
rect 31443 -4830 31477 -4796
rect 31535 -4830 31569 -4796
rect 31627 -4830 31661 -4796
rect 31719 -4830 31753 -4796
rect 31811 -4830 31845 -4796
rect 31903 -4830 31937 -4796
rect 31995 -4830 32029 -4796
rect 32087 -4830 32121 -4796
rect 32179 -4830 32213 -4796
rect 32271 -4830 32305 -4796
rect 32363 -4830 32397 -4796
rect 32455 -4830 32489 -4796
rect 32547 -4830 32581 -4796
rect 32639 -4830 32673 -4796
rect 32731 -4830 32765 -4796
rect 32823 -4830 32857 -4796
rect 32915 -4830 32949 -4796
rect 33007 -4830 33041 -4796
rect 33099 -4830 33133 -4796
rect 4255 -25711 4289 -7545
rect 7799 -25711 7833 -7545
rect 9970 -13267 10076 -13161
rect 12634 -13267 12740 -13161
rect 15296 -13267 15402 -13161
rect 9972 -18979 10064 -18885
rect 12640 -18979 12732 -18885
rect 15306 -18979 15398 -18885
rect 16526 -20487 16570 -20415
rect 16916 -20487 16960 -20415
rect 9972 -24875 10064 -24781
rect 12642 -24875 12734 -24781
rect 15308 -24875 15400 -24781
rect 4351 -25807 7737 -25773
rect 17876 -25710 17910 -7544
rect 21420 -25710 21454 -7544
rect 17972 -25806 21358 -25772
<< nsubdiffcont >>
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -27644 19274 -27112 19740
rect -96044 17274 -95512 17740
rect -27644 17274 -27112 17740
rect -96044 15274 -95512 15740
rect -27644 15274 -27112 15740
rect -96044 13274 -95512 13740
rect -27644 13274 -27112 13740
rect -96044 11274 -95512 11740
rect -27644 11274 -27112 11740
rect -96044 9274 -95512 9740
rect -27644 9274 -27112 9740
rect -96044 7274 -95512 7740
rect -27644 7274 -27112 7740
rect -96044 5274 -95512 5740
rect -27644 5274 -27112 5740
rect 1374 5776 1700 6016
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect 6262 5854 6588 6094
rect 11574 5642 11900 5882
rect 17010 5584 17336 5824
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect 26988 3304 27236 3550
rect 27988 3304 28236 3550
rect 28988 3304 29236 3550
rect 29988 3304 30236 3550
rect 30988 3304 31236 3550
rect 32242 3326 32484 3574
rect 32212 2660 32460 2904
rect 27926 930 28126 1128
rect 28182 928 28382 1128
rect 28422 930 28622 1130
rect 28656 928 28830 1128
rect 27926 656 28126 856
rect 27926 422 28126 622
rect 27926 182 28126 382
rect 27924 -48 28124 144
rect 27926 -288 28126 -88
rect 27924 -524 28124 -324
rect 8763 -968 8797 -934
rect 8855 -968 8889 -934
rect 8947 -968 8981 -934
rect 9039 -968 9073 -934
rect 9131 -968 9165 -934
rect 9223 -968 9257 -934
rect 9315 -968 9349 -934
rect 9407 -968 9441 -934
rect 9499 -968 9533 -934
rect 9591 -968 9625 -934
rect 9683 -968 9717 -934
rect 9775 -968 9809 -934
rect 9867 -968 9901 -934
rect 9959 -968 9993 -934
rect 10051 -968 10085 -934
rect 10143 -968 10177 -934
rect 10235 -968 10269 -934
rect 10327 -968 10361 -934
rect 10419 -968 10453 -934
rect 10511 -968 10545 -934
rect 10603 -968 10637 -934
rect 10695 -968 10729 -934
rect 10787 -968 10821 -934
rect 11229 -968 11263 -934
rect 11321 -968 11355 -934
rect 11413 -968 11447 -934
rect 11505 -968 11539 -934
rect 11597 -968 11631 -934
rect 11689 -968 11723 -934
rect 11781 -968 11815 -934
rect 11873 -968 11907 -934
rect 11965 -968 11999 -934
rect 12057 -968 12091 -934
rect 12149 -968 12183 -934
rect 12241 -968 12275 -934
rect 12333 -968 12367 -934
rect 12425 -968 12459 -934
rect 12517 -968 12551 -934
rect 12609 -968 12643 -934
rect 12701 -968 12735 -934
rect 12793 -968 12827 -934
rect 12885 -968 12919 -934
rect 12977 -968 13011 -934
rect 13069 -968 13103 -934
rect 13161 -968 13195 -934
rect 13253 -968 13287 -934
rect 28042 -936 28242 -736
rect 28348 -938 28548 -738
rect 28628 -938 28790 -738
rect 10181 -1770 10215 -1736
rect 10273 -1770 10307 -1736
rect 10365 -1770 10399 -1736
rect 11229 -1769 11263 -1735
rect 11321 -1769 11355 -1735
rect 11413 -1769 11447 -1735
rect 11505 -1769 11539 -1735
rect 11597 -1769 11631 -1735
rect 11689 -1769 11723 -1735
rect 11781 -1769 11815 -1735
rect 11873 -1769 11907 -1735
rect 11965 -1769 11999 -1735
rect 12057 -1769 12091 -1735
rect 12149 -1769 12183 -1735
rect 12241 -1769 12275 -1735
rect 12333 -1769 12367 -1735
rect 12425 -1769 12459 -1735
rect 12517 -1769 12551 -1735
rect 12609 -1769 12643 -1735
rect 12701 -1769 12735 -1735
rect 12793 -1769 12827 -1735
rect 12885 -1769 12919 -1735
rect 12977 -1769 13011 -1735
rect 13069 -1769 13103 -1735
rect 13161 -1769 13195 -1735
rect 13253 -1769 13287 -1735
rect -9129 -4238 -9095 -4204
rect -9037 -4238 -9003 -4204
rect -8945 -4238 -8911 -4204
rect -8853 -4238 -8819 -4204
rect -8761 -4238 -8727 -4204
rect -8669 -4238 -8635 -4204
rect -8577 -4238 -8543 -4204
rect -8485 -4238 -8451 -4204
rect -8393 -4238 -8359 -4204
rect -8301 -4238 -8267 -4204
rect -8209 -4238 -8175 -4204
rect -8117 -4238 -8083 -4204
rect -8025 -4238 -7991 -4204
rect -7933 -4238 -7899 -4204
rect -7841 -4238 -7807 -4204
rect -7749 -4238 -7715 -4204
rect -7657 -4238 -7623 -4204
rect -7565 -4238 -7531 -4204
rect -7473 -4238 -7439 -4204
rect -7381 -4238 -7347 -4204
rect -7289 -4238 -7255 -4204
rect -7197 -4238 -7163 -4204
rect -7105 -4238 -7071 -4204
rect -7013 -4238 -6979 -4204
rect -6921 -4238 -6887 -4204
rect -6829 -4238 -6795 -4204
rect -6737 -4238 -6703 -4204
rect -6645 -4238 -6611 -4204
rect -6553 -4238 -6519 -4204
rect -6461 -4238 -6427 -4204
rect -6369 -4238 -6335 -4204
rect -6277 -4238 -6243 -4204
rect -6185 -4238 -6151 -4204
rect -6093 -4238 -6059 -4204
rect -6001 -4238 -5967 -4204
rect -5909 -4238 -5875 -4204
rect -5817 -4238 -5783 -4204
rect -5725 -4238 -5691 -4204
rect -5633 -4238 -5599 -4204
rect -5541 -4238 -5507 -4204
rect -5449 -4238 -5415 -4204
rect -5357 -4238 -5323 -4204
rect -5265 -4238 -5231 -4204
rect -5173 -4238 -5139 -4204
rect -5081 -4238 -5047 -4204
rect -4989 -4238 -4955 -4204
rect -4897 -4238 -4863 -4204
rect -4805 -4238 -4771 -4204
rect -4713 -4238 -4679 -4204
rect -4621 -4238 -4587 -4204
rect -4529 -4238 -4495 -4204
rect -4437 -4238 -4403 -4204
rect -4345 -4238 -4311 -4204
rect -4253 -4238 -4219 -4204
rect -4161 -4238 -4127 -4204
rect -4069 -4238 -4035 -4204
rect -3977 -4238 -3943 -4204
rect -3885 -4238 -3851 -4204
rect -3793 -4238 -3759 -4204
rect -3701 -4238 -3667 -4204
rect -3609 -4238 -3575 -4204
rect -3517 -4238 -3483 -4204
rect -3425 -4238 -3391 -4204
rect -3333 -4238 -3299 -4204
rect -3241 -4238 -3207 -4204
rect -3149 -4238 -3115 -4204
rect -3057 -4238 -3023 -4204
rect -2965 -4238 -2931 -4204
rect -2873 -4238 -2839 -4204
rect -2781 -4238 -2747 -4204
rect -2689 -4238 -2655 -4204
rect -2597 -4238 -2563 -4204
rect -2505 -4238 -2471 -4204
rect -2413 -4238 -2379 -4204
rect -2321 -4238 -2287 -4204
rect -2229 -4238 -2195 -4204
rect -2137 -4238 -2103 -4204
rect -2045 -4238 -2011 -4204
rect -1953 -4238 -1919 -4204
rect -1861 -4238 -1827 -4204
rect -1769 -4238 -1735 -4204
rect -1677 -4238 -1643 -4204
rect -1585 -4238 -1551 -4204
rect -1493 -4238 -1459 -4204
rect -1401 -4238 -1367 -4204
rect -1309 -4238 -1275 -4204
rect -1217 -4238 -1183 -4204
rect -1125 -4238 -1091 -4204
rect -1033 -4238 -999 -4204
rect -941 -4238 -907 -4204
rect -849 -4238 -815 -4204
rect -757 -4238 -723 -4204
rect -665 -4238 -631 -4204
rect -573 -4238 -539 -4204
rect -481 -4238 -447 -4204
rect -389 -4238 -355 -4204
rect -297 -4238 -263 -4204
rect -205 -4238 -171 -4204
rect -113 -4238 -79 -4204
rect -21 -4238 13 -4204
rect 71 -4238 105 -4204
rect 163 -4238 197 -4204
rect 255 -4238 289 -4204
rect 347 -4238 381 -4204
rect 439 -4238 473 -4204
rect 531 -4238 565 -4204
rect 623 -4238 657 -4204
rect 715 -4238 749 -4204
rect 807 -4238 841 -4204
rect 899 -4238 933 -4204
rect 991 -4238 1025 -4204
rect 1083 -4238 1117 -4204
rect 1175 -4238 1209 -4204
rect 1267 -4238 1301 -4204
rect 1359 -4238 1393 -4204
rect 1451 -4238 1485 -4204
rect 1543 -4238 1577 -4204
rect 1635 -4238 1669 -4204
rect 1727 -4238 1761 -4204
rect 1819 -4238 1853 -4204
rect 1911 -4238 1945 -4204
rect 2003 -4238 2037 -4204
rect 2095 -4238 2129 -4204
rect 2187 -4238 2221 -4204
rect 2279 -4238 2313 -4204
rect 2371 -4238 2405 -4204
rect 2463 -4238 2497 -4204
rect 2555 -4238 2589 -4204
rect 2647 -4238 2681 -4204
rect 2739 -4238 2773 -4204
rect 2831 -4238 2865 -4204
rect 2923 -4238 2957 -4204
rect 3015 -4238 3049 -4204
rect 3107 -4238 3141 -4204
rect 3199 -4238 3233 -4204
rect 3291 -4238 3325 -4204
rect 3383 -4238 3417 -4204
rect 3475 -4238 3509 -4204
rect 3567 -4238 3601 -4204
rect 3659 -4238 3693 -4204
rect 3751 -4238 3785 -4204
rect 3843 -4238 3877 -4204
rect 3935 -4238 3969 -4204
rect 4027 -4238 4061 -4204
rect 4119 -4238 4153 -4204
rect 4211 -4238 4245 -4204
rect 4303 -4238 4337 -4204
rect 4395 -4238 4429 -4204
rect 4487 -4238 4521 -4204
rect 4579 -4238 4613 -4204
rect 4671 -4238 4705 -4204
rect 4763 -4238 4797 -4204
rect 4855 -4238 4889 -4204
rect 4947 -4238 4981 -4204
rect 5039 -4238 5073 -4204
rect 5131 -4238 5165 -4204
rect 5223 -4238 5257 -4204
rect 5315 -4238 5349 -4204
rect 5407 -4238 5441 -4204
rect 5499 -4238 5533 -4204
rect 5591 -4238 5625 -4204
rect 5683 -4238 5717 -4204
rect 5775 -4238 5809 -4204
rect 5867 -4238 5901 -4204
rect 5959 -4238 5993 -4204
rect 6051 -4238 6085 -4204
rect 6143 -4238 6177 -4204
rect 6235 -4238 6269 -4204
rect 6327 -4238 6361 -4204
rect 6419 -4238 6453 -4204
rect 6511 -4238 6545 -4204
rect 6603 -4238 6637 -4204
rect 6695 -4238 6729 -4204
rect 6787 -4238 6821 -4204
rect 6879 -4238 6913 -4204
rect 6971 -4238 7005 -4204
rect 7063 -4238 7097 -4204
rect 7155 -4238 7189 -4204
rect 7247 -4238 7281 -4204
rect 7339 -4238 7373 -4204
rect 7431 -4238 7465 -4204
rect 7523 -4238 7557 -4204
rect 7615 -4238 7649 -4204
rect 7707 -4238 7741 -4204
rect 7799 -4238 7833 -4204
rect 7891 -4238 7925 -4204
rect 7983 -4238 8017 -4204
rect 8075 -4238 8109 -4204
rect 8167 -4238 8201 -4204
rect 8259 -4238 8293 -4204
rect 8351 -4238 8385 -4204
rect 8443 -4238 8477 -4204
rect 8535 -4238 8569 -4204
rect 8627 -4238 8661 -4204
rect 8719 -4238 8753 -4204
rect 8811 -4238 8845 -4204
rect 8903 -4238 8937 -4204
rect 8995 -4238 9029 -4204
rect 9087 -4238 9121 -4204
rect 9179 -4238 9213 -4204
rect 9271 -4238 9305 -4204
rect 9363 -4238 9397 -4204
rect 9455 -4238 9489 -4204
rect 9547 -4238 9581 -4204
rect 9639 -4238 9673 -4204
rect 9731 -4238 9765 -4204
rect 9823 -4238 9857 -4204
rect 9915 -4238 9949 -4204
rect 10007 -4238 10041 -4204
rect 10099 -4238 10133 -4204
rect 10191 -4238 10225 -4204
rect 10283 -4238 10317 -4204
rect 10375 -4238 10409 -4204
rect 10467 -4238 10501 -4204
rect 10559 -4238 10593 -4204
rect 10651 -4238 10685 -4204
rect 10743 -4238 10777 -4204
rect 10835 -4238 10869 -4204
rect 10927 -4238 10961 -4204
rect 11019 -4238 11053 -4204
rect 11111 -4238 11145 -4204
rect 11203 -4238 11237 -4204
rect 11295 -4238 11329 -4204
rect 11387 -4238 11421 -4204
rect 11479 -4238 11513 -4204
rect 11571 -4238 11605 -4204
rect 11663 -4238 11697 -4204
rect 11755 -4238 11789 -4204
rect 11847 -4238 11881 -4204
rect 11939 -4238 11973 -4204
rect 12031 -4238 12065 -4204
rect 12123 -4238 12157 -4204
rect 12215 -4238 12249 -4204
rect 12307 -4238 12341 -4204
rect 12399 -4238 12433 -4204
rect 12491 -4238 12525 -4204
rect 12583 -4238 12617 -4204
rect 12675 -4238 12709 -4204
rect 12767 -4238 12801 -4204
rect 12859 -4238 12893 -4204
rect 12951 -4238 12985 -4204
rect 13043 -4238 13077 -4204
rect 13135 -4238 13169 -4204
rect 13227 -4238 13261 -4204
rect 13319 -4238 13353 -4204
rect 13411 -4238 13445 -4204
rect 13503 -4238 13537 -4204
rect 13595 -4238 13629 -4204
rect 13687 -4238 13721 -4204
rect 13779 -4238 13813 -4204
rect 13871 -4238 13905 -4204
rect 13963 -4238 13997 -4204
rect 14055 -4238 14089 -4204
rect 14147 -4238 14181 -4204
rect 14239 -4238 14273 -4204
rect 14331 -4238 14365 -4204
rect 14423 -4238 14457 -4204
rect 14515 -4238 14549 -4204
rect 14607 -4238 14641 -4204
rect 14699 -4238 14733 -4204
rect 14791 -4238 14825 -4204
rect 14883 -4238 14917 -4204
rect 14975 -4238 15009 -4204
rect 15067 -4238 15101 -4204
rect 15159 -4238 15193 -4204
rect 15251 -4238 15285 -4204
rect 15343 -4238 15377 -4204
rect 15435 -4238 15469 -4204
rect 15527 -4238 15561 -4204
rect 15619 -4238 15653 -4204
rect 15711 -4238 15745 -4204
rect 15803 -4238 15837 -4204
rect 15895 -4238 15929 -4204
rect 15987 -4238 16021 -4204
rect 16079 -4238 16113 -4204
rect 16171 -4238 16205 -4204
rect 16263 -4238 16297 -4204
rect 16355 -4238 16389 -4204
rect 16447 -4238 16481 -4204
rect 16539 -4238 16573 -4204
rect 16631 -4238 16665 -4204
rect 16723 -4238 16757 -4204
rect 16815 -4238 16849 -4204
rect 16907 -4238 16941 -4204
rect 16999 -4238 17033 -4204
rect 17091 -4238 17125 -4204
rect 17183 -4238 17217 -4204
rect 17275 -4238 17309 -4204
rect 17367 -4238 17401 -4204
rect 17459 -4238 17493 -4204
rect 17551 -4238 17585 -4204
rect 17643 -4238 17677 -4204
rect 17735 -4238 17769 -4204
rect 17827 -4238 17861 -4204
rect 17919 -4238 17953 -4204
rect 18011 -4238 18045 -4204
rect 18103 -4238 18137 -4204
rect 18195 -4238 18229 -4204
rect 18287 -4238 18321 -4204
rect 18379 -4238 18413 -4204
rect 18471 -4238 18505 -4204
rect 18563 -4238 18597 -4204
rect 18655 -4238 18689 -4204
rect 18747 -4238 18781 -4204
rect 18839 -4238 18873 -4204
rect 18931 -4238 18965 -4204
rect 19023 -4238 19057 -4204
rect 19115 -4238 19149 -4204
rect 19207 -4238 19241 -4204
rect 19299 -4238 19333 -4204
rect 19391 -4238 19425 -4204
rect 19483 -4238 19517 -4204
rect 19575 -4238 19609 -4204
rect 19667 -4238 19701 -4204
rect 19759 -4238 19793 -4204
rect 19851 -4238 19885 -4204
rect 19943 -4238 19977 -4204
rect 20035 -4238 20069 -4204
rect 20127 -4238 20161 -4204
rect 20219 -4238 20253 -4204
rect 20311 -4238 20345 -4204
rect 20403 -4238 20437 -4204
rect 20495 -4238 20529 -4204
rect 20587 -4238 20621 -4204
rect 20679 -4238 20713 -4204
rect 20771 -4238 20805 -4204
rect 20863 -4238 20897 -4204
rect 20955 -4238 20989 -4204
rect 21047 -4238 21081 -4204
rect 21139 -4238 21173 -4204
rect 21231 -4238 21265 -4204
rect 21323 -4238 21357 -4204
rect 21415 -4238 21449 -4204
rect 21507 -4238 21541 -4204
rect 21599 -4238 21633 -4204
rect 21691 -4238 21725 -4204
rect 21783 -4238 21817 -4204
rect 21875 -4238 21909 -4204
rect 21967 -4238 22001 -4204
rect 22059 -4238 22093 -4204
rect 22151 -4238 22185 -4204
rect 22243 -4238 22277 -4204
rect 22335 -4238 22369 -4204
rect 22427 -4238 22461 -4204
rect 22519 -4238 22553 -4204
rect 22611 -4238 22645 -4204
rect 22703 -4238 22737 -4204
rect 22795 -4238 22829 -4204
rect 22887 -4238 22921 -4204
rect 22979 -4238 23013 -4204
rect 23071 -4238 23105 -4204
rect 23163 -4238 23197 -4204
rect 23255 -4238 23289 -4204
rect 23347 -4238 23381 -4204
rect 23439 -4238 23473 -4204
rect 23531 -4238 23565 -4204
rect 23623 -4238 23657 -4204
rect 23715 -4238 23749 -4204
rect 23807 -4238 23841 -4204
rect 23899 -4238 23933 -4204
rect 23991 -4238 24025 -4204
rect 24083 -4238 24117 -4204
rect 24175 -4238 24209 -4204
rect 24267 -4238 24301 -4204
rect 24359 -4238 24393 -4204
rect 24451 -4238 24485 -4204
rect 24543 -4238 24577 -4204
rect 24635 -4238 24669 -4204
rect 24727 -4238 24761 -4204
rect 24819 -4238 24853 -4204
rect 24911 -4238 24945 -4204
rect 25003 -4238 25037 -4204
rect 25095 -4238 25129 -4204
rect 25187 -4238 25221 -4204
rect 25279 -4238 25313 -4204
rect 25371 -4238 25405 -4204
rect 25463 -4238 25497 -4204
rect 25555 -4238 25589 -4204
rect 25647 -4238 25681 -4204
rect 25739 -4238 25773 -4204
rect 25831 -4238 25865 -4204
rect 25923 -4238 25957 -4204
rect 26015 -4238 26049 -4204
rect 26107 -4238 26141 -4204
rect 26199 -4238 26233 -4204
rect 26291 -4238 26325 -4204
rect 26383 -4238 26417 -4204
rect 26475 -4238 26509 -4204
rect 26567 -4238 26601 -4204
rect 26659 -4238 26693 -4204
rect 26751 -4238 26785 -4204
rect 26843 -4238 26877 -4204
rect 26935 -4238 26969 -4204
rect 27027 -4238 27061 -4204
rect 27119 -4238 27153 -4204
rect 27211 -4238 27245 -4204
rect 27303 -4238 27337 -4204
rect 27395 -4238 27429 -4204
rect 27487 -4238 27521 -4204
rect 27579 -4238 27613 -4204
rect 27671 -4238 27705 -4204
rect 27763 -4238 27797 -4204
rect 27855 -4238 27889 -4204
rect 27947 -4238 27981 -4204
rect 28039 -4238 28073 -4204
rect 28131 -4238 28165 -4204
rect 28223 -4238 28257 -4204
rect 28315 -4238 28349 -4204
rect 28407 -4238 28441 -4204
rect 28499 -4238 28533 -4204
rect 28591 -4238 28625 -4204
rect 28683 -4238 28717 -4204
rect 28775 -4238 28809 -4204
rect 28867 -4238 28901 -4204
rect 28959 -4238 28993 -4204
rect 29051 -4238 29085 -4204
rect 29143 -4238 29177 -4204
rect 29235 -4238 29269 -4204
rect 29327 -4238 29361 -4204
rect 29419 -4238 29453 -4204
rect 29511 -4238 29545 -4204
rect 29603 -4238 29637 -4204
rect 29695 -4238 29729 -4204
rect 29787 -4238 29821 -4204
rect 29879 -4238 29913 -4204
rect 29971 -4238 30005 -4204
rect 30063 -4238 30097 -4204
rect 30155 -4238 30189 -4204
rect 30247 -4238 30281 -4204
rect 30339 -4238 30373 -4204
rect 30431 -4238 30465 -4204
rect 30523 -4238 30557 -4204
rect 30615 -4238 30649 -4204
rect 30707 -4238 30741 -4204
rect 30799 -4238 30833 -4204
rect 30891 -4238 30925 -4204
rect 30983 -4238 31017 -4204
rect 31075 -4238 31109 -4204
rect 31167 -4238 31201 -4204
rect 31259 -4238 31293 -4204
rect 31351 -4238 31385 -4204
rect 31443 -4238 31477 -4204
rect 31535 -4238 31569 -4204
rect 31627 -4238 31661 -4204
rect 31719 -4238 31753 -4204
rect 31811 -4238 31845 -4204
rect 31903 -4238 31937 -4204
rect 31995 -4238 32029 -4204
rect 32087 -4238 32121 -4204
rect 32179 -4238 32213 -4204
rect 32271 -4238 32305 -4204
rect 32363 -4238 32397 -4204
rect 32455 -4238 32489 -4204
rect 32547 -4238 32581 -4204
rect 32639 -4238 32673 -4204
rect 32731 -4238 32765 -4204
rect 32823 -4238 32857 -4204
rect 32915 -4238 32949 -4204
rect 33007 -4238 33041 -4204
rect 33099 -4238 33133 -4204
rect 10166 -7474 10794 -7379
rect 12946 -7478 13574 -7383
rect 9055 -8937 9192 -8675
rect 16474 -8956 16611 -8694
rect 9014 -14503 9151 -14241
rect 16428 -14510 16565 -14248
rect 8973 -20385 9109 -20124
rect 16248 -19893 16450 -19579
rect 16510 -19811 16566 -19749
rect 16900 -19813 16956 -19751
<< poly >>
rect -94172 20649 -93356 20665
rect -94172 20632 -94156 20649
rect -94564 20615 -94156 20632
rect -93372 20632 -93356 20649
rect -92514 20649 -91698 20665
rect -92514 20632 -92498 20649
rect -93372 20615 -92964 20632
rect -94564 20568 -92964 20615
rect -92906 20615 -92498 20632
rect -91714 20632 -91698 20649
rect -90856 20649 -90040 20665
rect -90856 20632 -90840 20649
rect -91714 20615 -91306 20632
rect -92906 20568 -91306 20615
rect -91248 20615 -90840 20632
rect -90056 20632 -90040 20649
rect -89198 20649 -88382 20665
rect -89198 20632 -89182 20649
rect -90056 20615 -89648 20632
rect -91248 20568 -89648 20615
rect -89590 20615 -89182 20632
rect -88398 20632 -88382 20649
rect -87540 20649 -86724 20665
rect -87540 20632 -87524 20649
rect -88398 20615 -87990 20632
rect -89590 20568 -87990 20615
rect -87932 20615 -87524 20632
rect -86740 20632 -86724 20649
rect -85882 20649 -85066 20665
rect -85882 20632 -85866 20649
rect -86740 20615 -86332 20632
rect -87932 20568 -86332 20615
rect -86274 20615 -85866 20632
rect -85082 20632 -85066 20649
rect -84224 20649 -83408 20665
rect -84224 20632 -84208 20649
rect -85082 20615 -84674 20632
rect -86274 20568 -84674 20615
rect -84616 20615 -84208 20632
rect -83424 20632 -83408 20649
rect -82566 20649 -81750 20665
rect -82566 20632 -82550 20649
rect -83424 20615 -83016 20632
rect -84616 20568 -83016 20615
rect -82958 20615 -82550 20632
rect -81766 20632 -81750 20649
rect -80908 20649 -80092 20665
rect -80908 20632 -80892 20649
rect -81766 20615 -81358 20632
rect -82958 20568 -81358 20615
rect -81300 20615 -80892 20632
rect -80108 20632 -80092 20649
rect -79250 20649 -78434 20665
rect -79250 20632 -79234 20649
rect -80108 20615 -79700 20632
rect -81300 20568 -79700 20615
rect -79642 20615 -79234 20632
rect -78450 20632 -78434 20649
rect -77592 20649 -76776 20665
rect -77592 20632 -77576 20649
rect -78450 20615 -78042 20632
rect -79642 20568 -78042 20615
rect -77984 20615 -77576 20632
rect -76792 20632 -76776 20649
rect -75934 20649 -75118 20665
rect -75934 20632 -75918 20649
rect -76792 20615 -76384 20632
rect -77984 20568 -76384 20615
rect -76326 20615 -75918 20632
rect -75134 20632 -75118 20649
rect -74276 20649 -73460 20665
rect -74276 20632 -74260 20649
rect -75134 20615 -74726 20632
rect -76326 20568 -74726 20615
rect -74668 20615 -74260 20632
rect -73476 20632 -73460 20649
rect -72618 20649 -71802 20665
rect -72618 20632 -72602 20649
rect -73476 20615 -73068 20632
rect -74668 20568 -73068 20615
rect -73010 20615 -72602 20632
rect -71818 20632 -71802 20649
rect -70960 20649 -70144 20665
rect -70960 20632 -70944 20649
rect -71818 20615 -71410 20632
rect -73010 20568 -71410 20615
rect -71352 20615 -70944 20632
rect -70160 20632 -70144 20649
rect -69302 20649 -68486 20665
rect -69302 20632 -69286 20649
rect -70160 20615 -69752 20632
rect -71352 20568 -69752 20615
rect -69694 20615 -69286 20632
rect -68502 20632 -68486 20649
rect -67644 20649 -66828 20665
rect -67644 20632 -67628 20649
rect -68502 20615 -68094 20632
rect -69694 20568 -68094 20615
rect -68036 20615 -67628 20632
rect -66844 20632 -66828 20649
rect -65986 20649 -65170 20665
rect -65986 20632 -65970 20649
rect -66844 20615 -66436 20632
rect -68036 20568 -66436 20615
rect -66378 20615 -65970 20632
rect -65186 20632 -65170 20649
rect -64328 20649 -63512 20665
rect -64328 20632 -64312 20649
rect -65186 20615 -64778 20632
rect -66378 20568 -64778 20615
rect -64720 20615 -64312 20632
rect -63528 20632 -63512 20649
rect -62670 20649 -61854 20665
rect -62670 20632 -62654 20649
rect -63528 20615 -63120 20632
rect -64720 20568 -63120 20615
rect -63062 20615 -62654 20632
rect -61870 20632 -61854 20649
rect -61012 20649 -60196 20665
rect -61012 20632 -60996 20649
rect -61870 20615 -61462 20632
rect -63062 20568 -61462 20615
rect -61404 20615 -60996 20632
rect -60212 20632 -60196 20649
rect -59354 20649 -58538 20665
rect -59354 20632 -59338 20649
rect -60212 20615 -59804 20632
rect -61404 20568 -59804 20615
rect -59746 20615 -59338 20632
rect -58554 20632 -58538 20649
rect -57696 20649 -56880 20665
rect -57696 20632 -57680 20649
rect -58554 20615 -58146 20632
rect -59746 20568 -58146 20615
rect -58088 20615 -57680 20632
rect -56896 20632 -56880 20649
rect -56038 20649 -55222 20665
rect -56038 20632 -56022 20649
rect -56896 20615 -56488 20632
rect -58088 20568 -56488 20615
rect -56430 20615 -56022 20632
rect -55238 20632 -55222 20649
rect -54380 20649 -53564 20665
rect -54380 20632 -54364 20649
rect -55238 20615 -54830 20632
rect -56430 20568 -54830 20615
rect -54772 20615 -54364 20632
rect -53580 20632 -53564 20649
rect -52722 20649 -51906 20665
rect -52722 20632 -52706 20649
rect -53580 20615 -53172 20632
rect -54772 20568 -53172 20615
rect -53114 20615 -52706 20632
rect -51922 20632 -51906 20649
rect -51064 20649 -50248 20665
rect -51064 20632 -51048 20649
rect -51922 20615 -51514 20632
rect -53114 20568 -51514 20615
rect -51456 20615 -51048 20632
rect -50264 20632 -50248 20649
rect -49406 20649 -48590 20665
rect -49406 20632 -49390 20649
rect -50264 20615 -49856 20632
rect -51456 20568 -49856 20615
rect -49798 20615 -49390 20632
rect -48606 20632 -48590 20649
rect -47748 20649 -46932 20665
rect -47748 20632 -47732 20649
rect -48606 20615 -48198 20632
rect -49798 20568 -48198 20615
rect -48140 20615 -47732 20632
rect -46948 20632 -46932 20649
rect -46090 20649 -45274 20665
rect -46090 20632 -46074 20649
rect -46948 20615 -46540 20632
rect -48140 20568 -46540 20615
rect -46482 20615 -46074 20632
rect -45290 20632 -45274 20649
rect -44432 20649 -43616 20665
rect -44432 20632 -44416 20649
rect -45290 20615 -44882 20632
rect -46482 20568 -44882 20615
rect -44824 20615 -44416 20632
rect -43632 20632 -43616 20649
rect -42774 20649 -41958 20665
rect -42774 20632 -42758 20649
rect -43632 20615 -43224 20632
rect -44824 20568 -43224 20615
rect -43166 20615 -42758 20632
rect -41974 20632 -41958 20649
rect -41116 20649 -40300 20665
rect -41116 20632 -41100 20649
rect -41974 20615 -41566 20632
rect -43166 20568 -41566 20615
rect -41508 20615 -41100 20632
rect -40316 20632 -40300 20649
rect -39458 20649 -38642 20665
rect -39458 20632 -39442 20649
rect -40316 20615 -39908 20632
rect -41508 20568 -39908 20615
rect -39850 20615 -39442 20632
rect -38658 20632 -38642 20649
rect -37800 20649 -36984 20665
rect -37800 20632 -37784 20649
rect -38658 20615 -38250 20632
rect -39850 20568 -38250 20615
rect -38192 20615 -37784 20632
rect -37000 20632 -36984 20649
rect -36142 20649 -35326 20665
rect -36142 20632 -36126 20649
rect -37000 20615 -36592 20632
rect -38192 20568 -36592 20615
rect -36534 20615 -36126 20632
rect -35342 20632 -35326 20649
rect -34484 20649 -33668 20665
rect -34484 20632 -34468 20649
rect -35342 20615 -34934 20632
rect -36534 20568 -34934 20615
rect -34876 20615 -34468 20632
rect -33684 20632 -33668 20649
rect -32826 20649 -32010 20665
rect -32826 20632 -32810 20649
rect -33684 20615 -33276 20632
rect -34876 20568 -33276 20615
rect -33218 20615 -32810 20632
rect -32026 20632 -32010 20649
rect -31168 20649 -30352 20665
rect -31168 20632 -31152 20649
rect -32026 20615 -31618 20632
rect -33218 20568 -31618 20615
rect -31560 20615 -31152 20632
rect -30368 20632 -30352 20649
rect -29510 20649 -28694 20665
rect -29510 20632 -29494 20649
rect -30368 20615 -29960 20632
rect -31560 20568 -29960 20615
rect -29902 20615 -29494 20632
rect -28710 20632 -28694 20649
rect -28710 20615 -28302 20632
rect -29902 20568 -28302 20615
rect -94564 19121 -92964 19168
rect -94564 19104 -94156 19121
rect -94172 19087 -94156 19104
rect -93372 19104 -92964 19121
rect -92906 19121 -91306 19168
rect -92906 19104 -92498 19121
rect -93372 19087 -93356 19104
rect -94172 19071 -93356 19087
rect -92514 19087 -92498 19104
rect -91714 19104 -91306 19121
rect -91248 19121 -89648 19168
rect -91248 19104 -90840 19121
rect -91714 19087 -91698 19104
rect -92514 19071 -91698 19087
rect -90856 19087 -90840 19104
rect -90056 19104 -89648 19121
rect -89590 19121 -87990 19168
rect -89590 19104 -89182 19121
rect -90056 19087 -90040 19104
rect -90856 19071 -90040 19087
rect -89198 19087 -89182 19104
rect -88398 19104 -87990 19121
rect -87932 19121 -86332 19168
rect -87932 19104 -87524 19121
rect -88398 19087 -88382 19104
rect -89198 19071 -88382 19087
rect -87540 19087 -87524 19104
rect -86740 19104 -86332 19121
rect -86274 19121 -84674 19168
rect -86274 19104 -85866 19121
rect -86740 19087 -86724 19104
rect -87540 19071 -86724 19087
rect -85882 19087 -85866 19104
rect -85082 19104 -84674 19121
rect -84616 19121 -83016 19168
rect -84616 19104 -84208 19121
rect -85082 19087 -85066 19104
rect -85882 19071 -85066 19087
rect -84224 19087 -84208 19104
rect -83424 19104 -83016 19121
rect -82958 19121 -81358 19168
rect -82958 19104 -82550 19121
rect -83424 19087 -83408 19104
rect -84224 19071 -83408 19087
rect -82566 19087 -82550 19104
rect -81766 19104 -81358 19121
rect -81300 19121 -79700 19168
rect -81300 19104 -80892 19121
rect -81766 19087 -81750 19104
rect -82566 19071 -81750 19087
rect -80908 19087 -80892 19104
rect -80108 19104 -79700 19121
rect -79642 19121 -78042 19168
rect -79642 19104 -79234 19121
rect -80108 19087 -80092 19104
rect -80908 19071 -80092 19087
rect -79250 19087 -79234 19104
rect -78450 19104 -78042 19121
rect -77984 19121 -76384 19168
rect -77984 19104 -77576 19121
rect -78450 19087 -78434 19104
rect -79250 19071 -78434 19087
rect -77592 19087 -77576 19104
rect -76792 19104 -76384 19121
rect -76326 19121 -74726 19168
rect -76326 19104 -75918 19121
rect -76792 19087 -76776 19104
rect -77592 19071 -76776 19087
rect -75934 19087 -75918 19104
rect -75134 19104 -74726 19121
rect -74668 19121 -73068 19168
rect -74668 19104 -74260 19121
rect -75134 19087 -75118 19104
rect -75934 19071 -75118 19087
rect -74276 19087 -74260 19104
rect -73476 19104 -73068 19121
rect -73010 19121 -71410 19168
rect -73010 19104 -72602 19121
rect -73476 19087 -73460 19104
rect -74276 19071 -73460 19087
rect -72618 19087 -72602 19104
rect -71818 19104 -71410 19121
rect -71352 19121 -69752 19168
rect -71352 19104 -70944 19121
rect -71818 19087 -71802 19104
rect -72618 19071 -71802 19087
rect -70960 19087 -70944 19104
rect -70160 19104 -69752 19121
rect -69694 19121 -68094 19168
rect -69694 19104 -69286 19121
rect -70160 19087 -70144 19104
rect -70960 19071 -70144 19087
rect -69302 19087 -69286 19104
rect -68502 19104 -68094 19121
rect -68036 19121 -66436 19168
rect -68036 19104 -67628 19121
rect -68502 19087 -68486 19104
rect -69302 19071 -68486 19087
rect -67644 19087 -67628 19104
rect -66844 19104 -66436 19121
rect -66378 19121 -64778 19168
rect -66378 19104 -65970 19121
rect -66844 19087 -66828 19104
rect -67644 19071 -66828 19087
rect -65986 19087 -65970 19104
rect -65186 19104 -64778 19121
rect -64720 19121 -63120 19168
rect -64720 19104 -64312 19121
rect -65186 19087 -65170 19104
rect -65986 19071 -65170 19087
rect -64328 19087 -64312 19104
rect -63528 19104 -63120 19121
rect -63062 19121 -61462 19168
rect -63062 19104 -62654 19121
rect -63528 19087 -63512 19104
rect -64328 19071 -63512 19087
rect -62670 19087 -62654 19104
rect -61870 19104 -61462 19121
rect -61404 19121 -59804 19168
rect -61404 19104 -60996 19121
rect -61870 19087 -61854 19104
rect -62670 19071 -61854 19087
rect -61012 19087 -60996 19104
rect -60212 19104 -59804 19121
rect -59746 19121 -58146 19168
rect -59746 19104 -59338 19121
rect -60212 19087 -60196 19104
rect -61012 19071 -60196 19087
rect -59354 19087 -59338 19104
rect -58554 19104 -58146 19121
rect -58088 19121 -56488 19168
rect -58088 19104 -57680 19121
rect -58554 19087 -58538 19104
rect -59354 19071 -58538 19087
rect -57696 19087 -57680 19104
rect -56896 19104 -56488 19121
rect -56430 19121 -54830 19168
rect -56430 19104 -56022 19121
rect -56896 19087 -56880 19104
rect -57696 19071 -56880 19087
rect -56038 19087 -56022 19104
rect -55238 19104 -54830 19121
rect -54772 19121 -53172 19168
rect -54772 19104 -54364 19121
rect -55238 19087 -55222 19104
rect -56038 19071 -55222 19087
rect -54380 19087 -54364 19104
rect -53580 19104 -53172 19121
rect -53114 19121 -51514 19168
rect -53114 19104 -52706 19121
rect -53580 19087 -53564 19104
rect -54380 19071 -53564 19087
rect -52722 19087 -52706 19104
rect -51922 19104 -51514 19121
rect -51456 19121 -49856 19168
rect -51456 19104 -51048 19121
rect -51922 19087 -51906 19104
rect -52722 19071 -51906 19087
rect -51064 19087 -51048 19104
rect -50264 19104 -49856 19121
rect -49798 19121 -48198 19168
rect -49798 19104 -49390 19121
rect -50264 19087 -50248 19104
rect -51064 19071 -50248 19087
rect -49406 19087 -49390 19104
rect -48606 19104 -48198 19121
rect -48140 19121 -46540 19168
rect -48140 19104 -47732 19121
rect -48606 19087 -48590 19104
rect -49406 19071 -48590 19087
rect -47748 19087 -47732 19104
rect -46948 19104 -46540 19121
rect -46482 19121 -44882 19168
rect -46482 19104 -46074 19121
rect -46948 19087 -46932 19104
rect -47748 19071 -46932 19087
rect -46090 19087 -46074 19104
rect -45290 19104 -44882 19121
rect -44824 19121 -43224 19168
rect -44824 19104 -44416 19121
rect -45290 19087 -45274 19104
rect -46090 19071 -45274 19087
rect -44432 19087 -44416 19104
rect -43632 19104 -43224 19121
rect -43166 19121 -41566 19168
rect -43166 19104 -42758 19121
rect -43632 19087 -43616 19104
rect -44432 19071 -43616 19087
rect -42774 19087 -42758 19104
rect -41974 19104 -41566 19121
rect -41508 19121 -39908 19168
rect -41508 19104 -41100 19121
rect -41974 19087 -41958 19104
rect -42774 19071 -41958 19087
rect -41116 19087 -41100 19104
rect -40316 19104 -39908 19121
rect -39850 19121 -38250 19168
rect -39850 19104 -39442 19121
rect -40316 19087 -40300 19104
rect -41116 19071 -40300 19087
rect -39458 19087 -39442 19104
rect -38658 19104 -38250 19121
rect -38192 19121 -36592 19168
rect -38192 19104 -37784 19121
rect -38658 19087 -38642 19104
rect -39458 19071 -38642 19087
rect -37800 19087 -37784 19104
rect -37000 19104 -36592 19121
rect -36534 19121 -34934 19168
rect -36534 19104 -36126 19121
rect -37000 19087 -36984 19104
rect -37800 19071 -36984 19087
rect -36142 19087 -36126 19104
rect -35342 19104 -34934 19121
rect -34876 19121 -33276 19168
rect -34876 19104 -34468 19121
rect -35342 19087 -35326 19104
rect -36142 19071 -35326 19087
rect -34484 19087 -34468 19104
rect -33684 19104 -33276 19121
rect -33218 19121 -31618 19168
rect -33218 19104 -32810 19121
rect -33684 19087 -33668 19104
rect -34484 19071 -33668 19087
rect -32826 19087 -32810 19104
rect -32026 19104 -31618 19121
rect -31560 19121 -29960 19168
rect -31560 19104 -31152 19121
rect -32026 19087 -32010 19104
rect -32826 19071 -32010 19087
rect -31168 19087 -31152 19104
rect -30368 19104 -29960 19121
rect -29902 19121 -28302 19168
rect -29902 19104 -29494 19121
rect -30368 19087 -30352 19104
rect -31168 19071 -30352 19087
rect -29510 19087 -29494 19104
rect -28710 19104 -28302 19121
rect -28710 19087 -28694 19104
rect -29510 19071 -28694 19087
rect -94172 19013 -93356 19029
rect -94172 18996 -94156 19013
rect -94564 18979 -94156 18996
rect -93372 18996 -93356 19013
rect -92514 19013 -91698 19029
rect -92514 18996 -92498 19013
rect -93372 18979 -92964 18996
rect -94564 18932 -92964 18979
rect -92906 18979 -92498 18996
rect -91714 18996 -91698 19013
rect -90856 19013 -90040 19029
rect -90856 18996 -90840 19013
rect -91714 18979 -91306 18996
rect -92906 18932 -91306 18979
rect -91248 18979 -90840 18996
rect -90056 18996 -90040 19013
rect -89198 19013 -88382 19029
rect -89198 18996 -89182 19013
rect -90056 18979 -89648 18996
rect -91248 18932 -89648 18979
rect -89590 18979 -89182 18996
rect -88398 18996 -88382 19013
rect -87540 19013 -86724 19029
rect -87540 18996 -87524 19013
rect -88398 18979 -87990 18996
rect -89590 18932 -87990 18979
rect -87932 18979 -87524 18996
rect -86740 18996 -86724 19013
rect -85882 19013 -85066 19029
rect -85882 18996 -85866 19013
rect -86740 18979 -86332 18996
rect -87932 18932 -86332 18979
rect -86274 18979 -85866 18996
rect -85082 18996 -85066 19013
rect -84224 19013 -83408 19029
rect -84224 18996 -84208 19013
rect -85082 18979 -84674 18996
rect -86274 18932 -84674 18979
rect -84616 18979 -84208 18996
rect -83424 18996 -83408 19013
rect -82566 19013 -81750 19029
rect -82566 18996 -82550 19013
rect -83424 18979 -83016 18996
rect -84616 18932 -83016 18979
rect -82958 18979 -82550 18996
rect -81766 18996 -81750 19013
rect -80908 19013 -80092 19029
rect -80908 18996 -80892 19013
rect -81766 18979 -81358 18996
rect -82958 18932 -81358 18979
rect -81300 18979 -80892 18996
rect -80108 18996 -80092 19013
rect -79250 19013 -78434 19029
rect -79250 18996 -79234 19013
rect -80108 18979 -79700 18996
rect -81300 18932 -79700 18979
rect -79642 18979 -79234 18996
rect -78450 18996 -78434 19013
rect -77592 19013 -76776 19029
rect -77592 18996 -77576 19013
rect -78450 18979 -78042 18996
rect -79642 18932 -78042 18979
rect -77984 18979 -77576 18996
rect -76792 18996 -76776 19013
rect -75934 19013 -75118 19029
rect -75934 18996 -75918 19013
rect -76792 18979 -76384 18996
rect -77984 18932 -76384 18979
rect -76326 18979 -75918 18996
rect -75134 18996 -75118 19013
rect -74276 19013 -73460 19029
rect -74276 18996 -74260 19013
rect -75134 18979 -74726 18996
rect -76326 18932 -74726 18979
rect -74668 18979 -74260 18996
rect -73476 18996 -73460 19013
rect -72618 19013 -71802 19029
rect -72618 18996 -72602 19013
rect -73476 18979 -73068 18996
rect -74668 18932 -73068 18979
rect -73010 18979 -72602 18996
rect -71818 18996 -71802 19013
rect -70960 19013 -70144 19029
rect -70960 18996 -70944 19013
rect -71818 18979 -71410 18996
rect -73010 18932 -71410 18979
rect -71352 18979 -70944 18996
rect -70160 18996 -70144 19013
rect -69302 19013 -68486 19029
rect -69302 18996 -69286 19013
rect -70160 18979 -69752 18996
rect -71352 18932 -69752 18979
rect -69694 18979 -69286 18996
rect -68502 18996 -68486 19013
rect -67644 19013 -66828 19029
rect -67644 18996 -67628 19013
rect -68502 18979 -68094 18996
rect -69694 18932 -68094 18979
rect -68036 18979 -67628 18996
rect -66844 18996 -66828 19013
rect -65986 19013 -65170 19029
rect -65986 18996 -65970 19013
rect -66844 18979 -66436 18996
rect -68036 18932 -66436 18979
rect -66378 18979 -65970 18996
rect -65186 18996 -65170 19013
rect -64328 19013 -63512 19029
rect -64328 18996 -64312 19013
rect -65186 18979 -64778 18996
rect -66378 18932 -64778 18979
rect -64720 18979 -64312 18996
rect -63528 18996 -63512 19013
rect -62670 19013 -61854 19029
rect -62670 18996 -62654 19013
rect -63528 18979 -63120 18996
rect -64720 18932 -63120 18979
rect -63062 18979 -62654 18996
rect -61870 18996 -61854 19013
rect -61012 19013 -60196 19029
rect -61012 18996 -60996 19013
rect -61870 18979 -61462 18996
rect -63062 18932 -61462 18979
rect -61404 18979 -60996 18996
rect -60212 18996 -60196 19013
rect -59354 19013 -58538 19029
rect -59354 18996 -59338 19013
rect -60212 18979 -59804 18996
rect -61404 18932 -59804 18979
rect -59746 18979 -59338 18996
rect -58554 18996 -58538 19013
rect -57696 19013 -56880 19029
rect -57696 18996 -57680 19013
rect -58554 18979 -58146 18996
rect -59746 18932 -58146 18979
rect -58088 18979 -57680 18996
rect -56896 18996 -56880 19013
rect -56038 19013 -55222 19029
rect -56038 18996 -56022 19013
rect -56896 18979 -56488 18996
rect -58088 18932 -56488 18979
rect -56430 18979 -56022 18996
rect -55238 18996 -55222 19013
rect -54380 19013 -53564 19029
rect -54380 18996 -54364 19013
rect -55238 18979 -54830 18996
rect -56430 18932 -54830 18979
rect -54772 18979 -54364 18996
rect -53580 18996 -53564 19013
rect -52722 19013 -51906 19029
rect -52722 18996 -52706 19013
rect -53580 18979 -53172 18996
rect -54772 18932 -53172 18979
rect -53114 18979 -52706 18996
rect -51922 18996 -51906 19013
rect -51064 19013 -50248 19029
rect -51064 18996 -51048 19013
rect -51922 18979 -51514 18996
rect -53114 18932 -51514 18979
rect -51456 18979 -51048 18996
rect -50264 18996 -50248 19013
rect -49406 19013 -48590 19029
rect -49406 18996 -49390 19013
rect -50264 18979 -49856 18996
rect -51456 18932 -49856 18979
rect -49798 18979 -49390 18996
rect -48606 18996 -48590 19013
rect -47748 19013 -46932 19029
rect -47748 18996 -47732 19013
rect -48606 18979 -48198 18996
rect -49798 18932 -48198 18979
rect -48140 18979 -47732 18996
rect -46948 18996 -46932 19013
rect -46090 19013 -45274 19029
rect -46090 18996 -46074 19013
rect -46948 18979 -46540 18996
rect -48140 18932 -46540 18979
rect -46482 18979 -46074 18996
rect -45290 18996 -45274 19013
rect -44432 19013 -43616 19029
rect -44432 18996 -44416 19013
rect -45290 18979 -44882 18996
rect -46482 18932 -44882 18979
rect -44824 18979 -44416 18996
rect -43632 18996 -43616 19013
rect -42774 19013 -41958 19029
rect -42774 18996 -42758 19013
rect -43632 18979 -43224 18996
rect -44824 18932 -43224 18979
rect -43166 18979 -42758 18996
rect -41974 18996 -41958 19013
rect -41116 19013 -40300 19029
rect -41116 18996 -41100 19013
rect -41974 18979 -41566 18996
rect -43166 18932 -41566 18979
rect -41508 18979 -41100 18996
rect -40316 18996 -40300 19013
rect -39458 19013 -38642 19029
rect -39458 18996 -39442 19013
rect -40316 18979 -39908 18996
rect -41508 18932 -39908 18979
rect -39850 18979 -39442 18996
rect -38658 18996 -38642 19013
rect -37800 19013 -36984 19029
rect -37800 18996 -37784 19013
rect -38658 18979 -38250 18996
rect -39850 18932 -38250 18979
rect -38192 18979 -37784 18996
rect -37000 18996 -36984 19013
rect -36142 19013 -35326 19029
rect -36142 18996 -36126 19013
rect -37000 18979 -36592 18996
rect -38192 18932 -36592 18979
rect -36534 18979 -36126 18996
rect -35342 18996 -35326 19013
rect -34484 19013 -33668 19029
rect -34484 18996 -34468 19013
rect -35342 18979 -34934 18996
rect -36534 18932 -34934 18979
rect -34876 18979 -34468 18996
rect -33684 18996 -33668 19013
rect -32826 19013 -32010 19029
rect -32826 18996 -32810 19013
rect -33684 18979 -33276 18996
rect -34876 18932 -33276 18979
rect -33218 18979 -32810 18996
rect -32026 18996 -32010 19013
rect -31168 19013 -30352 19029
rect -31168 18996 -31152 19013
rect -32026 18979 -31618 18996
rect -33218 18932 -31618 18979
rect -31560 18979 -31152 18996
rect -30368 18996 -30352 19013
rect -29510 19013 -28694 19029
rect -29510 18996 -29494 19013
rect -30368 18979 -29960 18996
rect -31560 18932 -29960 18979
rect -29902 18979 -29494 18996
rect -28710 18996 -28694 19013
rect -28710 18979 -28302 18996
rect -29902 18932 -28302 18979
rect -94564 17485 -92964 17532
rect -94564 17468 -94156 17485
rect -94172 17451 -94156 17468
rect -93372 17468 -92964 17485
rect -92906 17485 -91306 17532
rect -92906 17468 -92498 17485
rect -93372 17451 -93356 17468
rect -94172 17435 -93356 17451
rect -92514 17451 -92498 17468
rect -91714 17468 -91306 17485
rect -91248 17485 -89648 17532
rect -91248 17468 -90840 17485
rect -91714 17451 -91698 17468
rect -92514 17435 -91698 17451
rect -90856 17451 -90840 17468
rect -90056 17468 -89648 17485
rect -89590 17485 -87990 17532
rect -89590 17468 -89182 17485
rect -90056 17451 -90040 17468
rect -90856 17435 -90040 17451
rect -89198 17451 -89182 17468
rect -88398 17468 -87990 17485
rect -87932 17485 -86332 17532
rect -87932 17468 -87524 17485
rect -88398 17451 -88382 17468
rect -89198 17435 -88382 17451
rect -87540 17451 -87524 17468
rect -86740 17468 -86332 17485
rect -86274 17485 -84674 17532
rect -86274 17468 -85866 17485
rect -86740 17451 -86724 17468
rect -87540 17435 -86724 17451
rect -85882 17451 -85866 17468
rect -85082 17468 -84674 17485
rect -84616 17485 -83016 17532
rect -84616 17468 -84208 17485
rect -85082 17451 -85066 17468
rect -85882 17435 -85066 17451
rect -84224 17451 -84208 17468
rect -83424 17468 -83016 17485
rect -82958 17485 -81358 17532
rect -82958 17468 -82550 17485
rect -83424 17451 -83408 17468
rect -84224 17435 -83408 17451
rect -82566 17451 -82550 17468
rect -81766 17468 -81358 17485
rect -81300 17485 -79700 17532
rect -81300 17468 -80892 17485
rect -81766 17451 -81750 17468
rect -82566 17435 -81750 17451
rect -80908 17451 -80892 17468
rect -80108 17468 -79700 17485
rect -79642 17485 -78042 17532
rect -79642 17468 -79234 17485
rect -80108 17451 -80092 17468
rect -80908 17435 -80092 17451
rect -79250 17451 -79234 17468
rect -78450 17468 -78042 17485
rect -77984 17485 -76384 17532
rect -77984 17468 -77576 17485
rect -78450 17451 -78434 17468
rect -79250 17435 -78434 17451
rect -77592 17451 -77576 17468
rect -76792 17468 -76384 17485
rect -76326 17485 -74726 17532
rect -76326 17468 -75918 17485
rect -76792 17451 -76776 17468
rect -77592 17435 -76776 17451
rect -75934 17451 -75918 17468
rect -75134 17468 -74726 17485
rect -74668 17485 -73068 17532
rect -74668 17468 -74260 17485
rect -75134 17451 -75118 17468
rect -75934 17435 -75118 17451
rect -74276 17451 -74260 17468
rect -73476 17468 -73068 17485
rect -73010 17485 -71410 17532
rect -73010 17468 -72602 17485
rect -73476 17451 -73460 17468
rect -74276 17435 -73460 17451
rect -72618 17451 -72602 17468
rect -71818 17468 -71410 17485
rect -71352 17485 -69752 17532
rect -71352 17468 -70944 17485
rect -71818 17451 -71802 17468
rect -72618 17435 -71802 17451
rect -70960 17451 -70944 17468
rect -70160 17468 -69752 17485
rect -69694 17485 -68094 17532
rect -69694 17468 -69286 17485
rect -70160 17451 -70144 17468
rect -70960 17435 -70144 17451
rect -69302 17451 -69286 17468
rect -68502 17468 -68094 17485
rect -68036 17485 -66436 17532
rect -68036 17468 -67628 17485
rect -68502 17451 -68486 17468
rect -69302 17435 -68486 17451
rect -67644 17451 -67628 17468
rect -66844 17468 -66436 17485
rect -66378 17485 -64778 17532
rect -66378 17468 -65970 17485
rect -66844 17451 -66828 17468
rect -67644 17435 -66828 17451
rect -65986 17451 -65970 17468
rect -65186 17468 -64778 17485
rect -64720 17485 -63120 17532
rect -64720 17468 -64312 17485
rect -65186 17451 -65170 17468
rect -65986 17435 -65170 17451
rect -64328 17451 -64312 17468
rect -63528 17468 -63120 17485
rect -63062 17485 -61462 17532
rect -63062 17468 -62654 17485
rect -63528 17451 -63512 17468
rect -64328 17435 -63512 17451
rect -62670 17451 -62654 17468
rect -61870 17468 -61462 17485
rect -61404 17485 -59804 17532
rect -61404 17468 -60996 17485
rect -61870 17451 -61854 17468
rect -62670 17435 -61854 17451
rect -61012 17451 -60996 17468
rect -60212 17468 -59804 17485
rect -59746 17485 -58146 17532
rect -59746 17468 -59338 17485
rect -60212 17451 -60196 17468
rect -61012 17435 -60196 17451
rect -59354 17451 -59338 17468
rect -58554 17468 -58146 17485
rect -58088 17485 -56488 17532
rect -58088 17468 -57680 17485
rect -58554 17451 -58538 17468
rect -59354 17435 -58538 17451
rect -57696 17451 -57680 17468
rect -56896 17468 -56488 17485
rect -56430 17485 -54830 17532
rect -56430 17468 -56022 17485
rect -56896 17451 -56880 17468
rect -57696 17435 -56880 17451
rect -56038 17451 -56022 17468
rect -55238 17468 -54830 17485
rect -54772 17485 -53172 17532
rect -54772 17468 -54364 17485
rect -55238 17451 -55222 17468
rect -56038 17435 -55222 17451
rect -54380 17451 -54364 17468
rect -53580 17468 -53172 17485
rect -53114 17485 -51514 17532
rect -53114 17468 -52706 17485
rect -53580 17451 -53564 17468
rect -54380 17435 -53564 17451
rect -52722 17451 -52706 17468
rect -51922 17468 -51514 17485
rect -51456 17485 -49856 17532
rect -51456 17468 -51048 17485
rect -51922 17451 -51906 17468
rect -52722 17435 -51906 17451
rect -51064 17451 -51048 17468
rect -50264 17468 -49856 17485
rect -49798 17485 -48198 17532
rect -49798 17468 -49390 17485
rect -50264 17451 -50248 17468
rect -51064 17435 -50248 17451
rect -49406 17451 -49390 17468
rect -48606 17468 -48198 17485
rect -48140 17485 -46540 17532
rect -48140 17468 -47732 17485
rect -48606 17451 -48590 17468
rect -49406 17435 -48590 17451
rect -47748 17451 -47732 17468
rect -46948 17468 -46540 17485
rect -46482 17485 -44882 17532
rect -46482 17468 -46074 17485
rect -46948 17451 -46932 17468
rect -47748 17435 -46932 17451
rect -46090 17451 -46074 17468
rect -45290 17468 -44882 17485
rect -44824 17485 -43224 17532
rect -44824 17468 -44416 17485
rect -45290 17451 -45274 17468
rect -46090 17435 -45274 17451
rect -44432 17451 -44416 17468
rect -43632 17468 -43224 17485
rect -43166 17485 -41566 17532
rect -43166 17468 -42758 17485
rect -43632 17451 -43616 17468
rect -44432 17435 -43616 17451
rect -42774 17451 -42758 17468
rect -41974 17468 -41566 17485
rect -41508 17485 -39908 17532
rect -41508 17468 -41100 17485
rect -41974 17451 -41958 17468
rect -42774 17435 -41958 17451
rect -41116 17451 -41100 17468
rect -40316 17468 -39908 17485
rect -39850 17485 -38250 17532
rect -39850 17468 -39442 17485
rect -40316 17451 -40300 17468
rect -41116 17435 -40300 17451
rect -39458 17451 -39442 17468
rect -38658 17468 -38250 17485
rect -38192 17485 -36592 17532
rect -38192 17468 -37784 17485
rect -38658 17451 -38642 17468
rect -39458 17435 -38642 17451
rect -37800 17451 -37784 17468
rect -37000 17468 -36592 17485
rect -36534 17485 -34934 17532
rect -36534 17468 -36126 17485
rect -37000 17451 -36984 17468
rect -37800 17435 -36984 17451
rect -36142 17451 -36126 17468
rect -35342 17468 -34934 17485
rect -34876 17485 -33276 17532
rect -34876 17468 -34468 17485
rect -35342 17451 -35326 17468
rect -36142 17435 -35326 17451
rect -34484 17451 -34468 17468
rect -33684 17468 -33276 17485
rect -33218 17485 -31618 17532
rect -33218 17468 -32810 17485
rect -33684 17451 -33668 17468
rect -34484 17435 -33668 17451
rect -32826 17451 -32810 17468
rect -32026 17468 -31618 17485
rect -31560 17485 -29960 17532
rect -31560 17468 -31152 17485
rect -32026 17451 -32010 17468
rect -32826 17435 -32010 17451
rect -31168 17451 -31152 17468
rect -30368 17468 -29960 17485
rect -29902 17485 -28302 17532
rect -29902 17468 -29494 17485
rect -30368 17451 -30352 17468
rect -31168 17435 -30352 17451
rect -29510 17451 -29494 17468
rect -28710 17468 -28302 17485
rect -28710 17451 -28694 17468
rect -29510 17435 -28694 17451
rect -94170 17267 -93354 17283
rect -94170 17250 -94154 17267
rect -94562 17233 -94154 17250
rect -93370 17250 -93354 17267
rect -92512 17267 -91696 17283
rect -92512 17250 -92496 17267
rect -93370 17233 -92962 17250
rect -94562 17186 -92962 17233
rect -92904 17233 -92496 17250
rect -91712 17250 -91696 17267
rect -90854 17267 -90038 17283
rect -90854 17250 -90838 17267
rect -91712 17233 -91304 17250
rect -92904 17186 -91304 17233
rect -91246 17233 -90838 17250
rect -90054 17250 -90038 17267
rect -89196 17267 -88380 17283
rect -89196 17250 -89180 17267
rect -90054 17233 -89646 17250
rect -91246 17186 -89646 17233
rect -89588 17233 -89180 17250
rect -88396 17250 -88380 17267
rect -87538 17267 -86722 17283
rect -87538 17250 -87522 17267
rect -88396 17233 -87988 17250
rect -89588 17186 -87988 17233
rect -87930 17233 -87522 17250
rect -86738 17250 -86722 17267
rect -85880 17267 -85064 17283
rect -85880 17250 -85864 17267
rect -86738 17233 -86330 17250
rect -87930 17186 -86330 17233
rect -86272 17233 -85864 17250
rect -85080 17250 -85064 17267
rect -84222 17267 -83406 17283
rect -84222 17250 -84206 17267
rect -85080 17233 -84672 17250
rect -86272 17186 -84672 17233
rect -84614 17233 -84206 17250
rect -83422 17250 -83406 17267
rect -82564 17267 -81748 17283
rect -82564 17250 -82548 17267
rect -83422 17233 -83014 17250
rect -84614 17186 -83014 17233
rect -82956 17233 -82548 17250
rect -81764 17250 -81748 17267
rect -80906 17267 -80090 17283
rect -80906 17250 -80890 17267
rect -81764 17233 -81356 17250
rect -82956 17186 -81356 17233
rect -81298 17233 -80890 17250
rect -80106 17250 -80090 17267
rect -79248 17267 -78432 17283
rect -79248 17250 -79232 17267
rect -80106 17233 -79698 17250
rect -81298 17186 -79698 17233
rect -79640 17233 -79232 17250
rect -78448 17250 -78432 17267
rect -77590 17267 -76774 17283
rect -77590 17250 -77574 17267
rect -78448 17233 -78040 17250
rect -79640 17186 -78040 17233
rect -77982 17233 -77574 17250
rect -76790 17250 -76774 17267
rect -75932 17267 -75116 17283
rect -75932 17250 -75916 17267
rect -76790 17233 -76382 17250
rect -77982 17186 -76382 17233
rect -76324 17233 -75916 17250
rect -75132 17250 -75116 17267
rect -74274 17267 -73458 17283
rect -74274 17250 -74258 17267
rect -75132 17233 -74724 17250
rect -76324 17186 -74724 17233
rect -74666 17233 -74258 17250
rect -73474 17250 -73458 17267
rect -72616 17267 -71800 17283
rect -72616 17250 -72600 17267
rect -73474 17233 -73066 17250
rect -74666 17186 -73066 17233
rect -73008 17233 -72600 17250
rect -71816 17250 -71800 17267
rect -70958 17267 -70142 17283
rect -70958 17250 -70942 17267
rect -71816 17233 -71408 17250
rect -73008 17186 -71408 17233
rect -71350 17233 -70942 17250
rect -70158 17250 -70142 17267
rect -69300 17267 -68484 17283
rect -69300 17250 -69284 17267
rect -70158 17233 -69750 17250
rect -71350 17186 -69750 17233
rect -69692 17233 -69284 17250
rect -68500 17250 -68484 17267
rect -67642 17267 -66826 17283
rect -67642 17250 -67626 17267
rect -68500 17233 -68092 17250
rect -69692 17186 -68092 17233
rect -68034 17233 -67626 17250
rect -66842 17250 -66826 17267
rect -65984 17267 -65168 17283
rect -65984 17250 -65968 17267
rect -66842 17233 -66434 17250
rect -68034 17186 -66434 17233
rect -66376 17233 -65968 17250
rect -65184 17250 -65168 17267
rect -64326 17267 -63510 17283
rect -64326 17250 -64310 17267
rect -65184 17233 -64776 17250
rect -66376 17186 -64776 17233
rect -64718 17233 -64310 17250
rect -63526 17250 -63510 17267
rect -62668 17267 -61852 17283
rect -62668 17250 -62652 17267
rect -63526 17233 -63118 17250
rect -64718 17186 -63118 17233
rect -63060 17233 -62652 17250
rect -61868 17250 -61852 17267
rect -61010 17267 -60194 17283
rect -61010 17250 -60994 17267
rect -61868 17233 -61460 17250
rect -63060 17186 -61460 17233
rect -61402 17233 -60994 17250
rect -60210 17250 -60194 17267
rect -59352 17267 -58536 17283
rect -59352 17250 -59336 17267
rect -60210 17233 -59802 17250
rect -61402 17186 -59802 17233
rect -59744 17233 -59336 17250
rect -58552 17250 -58536 17267
rect -57694 17267 -56878 17283
rect -57694 17250 -57678 17267
rect -58552 17233 -58144 17250
rect -59744 17186 -58144 17233
rect -58086 17233 -57678 17250
rect -56894 17250 -56878 17267
rect -56036 17267 -55220 17283
rect -56036 17250 -56020 17267
rect -56894 17233 -56486 17250
rect -58086 17186 -56486 17233
rect -56428 17233 -56020 17250
rect -55236 17250 -55220 17267
rect -54378 17267 -53562 17283
rect -54378 17250 -54362 17267
rect -55236 17233 -54828 17250
rect -56428 17186 -54828 17233
rect -54770 17233 -54362 17250
rect -53578 17250 -53562 17267
rect -52720 17267 -51904 17283
rect -52720 17250 -52704 17267
rect -53578 17233 -53170 17250
rect -54770 17186 -53170 17233
rect -53112 17233 -52704 17250
rect -51920 17250 -51904 17267
rect -51062 17267 -50246 17283
rect -51062 17250 -51046 17267
rect -51920 17233 -51512 17250
rect -53112 17186 -51512 17233
rect -51454 17233 -51046 17250
rect -50262 17250 -50246 17267
rect -49404 17267 -48588 17283
rect -49404 17250 -49388 17267
rect -50262 17233 -49854 17250
rect -51454 17186 -49854 17233
rect -49796 17233 -49388 17250
rect -48604 17250 -48588 17267
rect -47746 17267 -46930 17283
rect -47746 17250 -47730 17267
rect -48604 17233 -48196 17250
rect -49796 17186 -48196 17233
rect -48138 17233 -47730 17250
rect -46946 17250 -46930 17267
rect -46088 17267 -45272 17283
rect -46088 17250 -46072 17267
rect -46946 17233 -46538 17250
rect -48138 17186 -46538 17233
rect -46480 17233 -46072 17250
rect -45288 17250 -45272 17267
rect -44430 17267 -43614 17283
rect -44430 17250 -44414 17267
rect -45288 17233 -44880 17250
rect -46480 17186 -44880 17233
rect -44822 17233 -44414 17250
rect -43630 17250 -43614 17267
rect -42772 17267 -41956 17283
rect -42772 17250 -42756 17267
rect -43630 17233 -43222 17250
rect -44822 17186 -43222 17233
rect -43164 17233 -42756 17250
rect -41972 17250 -41956 17267
rect -41114 17267 -40298 17283
rect -41114 17250 -41098 17267
rect -41972 17233 -41564 17250
rect -43164 17186 -41564 17233
rect -41506 17233 -41098 17250
rect -40314 17250 -40298 17267
rect -39456 17267 -38640 17283
rect -39456 17250 -39440 17267
rect -40314 17233 -39906 17250
rect -41506 17186 -39906 17233
rect -39848 17233 -39440 17250
rect -38656 17250 -38640 17267
rect -37798 17267 -36982 17283
rect -37798 17250 -37782 17267
rect -38656 17233 -38248 17250
rect -39848 17186 -38248 17233
rect -38190 17233 -37782 17250
rect -36998 17250 -36982 17267
rect -36140 17267 -35324 17283
rect -36140 17250 -36124 17267
rect -36998 17233 -36590 17250
rect -38190 17186 -36590 17233
rect -36532 17233 -36124 17250
rect -35340 17250 -35324 17267
rect -34482 17267 -33666 17283
rect -34482 17250 -34466 17267
rect -35340 17233 -34932 17250
rect -36532 17186 -34932 17233
rect -34874 17233 -34466 17250
rect -33682 17250 -33666 17267
rect -32824 17267 -32008 17283
rect -32824 17250 -32808 17267
rect -33682 17233 -33274 17250
rect -34874 17186 -33274 17233
rect -33216 17233 -32808 17250
rect -32024 17250 -32008 17267
rect -31166 17267 -30350 17283
rect -31166 17250 -31150 17267
rect -32024 17233 -31616 17250
rect -33216 17186 -31616 17233
rect -31558 17233 -31150 17250
rect -30366 17250 -30350 17267
rect -29508 17267 -28692 17283
rect -29508 17250 -29492 17267
rect -30366 17233 -29958 17250
rect -31558 17186 -29958 17233
rect -29900 17233 -29492 17250
rect -28708 17250 -28692 17267
rect -28708 17233 -28300 17250
rect -29900 17186 -28300 17233
rect -94562 15739 -92962 15786
rect -94562 15722 -94154 15739
rect -94170 15705 -94154 15722
rect -93370 15722 -92962 15739
rect -92904 15739 -91304 15786
rect -92904 15722 -92496 15739
rect -93370 15705 -93354 15722
rect -94170 15689 -93354 15705
rect -92512 15705 -92496 15722
rect -91712 15722 -91304 15739
rect -91246 15739 -89646 15786
rect -91246 15722 -90838 15739
rect -91712 15705 -91696 15722
rect -92512 15689 -91696 15705
rect -90854 15705 -90838 15722
rect -90054 15722 -89646 15739
rect -89588 15739 -87988 15786
rect -89588 15722 -89180 15739
rect -90054 15705 -90038 15722
rect -90854 15689 -90038 15705
rect -89196 15705 -89180 15722
rect -88396 15722 -87988 15739
rect -87930 15739 -86330 15786
rect -87930 15722 -87522 15739
rect -88396 15705 -88380 15722
rect -89196 15689 -88380 15705
rect -87538 15705 -87522 15722
rect -86738 15722 -86330 15739
rect -86272 15739 -84672 15786
rect -86272 15722 -85864 15739
rect -86738 15705 -86722 15722
rect -87538 15689 -86722 15705
rect -85880 15705 -85864 15722
rect -85080 15722 -84672 15739
rect -84614 15739 -83014 15786
rect -84614 15722 -84206 15739
rect -85080 15705 -85064 15722
rect -85880 15689 -85064 15705
rect -84222 15705 -84206 15722
rect -83422 15722 -83014 15739
rect -82956 15739 -81356 15786
rect -82956 15722 -82548 15739
rect -83422 15705 -83406 15722
rect -84222 15689 -83406 15705
rect -82564 15705 -82548 15722
rect -81764 15722 -81356 15739
rect -81298 15739 -79698 15786
rect -81298 15722 -80890 15739
rect -81764 15705 -81748 15722
rect -82564 15689 -81748 15705
rect -80906 15705 -80890 15722
rect -80106 15722 -79698 15739
rect -79640 15739 -78040 15786
rect -79640 15722 -79232 15739
rect -80106 15705 -80090 15722
rect -80906 15689 -80090 15705
rect -79248 15705 -79232 15722
rect -78448 15722 -78040 15739
rect -77982 15739 -76382 15786
rect -77982 15722 -77574 15739
rect -78448 15705 -78432 15722
rect -79248 15689 -78432 15705
rect -77590 15705 -77574 15722
rect -76790 15722 -76382 15739
rect -76324 15739 -74724 15786
rect -76324 15722 -75916 15739
rect -76790 15705 -76774 15722
rect -77590 15689 -76774 15705
rect -75932 15705 -75916 15722
rect -75132 15722 -74724 15739
rect -74666 15739 -73066 15786
rect -74666 15722 -74258 15739
rect -75132 15705 -75116 15722
rect -75932 15689 -75116 15705
rect -74274 15705 -74258 15722
rect -73474 15722 -73066 15739
rect -73008 15739 -71408 15786
rect -73008 15722 -72600 15739
rect -73474 15705 -73458 15722
rect -74274 15689 -73458 15705
rect -72616 15705 -72600 15722
rect -71816 15722 -71408 15739
rect -71350 15739 -69750 15786
rect -71350 15722 -70942 15739
rect -71816 15705 -71800 15722
rect -72616 15689 -71800 15705
rect -70958 15705 -70942 15722
rect -70158 15722 -69750 15739
rect -69692 15739 -68092 15786
rect -69692 15722 -69284 15739
rect -70158 15705 -70142 15722
rect -70958 15689 -70142 15705
rect -69300 15705 -69284 15722
rect -68500 15722 -68092 15739
rect -68034 15739 -66434 15786
rect -68034 15722 -67626 15739
rect -68500 15705 -68484 15722
rect -69300 15689 -68484 15705
rect -67642 15705 -67626 15722
rect -66842 15722 -66434 15739
rect -66376 15739 -64776 15786
rect -66376 15722 -65968 15739
rect -66842 15705 -66826 15722
rect -67642 15689 -66826 15705
rect -65984 15705 -65968 15722
rect -65184 15722 -64776 15739
rect -64718 15739 -63118 15786
rect -64718 15722 -64310 15739
rect -65184 15705 -65168 15722
rect -65984 15689 -65168 15705
rect -64326 15705 -64310 15722
rect -63526 15722 -63118 15739
rect -63060 15739 -61460 15786
rect -63060 15722 -62652 15739
rect -63526 15705 -63510 15722
rect -64326 15689 -63510 15705
rect -62668 15705 -62652 15722
rect -61868 15722 -61460 15739
rect -61402 15739 -59802 15786
rect -61402 15722 -60994 15739
rect -61868 15705 -61852 15722
rect -62668 15689 -61852 15705
rect -61010 15705 -60994 15722
rect -60210 15722 -59802 15739
rect -59744 15739 -58144 15786
rect -59744 15722 -59336 15739
rect -60210 15705 -60194 15722
rect -61010 15689 -60194 15705
rect -59352 15705 -59336 15722
rect -58552 15722 -58144 15739
rect -58086 15739 -56486 15786
rect -58086 15722 -57678 15739
rect -58552 15705 -58536 15722
rect -59352 15689 -58536 15705
rect -57694 15705 -57678 15722
rect -56894 15722 -56486 15739
rect -56428 15739 -54828 15786
rect -56428 15722 -56020 15739
rect -56894 15705 -56878 15722
rect -57694 15689 -56878 15705
rect -56036 15705 -56020 15722
rect -55236 15722 -54828 15739
rect -54770 15739 -53170 15786
rect -54770 15722 -54362 15739
rect -55236 15705 -55220 15722
rect -56036 15689 -55220 15705
rect -54378 15705 -54362 15722
rect -53578 15722 -53170 15739
rect -53112 15739 -51512 15786
rect -53112 15722 -52704 15739
rect -53578 15705 -53562 15722
rect -54378 15689 -53562 15705
rect -52720 15705 -52704 15722
rect -51920 15722 -51512 15739
rect -51454 15739 -49854 15786
rect -51454 15722 -51046 15739
rect -51920 15705 -51904 15722
rect -52720 15689 -51904 15705
rect -51062 15705 -51046 15722
rect -50262 15722 -49854 15739
rect -49796 15739 -48196 15786
rect -49796 15722 -49388 15739
rect -50262 15705 -50246 15722
rect -51062 15689 -50246 15705
rect -49404 15705 -49388 15722
rect -48604 15722 -48196 15739
rect -48138 15739 -46538 15786
rect -48138 15722 -47730 15739
rect -48604 15705 -48588 15722
rect -49404 15689 -48588 15705
rect -47746 15705 -47730 15722
rect -46946 15722 -46538 15739
rect -46480 15739 -44880 15786
rect -46480 15722 -46072 15739
rect -46946 15705 -46930 15722
rect -47746 15689 -46930 15705
rect -46088 15705 -46072 15722
rect -45288 15722 -44880 15739
rect -44822 15739 -43222 15786
rect -44822 15722 -44414 15739
rect -45288 15705 -45272 15722
rect -46088 15689 -45272 15705
rect -44430 15705 -44414 15722
rect -43630 15722 -43222 15739
rect -43164 15739 -41564 15786
rect -43164 15722 -42756 15739
rect -43630 15705 -43614 15722
rect -44430 15689 -43614 15705
rect -42772 15705 -42756 15722
rect -41972 15722 -41564 15739
rect -41506 15739 -39906 15786
rect -41506 15722 -41098 15739
rect -41972 15705 -41956 15722
rect -42772 15689 -41956 15705
rect -41114 15705 -41098 15722
rect -40314 15722 -39906 15739
rect -39848 15739 -38248 15786
rect -39848 15722 -39440 15739
rect -40314 15705 -40298 15722
rect -41114 15689 -40298 15705
rect -39456 15705 -39440 15722
rect -38656 15722 -38248 15739
rect -38190 15739 -36590 15786
rect -38190 15722 -37782 15739
rect -38656 15705 -38640 15722
rect -39456 15689 -38640 15705
rect -37798 15705 -37782 15722
rect -36998 15722 -36590 15739
rect -36532 15739 -34932 15786
rect -36532 15722 -36124 15739
rect -36998 15705 -36982 15722
rect -37798 15689 -36982 15705
rect -36140 15705 -36124 15722
rect -35340 15722 -34932 15739
rect -34874 15739 -33274 15786
rect -34874 15722 -34466 15739
rect -35340 15705 -35324 15722
rect -36140 15689 -35324 15705
rect -34482 15705 -34466 15722
rect -33682 15722 -33274 15739
rect -33216 15739 -31616 15786
rect -33216 15722 -32808 15739
rect -33682 15705 -33666 15722
rect -34482 15689 -33666 15705
rect -32824 15705 -32808 15722
rect -32024 15722 -31616 15739
rect -31558 15739 -29958 15786
rect -31558 15722 -31150 15739
rect -32024 15705 -32008 15722
rect -32824 15689 -32008 15705
rect -31166 15705 -31150 15722
rect -30366 15722 -29958 15739
rect -29900 15739 -28300 15786
rect -29900 15722 -29492 15739
rect -30366 15705 -30350 15722
rect -31166 15689 -30350 15705
rect -29508 15705 -29492 15722
rect -28708 15722 -28300 15739
rect -28708 15705 -28692 15722
rect -29508 15689 -28692 15705
rect -94170 15631 -93354 15647
rect -94170 15614 -94154 15631
rect -94562 15597 -94154 15614
rect -93370 15614 -93354 15631
rect -92512 15631 -91696 15647
rect -92512 15614 -92496 15631
rect -93370 15597 -92962 15614
rect -94562 15550 -92962 15597
rect -92904 15597 -92496 15614
rect -91712 15614 -91696 15631
rect -90854 15631 -90038 15647
rect -90854 15614 -90838 15631
rect -91712 15597 -91304 15614
rect -92904 15550 -91304 15597
rect -91246 15597 -90838 15614
rect -90054 15614 -90038 15631
rect -89196 15631 -88380 15647
rect -89196 15614 -89180 15631
rect -90054 15597 -89646 15614
rect -91246 15550 -89646 15597
rect -89588 15597 -89180 15614
rect -88396 15614 -88380 15631
rect -87538 15631 -86722 15647
rect -87538 15614 -87522 15631
rect -88396 15597 -87988 15614
rect -89588 15550 -87988 15597
rect -87930 15597 -87522 15614
rect -86738 15614 -86722 15631
rect -85880 15631 -85064 15647
rect -85880 15614 -85864 15631
rect -86738 15597 -86330 15614
rect -87930 15550 -86330 15597
rect -86272 15597 -85864 15614
rect -85080 15614 -85064 15631
rect -84222 15631 -83406 15647
rect -84222 15614 -84206 15631
rect -85080 15597 -84672 15614
rect -86272 15550 -84672 15597
rect -84614 15597 -84206 15614
rect -83422 15614 -83406 15631
rect -82564 15631 -81748 15647
rect -82564 15614 -82548 15631
rect -83422 15597 -83014 15614
rect -84614 15550 -83014 15597
rect -82956 15597 -82548 15614
rect -81764 15614 -81748 15631
rect -80906 15631 -80090 15647
rect -80906 15614 -80890 15631
rect -81764 15597 -81356 15614
rect -82956 15550 -81356 15597
rect -81298 15597 -80890 15614
rect -80106 15614 -80090 15631
rect -79248 15631 -78432 15647
rect -79248 15614 -79232 15631
rect -80106 15597 -79698 15614
rect -81298 15550 -79698 15597
rect -79640 15597 -79232 15614
rect -78448 15614 -78432 15631
rect -77590 15631 -76774 15647
rect -77590 15614 -77574 15631
rect -78448 15597 -78040 15614
rect -79640 15550 -78040 15597
rect -77982 15597 -77574 15614
rect -76790 15614 -76774 15631
rect -75932 15631 -75116 15647
rect -75932 15614 -75916 15631
rect -76790 15597 -76382 15614
rect -77982 15550 -76382 15597
rect -76324 15597 -75916 15614
rect -75132 15614 -75116 15631
rect -74274 15631 -73458 15647
rect -74274 15614 -74258 15631
rect -75132 15597 -74724 15614
rect -76324 15550 -74724 15597
rect -74666 15597 -74258 15614
rect -73474 15614 -73458 15631
rect -72616 15631 -71800 15647
rect -72616 15614 -72600 15631
rect -73474 15597 -73066 15614
rect -74666 15550 -73066 15597
rect -73008 15597 -72600 15614
rect -71816 15614 -71800 15631
rect -70958 15631 -70142 15647
rect -70958 15614 -70942 15631
rect -71816 15597 -71408 15614
rect -73008 15550 -71408 15597
rect -71350 15597 -70942 15614
rect -70158 15614 -70142 15631
rect -69300 15631 -68484 15647
rect -69300 15614 -69284 15631
rect -70158 15597 -69750 15614
rect -71350 15550 -69750 15597
rect -69692 15597 -69284 15614
rect -68500 15614 -68484 15631
rect -67642 15631 -66826 15647
rect -67642 15614 -67626 15631
rect -68500 15597 -68092 15614
rect -69692 15550 -68092 15597
rect -68034 15597 -67626 15614
rect -66842 15614 -66826 15631
rect -65984 15631 -65168 15647
rect -65984 15614 -65968 15631
rect -66842 15597 -66434 15614
rect -68034 15550 -66434 15597
rect -66376 15597 -65968 15614
rect -65184 15614 -65168 15631
rect -64326 15631 -63510 15647
rect -64326 15614 -64310 15631
rect -65184 15597 -64776 15614
rect -66376 15550 -64776 15597
rect -64718 15597 -64310 15614
rect -63526 15614 -63510 15631
rect -62668 15631 -61852 15647
rect -62668 15614 -62652 15631
rect -63526 15597 -63118 15614
rect -64718 15550 -63118 15597
rect -63060 15597 -62652 15614
rect -61868 15614 -61852 15631
rect -61010 15631 -60194 15647
rect -61010 15614 -60994 15631
rect -61868 15597 -61460 15614
rect -63060 15550 -61460 15597
rect -61402 15597 -60994 15614
rect -60210 15614 -60194 15631
rect -59352 15631 -58536 15647
rect -59352 15614 -59336 15631
rect -60210 15597 -59802 15614
rect -61402 15550 -59802 15597
rect -59744 15597 -59336 15614
rect -58552 15614 -58536 15631
rect -57694 15631 -56878 15647
rect -57694 15614 -57678 15631
rect -58552 15597 -58144 15614
rect -59744 15550 -58144 15597
rect -58086 15597 -57678 15614
rect -56894 15614 -56878 15631
rect -56036 15631 -55220 15647
rect -56036 15614 -56020 15631
rect -56894 15597 -56486 15614
rect -58086 15550 -56486 15597
rect -56428 15597 -56020 15614
rect -55236 15614 -55220 15631
rect -54378 15631 -53562 15647
rect -54378 15614 -54362 15631
rect -55236 15597 -54828 15614
rect -56428 15550 -54828 15597
rect -54770 15597 -54362 15614
rect -53578 15614 -53562 15631
rect -52720 15631 -51904 15647
rect -52720 15614 -52704 15631
rect -53578 15597 -53170 15614
rect -54770 15550 -53170 15597
rect -53112 15597 -52704 15614
rect -51920 15614 -51904 15631
rect -51062 15631 -50246 15647
rect -51062 15614 -51046 15631
rect -51920 15597 -51512 15614
rect -53112 15550 -51512 15597
rect -51454 15597 -51046 15614
rect -50262 15614 -50246 15631
rect -49404 15631 -48588 15647
rect -49404 15614 -49388 15631
rect -50262 15597 -49854 15614
rect -51454 15550 -49854 15597
rect -49796 15597 -49388 15614
rect -48604 15614 -48588 15631
rect -47746 15631 -46930 15647
rect -47746 15614 -47730 15631
rect -48604 15597 -48196 15614
rect -49796 15550 -48196 15597
rect -48138 15597 -47730 15614
rect -46946 15614 -46930 15631
rect -46088 15631 -45272 15647
rect -46088 15614 -46072 15631
rect -46946 15597 -46538 15614
rect -48138 15550 -46538 15597
rect -46480 15597 -46072 15614
rect -45288 15614 -45272 15631
rect -44430 15631 -43614 15647
rect -44430 15614 -44414 15631
rect -45288 15597 -44880 15614
rect -46480 15550 -44880 15597
rect -44822 15597 -44414 15614
rect -43630 15614 -43614 15631
rect -42772 15631 -41956 15647
rect -42772 15614 -42756 15631
rect -43630 15597 -43222 15614
rect -44822 15550 -43222 15597
rect -43164 15597 -42756 15614
rect -41972 15614 -41956 15631
rect -41114 15631 -40298 15647
rect -41114 15614 -41098 15631
rect -41972 15597 -41564 15614
rect -43164 15550 -41564 15597
rect -41506 15597 -41098 15614
rect -40314 15614 -40298 15631
rect -39456 15631 -38640 15647
rect -39456 15614 -39440 15631
rect -40314 15597 -39906 15614
rect -41506 15550 -39906 15597
rect -39848 15597 -39440 15614
rect -38656 15614 -38640 15631
rect -37798 15631 -36982 15647
rect -37798 15614 -37782 15631
rect -38656 15597 -38248 15614
rect -39848 15550 -38248 15597
rect -38190 15597 -37782 15614
rect -36998 15614 -36982 15631
rect -36140 15631 -35324 15647
rect -36140 15614 -36124 15631
rect -36998 15597 -36590 15614
rect -38190 15550 -36590 15597
rect -36532 15597 -36124 15614
rect -35340 15614 -35324 15631
rect -34482 15631 -33666 15647
rect -34482 15614 -34466 15631
rect -35340 15597 -34932 15614
rect -36532 15550 -34932 15597
rect -34874 15597 -34466 15614
rect -33682 15614 -33666 15631
rect -32824 15631 -32008 15647
rect -32824 15614 -32808 15631
rect -33682 15597 -33274 15614
rect -34874 15550 -33274 15597
rect -33216 15597 -32808 15614
rect -32024 15614 -32008 15631
rect -31166 15631 -30350 15647
rect -31166 15614 -31150 15631
rect -32024 15597 -31616 15614
rect -33216 15550 -31616 15597
rect -31558 15597 -31150 15614
rect -30366 15614 -30350 15631
rect -29508 15631 -28692 15647
rect -29508 15614 -29492 15631
rect -30366 15597 -29958 15614
rect -31558 15550 -29958 15597
rect -29900 15597 -29492 15614
rect -28708 15614 -28692 15631
rect -28708 15597 -28300 15614
rect -29900 15550 -28300 15597
rect -94562 14103 -92962 14150
rect -94562 14086 -94154 14103
rect -94170 14069 -94154 14086
rect -93370 14086 -92962 14103
rect -92904 14103 -91304 14150
rect -92904 14086 -92496 14103
rect -93370 14069 -93354 14086
rect -94170 14053 -93354 14069
rect -92512 14069 -92496 14086
rect -91712 14086 -91304 14103
rect -91246 14103 -89646 14150
rect -91246 14086 -90838 14103
rect -91712 14069 -91696 14086
rect -92512 14053 -91696 14069
rect -90854 14069 -90838 14086
rect -90054 14086 -89646 14103
rect -89588 14103 -87988 14150
rect -89588 14086 -89180 14103
rect -90054 14069 -90038 14086
rect -90854 14053 -90038 14069
rect -89196 14069 -89180 14086
rect -88396 14086 -87988 14103
rect -87930 14103 -86330 14150
rect -87930 14086 -87522 14103
rect -88396 14069 -88380 14086
rect -89196 14053 -88380 14069
rect -87538 14069 -87522 14086
rect -86738 14086 -86330 14103
rect -86272 14103 -84672 14150
rect -86272 14086 -85864 14103
rect -86738 14069 -86722 14086
rect -87538 14053 -86722 14069
rect -85880 14069 -85864 14086
rect -85080 14086 -84672 14103
rect -84614 14103 -83014 14150
rect -84614 14086 -84206 14103
rect -85080 14069 -85064 14086
rect -85880 14053 -85064 14069
rect -84222 14069 -84206 14086
rect -83422 14086 -83014 14103
rect -82956 14103 -81356 14150
rect -82956 14086 -82548 14103
rect -83422 14069 -83406 14086
rect -84222 14053 -83406 14069
rect -82564 14069 -82548 14086
rect -81764 14086 -81356 14103
rect -81298 14103 -79698 14150
rect -81298 14086 -80890 14103
rect -81764 14069 -81748 14086
rect -82564 14053 -81748 14069
rect -80906 14069 -80890 14086
rect -80106 14086 -79698 14103
rect -79640 14103 -78040 14150
rect -79640 14086 -79232 14103
rect -80106 14069 -80090 14086
rect -80906 14053 -80090 14069
rect -79248 14069 -79232 14086
rect -78448 14086 -78040 14103
rect -77982 14103 -76382 14150
rect -77982 14086 -77574 14103
rect -78448 14069 -78432 14086
rect -79248 14053 -78432 14069
rect -77590 14069 -77574 14086
rect -76790 14086 -76382 14103
rect -76324 14103 -74724 14150
rect -76324 14086 -75916 14103
rect -76790 14069 -76774 14086
rect -77590 14053 -76774 14069
rect -75932 14069 -75916 14086
rect -75132 14086 -74724 14103
rect -74666 14103 -73066 14150
rect -74666 14086 -74258 14103
rect -75132 14069 -75116 14086
rect -75932 14053 -75116 14069
rect -74274 14069 -74258 14086
rect -73474 14086 -73066 14103
rect -73008 14103 -71408 14150
rect -73008 14086 -72600 14103
rect -73474 14069 -73458 14086
rect -74274 14053 -73458 14069
rect -72616 14069 -72600 14086
rect -71816 14086 -71408 14103
rect -71350 14103 -69750 14150
rect -71350 14086 -70942 14103
rect -71816 14069 -71800 14086
rect -72616 14053 -71800 14069
rect -70958 14069 -70942 14086
rect -70158 14086 -69750 14103
rect -69692 14103 -68092 14150
rect -69692 14086 -69284 14103
rect -70158 14069 -70142 14086
rect -70958 14053 -70142 14069
rect -69300 14069 -69284 14086
rect -68500 14086 -68092 14103
rect -68034 14103 -66434 14150
rect -68034 14086 -67626 14103
rect -68500 14069 -68484 14086
rect -69300 14053 -68484 14069
rect -67642 14069 -67626 14086
rect -66842 14086 -66434 14103
rect -66376 14103 -64776 14150
rect -66376 14086 -65968 14103
rect -66842 14069 -66826 14086
rect -67642 14053 -66826 14069
rect -65984 14069 -65968 14086
rect -65184 14086 -64776 14103
rect -64718 14103 -63118 14150
rect -64718 14086 -64310 14103
rect -65184 14069 -65168 14086
rect -65984 14053 -65168 14069
rect -64326 14069 -64310 14086
rect -63526 14086 -63118 14103
rect -63060 14103 -61460 14150
rect -63060 14086 -62652 14103
rect -63526 14069 -63510 14086
rect -64326 14053 -63510 14069
rect -62668 14069 -62652 14086
rect -61868 14086 -61460 14103
rect -61402 14103 -59802 14150
rect -61402 14086 -60994 14103
rect -61868 14069 -61852 14086
rect -62668 14053 -61852 14069
rect -61010 14069 -60994 14086
rect -60210 14086 -59802 14103
rect -59744 14103 -58144 14150
rect -59744 14086 -59336 14103
rect -60210 14069 -60194 14086
rect -61010 14053 -60194 14069
rect -59352 14069 -59336 14086
rect -58552 14086 -58144 14103
rect -58086 14103 -56486 14150
rect -58086 14086 -57678 14103
rect -58552 14069 -58536 14086
rect -59352 14053 -58536 14069
rect -57694 14069 -57678 14086
rect -56894 14086 -56486 14103
rect -56428 14103 -54828 14150
rect -56428 14086 -56020 14103
rect -56894 14069 -56878 14086
rect -57694 14053 -56878 14069
rect -56036 14069 -56020 14086
rect -55236 14086 -54828 14103
rect -54770 14103 -53170 14150
rect -54770 14086 -54362 14103
rect -55236 14069 -55220 14086
rect -56036 14053 -55220 14069
rect -54378 14069 -54362 14086
rect -53578 14086 -53170 14103
rect -53112 14103 -51512 14150
rect -53112 14086 -52704 14103
rect -53578 14069 -53562 14086
rect -54378 14053 -53562 14069
rect -52720 14069 -52704 14086
rect -51920 14086 -51512 14103
rect -51454 14103 -49854 14150
rect -51454 14086 -51046 14103
rect -51920 14069 -51904 14086
rect -52720 14053 -51904 14069
rect -51062 14069 -51046 14086
rect -50262 14086 -49854 14103
rect -49796 14103 -48196 14150
rect -49796 14086 -49388 14103
rect -50262 14069 -50246 14086
rect -51062 14053 -50246 14069
rect -49404 14069 -49388 14086
rect -48604 14086 -48196 14103
rect -48138 14103 -46538 14150
rect -48138 14086 -47730 14103
rect -48604 14069 -48588 14086
rect -49404 14053 -48588 14069
rect -47746 14069 -47730 14086
rect -46946 14086 -46538 14103
rect -46480 14103 -44880 14150
rect -46480 14086 -46072 14103
rect -46946 14069 -46930 14086
rect -47746 14053 -46930 14069
rect -46088 14069 -46072 14086
rect -45288 14086 -44880 14103
rect -44822 14103 -43222 14150
rect -44822 14086 -44414 14103
rect -45288 14069 -45272 14086
rect -46088 14053 -45272 14069
rect -44430 14069 -44414 14086
rect -43630 14086 -43222 14103
rect -43164 14103 -41564 14150
rect -43164 14086 -42756 14103
rect -43630 14069 -43614 14086
rect -44430 14053 -43614 14069
rect -42772 14069 -42756 14086
rect -41972 14086 -41564 14103
rect -41506 14103 -39906 14150
rect -41506 14086 -41098 14103
rect -41972 14069 -41956 14086
rect -42772 14053 -41956 14069
rect -41114 14069 -41098 14086
rect -40314 14086 -39906 14103
rect -39848 14103 -38248 14150
rect -39848 14086 -39440 14103
rect -40314 14069 -40298 14086
rect -41114 14053 -40298 14069
rect -39456 14069 -39440 14086
rect -38656 14086 -38248 14103
rect -38190 14103 -36590 14150
rect -38190 14086 -37782 14103
rect -38656 14069 -38640 14086
rect -39456 14053 -38640 14069
rect -37798 14069 -37782 14086
rect -36998 14086 -36590 14103
rect -36532 14103 -34932 14150
rect -36532 14086 -36124 14103
rect -36998 14069 -36982 14086
rect -37798 14053 -36982 14069
rect -36140 14069 -36124 14086
rect -35340 14086 -34932 14103
rect -34874 14103 -33274 14150
rect -34874 14086 -34466 14103
rect -35340 14069 -35324 14086
rect -36140 14053 -35324 14069
rect -34482 14069 -34466 14086
rect -33682 14086 -33274 14103
rect -33216 14103 -31616 14150
rect -33216 14086 -32808 14103
rect -33682 14069 -33666 14086
rect -34482 14053 -33666 14069
rect -32824 14069 -32808 14086
rect -32024 14086 -31616 14103
rect -31558 14103 -29958 14150
rect -31558 14086 -31150 14103
rect -32024 14069 -32008 14086
rect -32824 14053 -32008 14069
rect -31166 14069 -31150 14086
rect -30366 14086 -29958 14103
rect -29900 14103 -28300 14150
rect -29900 14086 -29492 14103
rect -30366 14069 -30350 14086
rect -31166 14053 -30350 14069
rect -29508 14069 -29492 14086
rect -28708 14086 -28300 14103
rect -28708 14069 -28692 14086
rect -29508 14053 -28692 14069
rect -94170 13995 -93354 14011
rect -94170 13978 -94154 13995
rect -94562 13961 -94154 13978
rect -93370 13978 -93354 13995
rect -92512 13995 -91696 14011
rect -92512 13978 -92496 13995
rect -93370 13961 -92962 13978
rect -94562 13914 -92962 13961
rect -92904 13961 -92496 13978
rect -91712 13978 -91696 13995
rect -90854 13995 -90038 14011
rect -90854 13978 -90838 13995
rect -91712 13961 -91304 13978
rect -92904 13914 -91304 13961
rect -91246 13961 -90838 13978
rect -90054 13978 -90038 13995
rect -89196 13995 -88380 14011
rect -89196 13978 -89180 13995
rect -90054 13961 -89646 13978
rect -91246 13914 -89646 13961
rect -89588 13961 -89180 13978
rect -88396 13978 -88380 13995
rect -87538 13995 -86722 14011
rect -87538 13978 -87522 13995
rect -88396 13961 -87988 13978
rect -89588 13914 -87988 13961
rect -87930 13961 -87522 13978
rect -86738 13978 -86722 13995
rect -85880 13995 -85064 14011
rect -85880 13978 -85864 13995
rect -86738 13961 -86330 13978
rect -87930 13914 -86330 13961
rect -86272 13961 -85864 13978
rect -85080 13978 -85064 13995
rect -84222 13995 -83406 14011
rect -84222 13978 -84206 13995
rect -85080 13961 -84672 13978
rect -86272 13914 -84672 13961
rect -84614 13961 -84206 13978
rect -83422 13978 -83406 13995
rect -82564 13995 -81748 14011
rect -82564 13978 -82548 13995
rect -83422 13961 -83014 13978
rect -84614 13914 -83014 13961
rect -82956 13961 -82548 13978
rect -81764 13978 -81748 13995
rect -80906 13995 -80090 14011
rect -80906 13978 -80890 13995
rect -81764 13961 -81356 13978
rect -82956 13914 -81356 13961
rect -81298 13961 -80890 13978
rect -80106 13978 -80090 13995
rect -79248 13995 -78432 14011
rect -79248 13978 -79232 13995
rect -80106 13961 -79698 13978
rect -81298 13914 -79698 13961
rect -79640 13961 -79232 13978
rect -78448 13978 -78432 13995
rect -77590 13995 -76774 14011
rect -77590 13978 -77574 13995
rect -78448 13961 -78040 13978
rect -79640 13914 -78040 13961
rect -77982 13961 -77574 13978
rect -76790 13978 -76774 13995
rect -75932 13995 -75116 14011
rect -75932 13978 -75916 13995
rect -76790 13961 -76382 13978
rect -77982 13914 -76382 13961
rect -76324 13961 -75916 13978
rect -75132 13978 -75116 13995
rect -74274 13995 -73458 14011
rect -74274 13978 -74258 13995
rect -75132 13961 -74724 13978
rect -76324 13914 -74724 13961
rect -74666 13961 -74258 13978
rect -73474 13978 -73458 13995
rect -72616 13995 -71800 14011
rect -72616 13978 -72600 13995
rect -73474 13961 -73066 13978
rect -74666 13914 -73066 13961
rect -73008 13961 -72600 13978
rect -71816 13978 -71800 13995
rect -70958 13995 -70142 14011
rect -70958 13978 -70942 13995
rect -71816 13961 -71408 13978
rect -73008 13914 -71408 13961
rect -71350 13961 -70942 13978
rect -70158 13978 -70142 13995
rect -69300 13995 -68484 14011
rect -69300 13978 -69284 13995
rect -70158 13961 -69750 13978
rect -71350 13914 -69750 13961
rect -69692 13961 -69284 13978
rect -68500 13978 -68484 13995
rect -67642 13995 -66826 14011
rect -67642 13978 -67626 13995
rect -68500 13961 -68092 13978
rect -69692 13914 -68092 13961
rect -68034 13961 -67626 13978
rect -66842 13978 -66826 13995
rect -65984 13995 -65168 14011
rect -65984 13978 -65968 13995
rect -66842 13961 -66434 13978
rect -68034 13914 -66434 13961
rect -66376 13961 -65968 13978
rect -65184 13978 -65168 13995
rect -64326 13995 -63510 14011
rect -64326 13978 -64310 13995
rect -65184 13961 -64776 13978
rect -66376 13914 -64776 13961
rect -64718 13961 -64310 13978
rect -63526 13978 -63510 13995
rect -62668 13995 -61852 14011
rect -62668 13978 -62652 13995
rect -63526 13961 -63118 13978
rect -64718 13914 -63118 13961
rect -63060 13961 -62652 13978
rect -61868 13978 -61852 13995
rect -61010 13995 -60194 14011
rect -61010 13978 -60994 13995
rect -61868 13961 -61460 13978
rect -63060 13914 -61460 13961
rect -61402 13961 -60994 13978
rect -60210 13978 -60194 13995
rect -59352 13995 -58536 14011
rect -59352 13978 -59336 13995
rect -60210 13961 -59802 13978
rect -61402 13914 -59802 13961
rect -59744 13961 -59336 13978
rect -58552 13978 -58536 13995
rect -57694 13995 -56878 14011
rect -57694 13978 -57678 13995
rect -58552 13961 -58144 13978
rect -59744 13914 -58144 13961
rect -58086 13961 -57678 13978
rect -56894 13978 -56878 13995
rect -56036 13995 -55220 14011
rect -56036 13978 -56020 13995
rect -56894 13961 -56486 13978
rect -58086 13914 -56486 13961
rect -56428 13961 -56020 13978
rect -55236 13978 -55220 13995
rect -54378 13995 -53562 14011
rect -54378 13978 -54362 13995
rect -55236 13961 -54828 13978
rect -56428 13914 -54828 13961
rect -54770 13961 -54362 13978
rect -53578 13978 -53562 13995
rect -52720 13995 -51904 14011
rect -52720 13978 -52704 13995
rect -53578 13961 -53170 13978
rect -54770 13914 -53170 13961
rect -53112 13961 -52704 13978
rect -51920 13978 -51904 13995
rect -51062 13995 -50246 14011
rect -51062 13978 -51046 13995
rect -51920 13961 -51512 13978
rect -53112 13914 -51512 13961
rect -51454 13961 -51046 13978
rect -50262 13978 -50246 13995
rect -49404 13995 -48588 14011
rect -49404 13978 -49388 13995
rect -50262 13961 -49854 13978
rect -51454 13914 -49854 13961
rect -49796 13961 -49388 13978
rect -48604 13978 -48588 13995
rect -47746 13995 -46930 14011
rect -47746 13978 -47730 13995
rect -48604 13961 -48196 13978
rect -49796 13914 -48196 13961
rect -48138 13961 -47730 13978
rect -46946 13978 -46930 13995
rect -46088 13995 -45272 14011
rect -46088 13978 -46072 13995
rect -46946 13961 -46538 13978
rect -48138 13914 -46538 13961
rect -46480 13961 -46072 13978
rect -45288 13978 -45272 13995
rect -44430 13995 -43614 14011
rect -44430 13978 -44414 13995
rect -45288 13961 -44880 13978
rect -46480 13914 -44880 13961
rect -44822 13961 -44414 13978
rect -43630 13978 -43614 13995
rect -42772 13995 -41956 14011
rect -42772 13978 -42756 13995
rect -43630 13961 -43222 13978
rect -44822 13914 -43222 13961
rect -43164 13961 -42756 13978
rect -41972 13978 -41956 13995
rect -41114 13995 -40298 14011
rect -41114 13978 -41098 13995
rect -41972 13961 -41564 13978
rect -43164 13914 -41564 13961
rect -41506 13961 -41098 13978
rect -40314 13978 -40298 13995
rect -39456 13995 -38640 14011
rect -39456 13978 -39440 13995
rect -40314 13961 -39906 13978
rect -41506 13914 -39906 13961
rect -39848 13961 -39440 13978
rect -38656 13978 -38640 13995
rect -37798 13995 -36982 14011
rect -37798 13978 -37782 13995
rect -38656 13961 -38248 13978
rect -39848 13914 -38248 13961
rect -38190 13961 -37782 13978
rect -36998 13978 -36982 13995
rect -36140 13995 -35324 14011
rect -36140 13978 -36124 13995
rect -36998 13961 -36590 13978
rect -38190 13914 -36590 13961
rect -36532 13961 -36124 13978
rect -35340 13978 -35324 13995
rect -34482 13995 -33666 14011
rect -34482 13978 -34466 13995
rect -35340 13961 -34932 13978
rect -36532 13914 -34932 13961
rect -34874 13961 -34466 13978
rect -33682 13978 -33666 13995
rect -32824 13995 -32008 14011
rect -32824 13978 -32808 13995
rect -33682 13961 -33274 13978
rect -34874 13914 -33274 13961
rect -33216 13961 -32808 13978
rect -32024 13978 -32008 13995
rect -31166 13995 -30350 14011
rect -31166 13978 -31150 13995
rect -32024 13961 -31616 13978
rect -33216 13914 -31616 13961
rect -31558 13961 -31150 13978
rect -30366 13978 -30350 13995
rect -29508 13995 -28692 14011
rect -29508 13978 -29492 13995
rect -30366 13961 -29958 13978
rect -31558 13914 -29958 13961
rect -29900 13961 -29492 13978
rect -28708 13978 -28692 13995
rect -28708 13961 -28300 13978
rect -29900 13914 -28300 13961
rect -94562 12467 -92962 12514
rect -94562 12450 -94154 12467
rect -94170 12433 -94154 12450
rect -93370 12450 -92962 12467
rect -92904 12467 -91304 12514
rect -92904 12450 -92496 12467
rect -93370 12433 -93354 12450
rect -94170 12417 -93354 12433
rect -92512 12433 -92496 12450
rect -91712 12450 -91304 12467
rect -91246 12467 -89646 12514
rect -91246 12450 -90838 12467
rect -91712 12433 -91696 12450
rect -92512 12417 -91696 12433
rect -90854 12433 -90838 12450
rect -90054 12450 -89646 12467
rect -89588 12467 -87988 12514
rect -89588 12450 -89180 12467
rect -90054 12433 -90038 12450
rect -90854 12417 -90038 12433
rect -89196 12433 -89180 12450
rect -88396 12450 -87988 12467
rect -87930 12467 -86330 12514
rect -87930 12450 -87522 12467
rect -88396 12433 -88380 12450
rect -89196 12417 -88380 12433
rect -87538 12433 -87522 12450
rect -86738 12450 -86330 12467
rect -86272 12467 -84672 12514
rect -86272 12450 -85864 12467
rect -86738 12433 -86722 12450
rect -87538 12417 -86722 12433
rect -85880 12433 -85864 12450
rect -85080 12450 -84672 12467
rect -84614 12467 -83014 12514
rect -84614 12450 -84206 12467
rect -85080 12433 -85064 12450
rect -85880 12417 -85064 12433
rect -84222 12433 -84206 12450
rect -83422 12450 -83014 12467
rect -82956 12467 -81356 12514
rect -82956 12450 -82548 12467
rect -83422 12433 -83406 12450
rect -84222 12417 -83406 12433
rect -82564 12433 -82548 12450
rect -81764 12450 -81356 12467
rect -81298 12467 -79698 12514
rect -81298 12450 -80890 12467
rect -81764 12433 -81748 12450
rect -82564 12417 -81748 12433
rect -80906 12433 -80890 12450
rect -80106 12450 -79698 12467
rect -79640 12467 -78040 12514
rect -79640 12450 -79232 12467
rect -80106 12433 -80090 12450
rect -80906 12417 -80090 12433
rect -79248 12433 -79232 12450
rect -78448 12450 -78040 12467
rect -77982 12467 -76382 12514
rect -77982 12450 -77574 12467
rect -78448 12433 -78432 12450
rect -79248 12417 -78432 12433
rect -77590 12433 -77574 12450
rect -76790 12450 -76382 12467
rect -76324 12467 -74724 12514
rect -76324 12450 -75916 12467
rect -76790 12433 -76774 12450
rect -77590 12417 -76774 12433
rect -75932 12433 -75916 12450
rect -75132 12450 -74724 12467
rect -74666 12467 -73066 12514
rect -74666 12450 -74258 12467
rect -75132 12433 -75116 12450
rect -75932 12417 -75116 12433
rect -74274 12433 -74258 12450
rect -73474 12450 -73066 12467
rect -73008 12467 -71408 12514
rect -73008 12450 -72600 12467
rect -73474 12433 -73458 12450
rect -74274 12417 -73458 12433
rect -72616 12433 -72600 12450
rect -71816 12450 -71408 12467
rect -71350 12467 -69750 12514
rect -71350 12450 -70942 12467
rect -71816 12433 -71800 12450
rect -72616 12417 -71800 12433
rect -70958 12433 -70942 12450
rect -70158 12450 -69750 12467
rect -69692 12467 -68092 12514
rect -69692 12450 -69284 12467
rect -70158 12433 -70142 12450
rect -70958 12417 -70142 12433
rect -69300 12433 -69284 12450
rect -68500 12450 -68092 12467
rect -68034 12467 -66434 12514
rect -68034 12450 -67626 12467
rect -68500 12433 -68484 12450
rect -69300 12417 -68484 12433
rect -67642 12433 -67626 12450
rect -66842 12450 -66434 12467
rect -66376 12467 -64776 12514
rect -66376 12450 -65968 12467
rect -66842 12433 -66826 12450
rect -67642 12417 -66826 12433
rect -65984 12433 -65968 12450
rect -65184 12450 -64776 12467
rect -64718 12467 -63118 12514
rect -64718 12450 -64310 12467
rect -65184 12433 -65168 12450
rect -65984 12417 -65168 12433
rect -64326 12433 -64310 12450
rect -63526 12450 -63118 12467
rect -63060 12467 -61460 12514
rect -63060 12450 -62652 12467
rect -63526 12433 -63510 12450
rect -64326 12417 -63510 12433
rect -62668 12433 -62652 12450
rect -61868 12450 -61460 12467
rect -61402 12467 -59802 12514
rect -61402 12450 -60994 12467
rect -61868 12433 -61852 12450
rect -62668 12417 -61852 12433
rect -61010 12433 -60994 12450
rect -60210 12450 -59802 12467
rect -59744 12467 -58144 12514
rect -59744 12450 -59336 12467
rect -60210 12433 -60194 12450
rect -61010 12417 -60194 12433
rect -59352 12433 -59336 12450
rect -58552 12450 -58144 12467
rect -58086 12467 -56486 12514
rect -58086 12450 -57678 12467
rect -58552 12433 -58536 12450
rect -59352 12417 -58536 12433
rect -57694 12433 -57678 12450
rect -56894 12450 -56486 12467
rect -56428 12467 -54828 12514
rect -56428 12450 -56020 12467
rect -56894 12433 -56878 12450
rect -57694 12417 -56878 12433
rect -56036 12433 -56020 12450
rect -55236 12450 -54828 12467
rect -54770 12467 -53170 12514
rect -54770 12450 -54362 12467
rect -55236 12433 -55220 12450
rect -56036 12417 -55220 12433
rect -54378 12433 -54362 12450
rect -53578 12450 -53170 12467
rect -53112 12467 -51512 12514
rect -53112 12450 -52704 12467
rect -53578 12433 -53562 12450
rect -54378 12417 -53562 12433
rect -52720 12433 -52704 12450
rect -51920 12450 -51512 12467
rect -51454 12467 -49854 12514
rect -51454 12450 -51046 12467
rect -51920 12433 -51904 12450
rect -52720 12417 -51904 12433
rect -51062 12433 -51046 12450
rect -50262 12450 -49854 12467
rect -49796 12467 -48196 12514
rect -49796 12450 -49388 12467
rect -50262 12433 -50246 12450
rect -51062 12417 -50246 12433
rect -49404 12433 -49388 12450
rect -48604 12450 -48196 12467
rect -48138 12467 -46538 12514
rect -48138 12450 -47730 12467
rect -48604 12433 -48588 12450
rect -49404 12417 -48588 12433
rect -47746 12433 -47730 12450
rect -46946 12450 -46538 12467
rect -46480 12467 -44880 12514
rect -46480 12450 -46072 12467
rect -46946 12433 -46930 12450
rect -47746 12417 -46930 12433
rect -46088 12433 -46072 12450
rect -45288 12450 -44880 12467
rect -44822 12467 -43222 12514
rect -44822 12450 -44414 12467
rect -45288 12433 -45272 12450
rect -46088 12417 -45272 12433
rect -44430 12433 -44414 12450
rect -43630 12450 -43222 12467
rect -43164 12467 -41564 12514
rect -43164 12450 -42756 12467
rect -43630 12433 -43614 12450
rect -44430 12417 -43614 12433
rect -42772 12433 -42756 12450
rect -41972 12450 -41564 12467
rect -41506 12467 -39906 12514
rect -41506 12450 -41098 12467
rect -41972 12433 -41956 12450
rect -42772 12417 -41956 12433
rect -41114 12433 -41098 12450
rect -40314 12450 -39906 12467
rect -39848 12467 -38248 12514
rect -39848 12450 -39440 12467
rect -40314 12433 -40298 12450
rect -41114 12417 -40298 12433
rect -39456 12433 -39440 12450
rect -38656 12450 -38248 12467
rect -38190 12467 -36590 12514
rect -38190 12450 -37782 12467
rect -38656 12433 -38640 12450
rect -39456 12417 -38640 12433
rect -37798 12433 -37782 12450
rect -36998 12450 -36590 12467
rect -36532 12467 -34932 12514
rect -36532 12450 -36124 12467
rect -36998 12433 -36982 12450
rect -37798 12417 -36982 12433
rect -36140 12433 -36124 12450
rect -35340 12450 -34932 12467
rect -34874 12467 -33274 12514
rect -34874 12450 -34466 12467
rect -35340 12433 -35324 12450
rect -36140 12417 -35324 12433
rect -34482 12433 -34466 12450
rect -33682 12450 -33274 12467
rect -33216 12467 -31616 12514
rect -33216 12450 -32808 12467
rect -33682 12433 -33666 12450
rect -34482 12417 -33666 12433
rect -32824 12433 -32808 12450
rect -32024 12450 -31616 12467
rect -31558 12467 -29958 12514
rect -31558 12450 -31150 12467
rect -32024 12433 -32008 12450
rect -32824 12417 -32008 12433
rect -31166 12433 -31150 12450
rect -30366 12450 -29958 12467
rect -29900 12467 -28300 12514
rect -29900 12450 -29492 12467
rect -30366 12433 -30350 12450
rect -31166 12417 -30350 12433
rect -29508 12433 -29492 12450
rect -28708 12450 -28300 12467
rect -28708 12433 -28692 12450
rect -29508 12417 -28692 12433
rect -94170 12359 -93354 12375
rect -94170 12342 -94154 12359
rect -94562 12325 -94154 12342
rect -93370 12342 -93354 12359
rect -92512 12359 -91696 12375
rect -92512 12342 -92496 12359
rect -93370 12325 -92962 12342
rect -94562 12278 -92962 12325
rect -92904 12325 -92496 12342
rect -91712 12342 -91696 12359
rect -90854 12359 -90038 12375
rect -90854 12342 -90838 12359
rect -91712 12325 -91304 12342
rect -92904 12278 -91304 12325
rect -91246 12325 -90838 12342
rect -90054 12342 -90038 12359
rect -89196 12359 -88380 12375
rect -89196 12342 -89180 12359
rect -90054 12325 -89646 12342
rect -91246 12278 -89646 12325
rect -89588 12325 -89180 12342
rect -88396 12342 -88380 12359
rect -87538 12359 -86722 12375
rect -87538 12342 -87522 12359
rect -88396 12325 -87988 12342
rect -89588 12278 -87988 12325
rect -87930 12325 -87522 12342
rect -86738 12342 -86722 12359
rect -85880 12359 -85064 12375
rect -85880 12342 -85864 12359
rect -86738 12325 -86330 12342
rect -87930 12278 -86330 12325
rect -86272 12325 -85864 12342
rect -85080 12342 -85064 12359
rect -84222 12359 -83406 12375
rect -84222 12342 -84206 12359
rect -85080 12325 -84672 12342
rect -86272 12278 -84672 12325
rect -84614 12325 -84206 12342
rect -83422 12342 -83406 12359
rect -82564 12359 -81748 12375
rect -82564 12342 -82548 12359
rect -83422 12325 -83014 12342
rect -84614 12278 -83014 12325
rect -82956 12325 -82548 12342
rect -81764 12342 -81748 12359
rect -80906 12359 -80090 12375
rect -80906 12342 -80890 12359
rect -81764 12325 -81356 12342
rect -82956 12278 -81356 12325
rect -81298 12325 -80890 12342
rect -80106 12342 -80090 12359
rect -79248 12359 -78432 12375
rect -79248 12342 -79232 12359
rect -80106 12325 -79698 12342
rect -81298 12278 -79698 12325
rect -79640 12325 -79232 12342
rect -78448 12342 -78432 12359
rect -77590 12359 -76774 12375
rect -77590 12342 -77574 12359
rect -78448 12325 -78040 12342
rect -79640 12278 -78040 12325
rect -77982 12325 -77574 12342
rect -76790 12342 -76774 12359
rect -75932 12359 -75116 12375
rect -75932 12342 -75916 12359
rect -76790 12325 -76382 12342
rect -77982 12278 -76382 12325
rect -76324 12325 -75916 12342
rect -75132 12342 -75116 12359
rect -74274 12359 -73458 12375
rect -74274 12342 -74258 12359
rect -75132 12325 -74724 12342
rect -76324 12278 -74724 12325
rect -74666 12325 -74258 12342
rect -73474 12342 -73458 12359
rect -72616 12359 -71800 12375
rect -72616 12342 -72600 12359
rect -73474 12325 -73066 12342
rect -74666 12278 -73066 12325
rect -73008 12325 -72600 12342
rect -71816 12342 -71800 12359
rect -70958 12359 -70142 12375
rect -70958 12342 -70942 12359
rect -71816 12325 -71408 12342
rect -73008 12278 -71408 12325
rect -71350 12325 -70942 12342
rect -70158 12342 -70142 12359
rect -69300 12359 -68484 12375
rect -69300 12342 -69284 12359
rect -70158 12325 -69750 12342
rect -71350 12278 -69750 12325
rect -69692 12325 -69284 12342
rect -68500 12342 -68484 12359
rect -67642 12359 -66826 12375
rect -67642 12342 -67626 12359
rect -68500 12325 -68092 12342
rect -69692 12278 -68092 12325
rect -68034 12325 -67626 12342
rect -66842 12342 -66826 12359
rect -65984 12359 -65168 12375
rect -65984 12342 -65968 12359
rect -66842 12325 -66434 12342
rect -68034 12278 -66434 12325
rect -66376 12325 -65968 12342
rect -65184 12342 -65168 12359
rect -64326 12359 -63510 12375
rect -64326 12342 -64310 12359
rect -65184 12325 -64776 12342
rect -66376 12278 -64776 12325
rect -64718 12325 -64310 12342
rect -63526 12342 -63510 12359
rect -62668 12359 -61852 12375
rect -62668 12342 -62652 12359
rect -63526 12325 -63118 12342
rect -64718 12278 -63118 12325
rect -63060 12325 -62652 12342
rect -61868 12342 -61852 12359
rect -61010 12359 -60194 12375
rect -61010 12342 -60994 12359
rect -61868 12325 -61460 12342
rect -63060 12278 -61460 12325
rect -61402 12325 -60994 12342
rect -60210 12342 -60194 12359
rect -59352 12359 -58536 12375
rect -59352 12342 -59336 12359
rect -60210 12325 -59802 12342
rect -61402 12278 -59802 12325
rect -59744 12325 -59336 12342
rect -58552 12342 -58536 12359
rect -57694 12359 -56878 12375
rect -57694 12342 -57678 12359
rect -58552 12325 -58144 12342
rect -59744 12278 -58144 12325
rect -58086 12325 -57678 12342
rect -56894 12342 -56878 12359
rect -56036 12359 -55220 12375
rect -56036 12342 -56020 12359
rect -56894 12325 -56486 12342
rect -58086 12278 -56486 12325
rect -56428 12325 -56020 12342
rect -55236 12342 -55220 12359
rect -54378 12359 -53562 12375
rect -54378 12342 -54362 12359
rect -55236 12325 -54828 12342
rect -56428 12278 -54828 12325
rect -54770 12325 -54362 12342
rect -53578 12342 -53562 12359
rect -52720 12359 -51904 12375
rect -52720 12342 -52704 12359
rect -53578 12325 -53170 12342
rect -54770 12278 -53170 12325
rect -53112 12325 -52704 12342
rect -51920 12342 -51904 12359
rect -51062 12359 -50246 12375
rect -51062 12342 -51046 12359
rect -51920 12325 -51512 12342
rect -53112 12278 -51512 12325
rect -51454 12325 -51046 12342
rect -50262 12342 -50246 12359
rect -49404 12359 -48588 12375
rect -49404 12342 -49388 12359
rect -50262 12325 -49854 12342
rect -51454 12278 -49854 12325
rect -49796 12325 -49388 12342
rect -48604 12342 -48588 12359
rect -47746 12359 -46930 12375
rect -47746 12342 -47730 12359
rect -48604 12325 -48196 12342
rect -49796 12278 -48196 12325
rect -48138 12325 -47730 12342
rect -46946 12342 -46930 12359
rect -46088 12359 -45272 12375
rect -46088 12342 -46072 12359
rect -46946 12325 -46538 12342
rect -48138 12278 -46538 12325
rect -46480 12325 -46072 12342
rect -45288 12342 -45272 12359
rect -44430 12359 -43614 12375
rect -44430 12342 -44414 12359
rect -45288 12325 -44880 12342
rect -46480 12278 -44880 12325
rect -44822 12325 -44414 12342
rect -43630 12342 -43614 12359
rect -42772 12359 -41956 12375
rect -42772 12342 -42756 12359
rect -43630 12325 -43222 12342
rect -44822 12278 -43222 12325
rect -43164 12325 -42756 12342
rect -41972 12342 -41956 12359
rect -41114 12359 -40298 12375
rect -41114 12342 -41098 12359
rect -41972 12325 -41564 12342
rect -43164 12278 -41564 12325
rect -41506 12325 -41098 12342
rect -40314 12342 -40298 12359
rect -39456 12359 -38640 12375
rect -39456 12342 -39440 12359
rect -40314 12325 -39906 12342
rect -41506 12278 -39906 12325
rect -39848 12325 -39440 12342
rect -38656 12342 -38640 12359
rect -37798 12359 -36982 12375
rect -37798 12342 -37782 12359
rect -38656 12325 -38248 12342
rect -39848 12278 -38248 12325
rect -38190 12325 -37782 12342
rect -36998 12342 -36982 12359
rect -36140 12359 -35324 12375
rect -36140 12342 -36124 12359
rect -36998 12325 -36590 12342
rect -38190 12278 -36590 12325
rect -36532 12325 -36124 12342
rect -35340 12342 -35324 12359
rect -34482 12359 -33666 12375
rect -34482 12342 -34466 12359
rect -35340 12325 -34932 12342
rect -36532 12278 -34932 12325
rect -34874 12325 -34466 12342
rect -33682 12342 -33666 12359
rect -32824 12359 -32008 12375
rect -32824 12342 -32808 12359
rect -33682 12325 -33274 12342
rect -34874 12278 -33274 12325
rect -33216 12325 -32808 12342
rect -32024 12342 -32008 12359
rect -31166 12359 -30350 12375
rect -31166 12342 -31150 12359
rect -32024 12325 -31616 12342
rect -33216 12278 -31616 12325
rect -31558 12325 -31150 12342
rect -30366 12342 -30350 12359
rect -29508 12359 -28692 12375
rect -29508 12342 -29492 12359
rect -30366 12325 -29958 12342
rect -31558 12278 -29958 12325
rect -29900 12325 -29492 12342
rect -28708 12342 -28692 12359
rect -28708 12325 -28300 12342
rect -29900 12278 -28300 12325
rect -94562 10831 -92962 10878
rect -94562 10814 -94154 10831
rect -94170 10797 -94154 10814
rect -93370 10814 -92962 10831
rect -92904 10831 -91304 10878
rect -92904 10814 -92496 10831
rect -93370 10797 -93354 10814
rect -94170 10781 -93354 10797
rect -92512 10797 -92496 10814
rect -91712 10814 -91304 10831
rect -91246 10831 -89646 10878
rect -91246 10814 -90838 10831
rect -91712 10797 -91696 10814
rect -92512 10781 -91696 10797
rect -90854 10797 -90838 10814
rect -90054 10814 -89646 10831
rect -89588 10831 -87988 10878
rect -89588 10814 -89180 10831
rect -90054 10797 -90038 10814
rect -90854 10781 -90038 10797
rect -89196 10797 -89180 10814
rect -88396 10814 -87988 10831
rect -87930 10831 -86330 10878
rect -87930 10814 -87522 10831
rect -88396 10797 -88380 10814
rect -89196 10781 -88380 10797
rect -87538 10797 -87522 10814
rect -86738 10814 -86330 10831
rect -86272 10831 -84672 10878
rect -86272 10814 -85864 10831
rect -86738 10797 -86722 10814
rect -87538 10781 -86722 10797
rect -85880 10797 -85864 10814
rect -85080 10814 -84672 10831
rect -84614 10831 -83014 10878
rect -84614 10814 -84206 10831
rect -85080 10797 -85064 10814
rect -85880 10781 -85064 10797
rect -84222 10797 -84206 10814
rect -83422 10814 -83014 10831
rect -82956 10831 -81356 10878
rect -82956 10814 -82548 10831
rect -83422 10797 -83406 10814
rect -84222 10781 -83406 10797
rect -82564 10797 -82548 10814
rect -81764 10814 -81356 10831
rect -81298 10831 -79698 10878
rect -81298 10814 -80890 10831
rect -81764 10797 -81748 10814
rect -82564 10781 -81748 10797
rect -80906 10797 -80890 10814
rect -80106 10814 -79698 10831
rect -79640 10831 -78040 10878
rect -79640 10814 -79232 10831
rect -80106 10797 -80090 10814
rect -80906 10781 -80090 10797
rect -79248 10797 -79232 10814
rect -78448 10814 -78040 10831
rect -77982 10831 -76382 10878
rect -77982 10814 -77574 10831
rect -78448 10797 -78432 10814
rect -79248 10781 -78432 10797
rect -77590 10797 -77574 10814
rect -76790 10814 -76382 10831
rect -76324 10831 -74724 10878
rect -76324 10814 -75916 10831
rect -76790 10797 -76774 10814
rect -77590 10781 -76774 10797
rect -75932 10797 -75916 10814
rect -75132 10814 -74724 10831
rect -74666 10831 -73066 10878
rect -74666 10814 -74258 10831
rect -75132 10797 -75116 10814
rect -75932 10781 -75116 10797
rect -74274 10797 -74258 10814
rect -73474 10814 -73066 10831
rect -73008 10831 -71408 10878
rect -73008 10814 -72600 10831
rect -73474 10797 -73458 10814
rect -74274 10781 -73458 10797
rect -72616 10797 -72600 10814
rect -71816 10814 -71408 10831
rect -71350 10831 -69750 10878
rect -71350 10814 -70942 10831
rect -71816 10797 -71800 10814
rect -72616 10781 -71800 10797
rect -70958 10797 -70942 10814
rect -70158 10814 -69750 10831
rect -69692 10831 -68092 10878
rect -69692 10814 -69284 10831
rect -70158 10797 -70142 10814
rect -70958 10781 -70142 10797
rect -69300 10797 -69284 10814
rect -68500 10814 -68092 10831
rect -68034 10831 -66434 10878
rect -68034 10814 -67626 10831
rect -68500 10797 -68484 10814
rect -69300 10781 -68484 10797
rect -67642 10797 -67626 10814
rect -66842 10814 -66434 10831
rect -66376 10831 -64776 10878
rect -66376 10814 -65968 10831
rect -66842 10797 -66826 10814
rect -67642 10781 -66826 10797
rect -65984 10797 -65968 10814
rect -65184 10814 -64776 10831
rect -64718 10831 -63118 10878
rect -64718 10814 -64310 10831
rect -65184 10797 -65168 10814
rect -65984 10781 -65168 10797
rect -64326 10797 -64310 10814
rect -63526 10814 -63118 10831
rect -63060 10831 -61460 10878
rect -63060 10814 -62652 10831
rect -63526 10797 -63510 10814
rect -64326 10781 -63510 10797
rect -62668 10797 -62652 10814
rect -61868 10814 -61460 10831
rect -61402 10831 -59802 10878
rect -61402 10814 -60994 10831
rect -61868 10797 -61852 10814
rect -62668 10781 -61852 10797
rect -61010 10797 -60994 10814
rect -60210 10814 -59802 10831
rect -59744 10831 -58144 10878
rect -59744 10814 -59336 10831
rect -60210 10797 -60194 10814
rect -61010 10781 -60194 10797
rect -59352 10797 -59336 10814
rect -58552 10814 -58144 10831
rect -58086 10831 -56486 10878
rect -58086 10814 -57678 10831
rect -58552 10797 -58536 10814
rect -59352 10781 -58536 10797
rect -57694 10797 -57678 10814
rect -56894 10814 -56486 10831
rect -56428 10831 -54828 10878
rect -56428 10814 -56020 10831
rect -56894 10797 -56878 10814
rect -57694 10781 -56878 10797
rect -56036 10797 -56020 10814
rect -55236 10814 -54828 10831
rect -54770 10831 -53170 10878
rect -54770 10814 -54362 10831
rect -55236 10797 -55220 10814
rect -56036 10781 -55220 10797
rect -54378 10797 -54362 10814
rect -53578 10814 -53170 10831
rect -53112 10831 -51512 10878
rect -53112 10814 -52704 10831
rect -53578 10797 -53562 10814
rect -54378 10781 -53562 10797
rect -52720 10797 -52704 10814
rect -51920 10814 -51512 10831
rect -51454 10831 -49854 10878
rect -51454 10814 -51046 10831
rect -51920 10797 -51904 10814
rect -52720 10781 -51904 10797
rect -51062 10797 -51046 10814
rect -50262 10814 -49854 10831
rect -49796 10831 -48196 10878
rect -49796 10814 -49388 10831
rect -50262 10797 -50246 10814
rect -51062 10781 -50246 10797
rect -49404 10797 -49388 10814
rect -48604 10814 -48196 10831
rect -48138 10831 -46538 10878
rect -48138 10814 -47730 10831
rect -48604 10797 -48588 10814
rect -49404 10781 -48588 10797
rect -47746 10797 -47730 10814
rect -46946 10814 -46538 10831
rect -46480 10831 -44880 10878
rect -46480 10814 -46072 10831
rect -46946 10797 -46930 10814
rect -47746 10781 -46930 10797
rect -46088 10797 -46072 10814
rect -45288 10814 -44880 10831
rect -44822 10831 -43222 10878
rect -44822 10814 -44414 10831
rect -45288 10797 -45272 10814
rect -46088 10781 -45272 10797
rect -44430 10797 -44414 10814
rect -43630 10814 -43222 10831
rect -43164 10831 -41564 10878
rect -43164 10814 -42756 10831
rect -43630 10797 -43614 10814
rect -44430 10781 -43614 10797
rect -42772 10797 -42756 10814
rect -41972 10814 -41564 10831
rect -41506 10831 -39906 10878
rect -41506 10814 -41098 10831
rect -41972 10797 -41956 10814
rect -42772 10781 -41956 10797
rect -41114 10797 -41098 10814
rect -40314 10814 -39906 10831
rect -39848 10831 -38248 10878
rect -39848 10814 -39440 10831
rect -40314 10797 -40298 10814
rect -41114 10781 -40298 10797
rect -39456 10797 -39440 10814
rect -38656 10814 -38248 10831
rect -38190 10831 -36590 10878
rect -38190 10814 -37782 10831
rect -38656 10797 -38640 10814
rect -39456 10781 -38640 10797
rect -37798 10797 -37782 10814
rect -36998 10814 -36590 10831
rect -36532 10831 -34932 10878
rect -36532 10814 -36124 10831
rect -36998 10797 -36982 10814
rect -37798 10781 -36982 10797
rect -36140 10797 -36124 10814
rect -35340 10814 -34932 10831
rect -34874 10831 -33274 10878
rect -34874 10814 -34466 10831
rect -35340 10797 -35324 10814
rect -36140 10781 -35324 10797
rect -34482 10797 -34466 10814
rect -33682 10814 -33274 10831
rect -33216 10831 -31616 10878
rect -33216 10814 -32808 10831
rect -33682 10797 -33666 10814
rect -34482 10781 -33666 10797
rect -32824 10797 -32808 10814
rect -32024 10814 -31616 10831
rect -31558 10831 -29958 10878
rect -31558 10814 -31150 10831
rect -32024 10797 -32008 10814
rect -32824 10781 -32008 10797
rect -31166 10797 -31150 10814
rect -30366 10814 -29958 10831
rect -29900 10831 -28300 10878
rect -29900 10814 -29492 10831
rect -30366 10797 -30350 10814
rect -31166 10781 -30350 10797
rect -29508 10797 -29492 10814
rect -28708 10814 -28300 10831
rect -28708 10797 -28692 10814
rect -29508 10781 -28692 10797
rect -94170 10721 -93354 10737
rect -94170 10704 -94154 10721
rect -94562 10687 -94154 10704
rect -93370 10704 -93354 10721
rect -92512 10721 -91696 10737
rect -92512 10704 -92496 10721
rect -93370 10687 -92962 10704
rect -94562 10640 -92962 10687
rect -92904 10687 -92496 10704
rect -91712 10704 -91696 10721
rect -90854 10721 -90038 10737
rect -90854 10704 -90838 10721
rect -91712 10687 -91304 10704
rect -92904 10640 -91304 10687
rect -91246 10687 -90838 10704
rect -90054 10704 -90038 10721
rect -89196 10721 -88380 10737
rect -89196 10704 -89180 10721
rect -90054 10687 -89646 10704
rect -91246 10640 -89646 10687
rect -89588 10687 -89180 10704
rect -88396 10704 -88380 10721
rect -87538 10721 -86722 10737
rect -87538 10704 -87522 10721
rect -88396 10687 -87988 10704
rect -89588 10640 -87988 10687
rect -87930 10687 -87522 10704
rect -86738 10704 -86722 10721
rect -85880 10721 -85064 10737
rect -85880 10704 -85864 10721
rect -86738 10687 -86330 10704
rect -87930 10640 -86330 10687
rect -86272 10687 -85864 10704
rect -85080 10704 -85064 10721
rect -84222 10721 -83406 10737
rect -84222 10704 -84206 10721
rect -85080 10687 -84672 10704
rect -86272 10640 -84672 10687
rect -84614 10687 -84206 10704
rect -83422 10704 -83406 10721
rect -82564 10721 -81748 10737
rect -82564 10704 -82548 10721
rect -83422 10687 -83014 10704
rect -84614 10640 -83014 10687
rect -82956 10687 -82548 10704
rect -81764 10704 -81748 10721
rect -80906 10721 -80090 10737
rect -80906 10704 -80890 10721
rect -81764 10687 -81356 10704
rect -82956 10640 -81356 10687
rect -81298 10687 -80890 10704
rect -80106 10704 -80090 10721
rect -79248 10721 -78432 10737
rect -79248 10704 -79232 10721
rect -80106 10687 -79698 10704
rect -81298 10640 -79698 10687
rect -79640 10687 -79232 10704
rect -78448 10704 -78432 10721
rect -77590 10721 -76774 10737
rect -77590 10704 -77574 10721
rect -78448 10687 -78040 10704
rect -79640 10640 -78040 10687
rect -77982 10687 -77574 10704
rect -76790 10704 -76774 10721
rect -75932 10721 -75116 10737
rect -75932 10704 -75916 10721
rect -76790 10687 -76382 10704
rect -77982 10640 -76382 10687
rect -76324 10687 -75916 10704
rect -75132 10704 -75116 10721
rect -74274 10721 -73458 10737
rect -74274 10704 -74258 10721
rect -75132 10687 -74724 10704
rect -76324 10640 -74724 10687
rect -74666 10687 -74258 10704
rect -73474 10704 -73458 10721
rect -72616 10721 -71800 10737
rect -72616 10704 -72600 10721
rect -73474 10687 -73066 10704
rect -74666 10640 -73066 10687
rect -73008 10687 -72600 10704
rect -71816 10704 -71800 10721
rect -70958 10721 -70142 10737
rect -70958 10704 -70942 10721
rect -71816 10687 -71408 10704
rect -73008 10640 -71408 10687
rect -71350 10687 -70942 10704
rect -70158 10704 -70142 10721
rect -69300 10721 -68484 10737
rect -69300 10704 -69284 10721
rect -70158 10687 -69750 10704
rect -71350 10640 -69750 10687
rect -69692 10687 -69284 10704
rect -68500 10704 -68484 10721
rect -67642 10721 -66826 10737
rect -67642 10704 -67626 10721
rect -68500 10687 -68092 10704
rect -69692 10640 -68092 10687
rect -68034 10687 -67626 10704
rect -66842 10704 -66826 10721
rect -65984 10721 -65168 10737
rect -65984 10704 -65968 10721
rect -66842 10687 -66434 10704
rect -68034 10640 -66434 10687
rect -66376 10687 -65968 10704
rect -65184 10704 -65168 10721
rect -64326 10721 -63510 10737
rect -64326 10704 -64310 10721
rect -65184 10687 -64776 10704
rect -66376 10640 -64776 10687
rect -64718 10687 -64310 10704
rect -63526 10704 -63510 10721
rect -62668 10721 -61852 10737
rect -62668 10704 -62652 10721
rect -63526 10687 -63118 10704
rect -64718 10640 -63118 10687
rect -63060 10687 -62652 10704
rect -61868 10704 -61852 10721
rect -61010 10721 -60194 10737
rect -61010 10704 -60994 10721
rect -61868 10687 -61460 10704
rect -63060 10640 -61460 10687
rect -61402 10687 -60994 10704
rect -60210 10704 -60194 10721
rect -59352 10721 -58536 10737
rect -59352 10704 -59336 10721
rect -60210 10687 -59802 10704
rect -61402 10640 -59802 10687
rect -59744 10687 -59336 10704
rect -58552 10704 -58536 10721
rect -57694 10721 -56878 10737
rect -57694 10704 -57678 10721
rect -58552 10687 -58144 10704
rect -59744 10640 -58144 10687
rect -58086 10687 -57678 10704
rect -56894 10704 -56878 10721
rect -56036 10721 -55220 10737
rect -56036 10704 -56020 10721
rect -56894 10687 -56486 10704
rect -58086 10640 -56486 10687
rect -56428 10687 -56020 10704
rect -55236 10704 -55220 10721
rect -54378 10721 -53562 10737
rect -54378 10704 -54362 10721
rect -55236 10687 -54828 10704
rect -56428 10640 -54828 10687
rect -54770 10687 -54362 10704
rect -53578 10704 -53562 10721
rect -52720 10721 -51904 10737
rect -52720 10704 -52704 10721
rect -53578 10687 -53170 10704
rect -54770 10640 -53170 10687
rect -53112 10687 -52704 10704
rect -51920 10704 -51904 10721
rect -51062 10721 -50246 10737
rect -51062 10704 -51046 10721
rect -51920 10687 -51512 10704
rect -53112 10640 -51512 10687
rect -51454 10687 -51046 10704
rect -50262 10704 -50246 10721
rect -49404 10721 -48588 10737
rect -49404 10704 -49388 10721
rect -50262 10687 -49854 10704
rect -51454 10640 -49854 10687
rect -49796 10687 -49388 10704
rect -48604 10704 -48588 10721
rect -47746 10721 -46930 10737
rect -47746 10704 -47730 10721
rect -48604 10687 -48196 10704
rect -49796 10640 -48196 10687
rect -48138 10687 -47730 10704
rect -46946 10704 -46930 10721
rect -46088 10721 -45272 10737
rect -46088 10704 -46072 10721
rect -46946 10687 -46538 10704
rect -48138 10640 -46538 10687
rect -46480 10687 -46072 10704
rect -45288 10704 -45272 10721
rect -44430 10721 -43614 10737
rect -44430 10704 -44414 10721
rect -45288 10687 -44880 10704
rect -46480 10640 -44880 10687
rect -44822 10687 -44414 10704
rect -43630 10704 -43614 10721
rect -42772 10721 -41956 10737
rect -42772 10704 -42756 10721
rect -43630 10687 -43222 10704
rect -44822 10640 -43222 10687
rect -43164 10687 -42756 10704
rect -41972 10704 -41956 10721
rect -41114 10721 -40298 10737
rect -41114 10704 -41098 10721
rect -41972 10687 -41564 10704
rect -43164 10640 -41564 10687
rect -41506 10687 -41098 10704
rect -40314 10704 -40298 10721
rect -39456 10721 -38640 10737
rect -39456 10704 -39440 10721
rect -40314 10687 -39906 10704
rect -41506 10640 -39906 10687
rect -39848 10687 -39440 10704
rect -38656 10704 -38640 10721
rect -37798 10721 -36982 10737
rect -37798 10704 -37782 10721
rect -38656 10687 -38248 10704
rect -39848 10640 -38248 10687
rect -38190 10687 -37782 10704
rect -36998 10704 -36982 10721
rect -36140 10721 -35324 10737
rect -36140 10704 -36124 10721
rect -36998 10687 -36590 10704
rect -38190 10640 -36590 10687
rect -36532 10687 -36124 10704
rect -35340 10704 -35324 10721
rect -34482 10721 -33666 10737
rect -34482 10704 -34466 10721
rect -35340 10687 -34932 10704
rect -36532 10640 -34932 10687
rect -34874 10687 -34466 10704
rect -33682 10704 -33666 10721
rect -32824 10721 -32008 10737
rect -32824 10704 -32808 10721
rect -33682 10687 -33274 10704
rect -34874 10640 -33274 10687
rect -33216 10687 -32808 10704
rect -32024 10704 -32008 10721
rect -31166 10721 -30350 10737
rect -31166 10704 -31150 10721
rect -32024 10687 -31616 10704
rect -33216 10640 -31616 10687
rect -31558 10687 -31150 10704
rect -30366 10704 -30350 10721
rect -29508 10721 -28692 10737
rect -29508 10704 -29492 10721
rect -30366 10687 -29958 10704
rect -31558 10640 -29958 10687
rect -29900 10687 -29492 10704
rect -28708 10704 -28692 10721
rect -28708 10687 -28300 10704
rect -29900 10640 -28300 10687
rect -94562 9193 -92962 9240
rect -94562 9176 -94154 9193
rect -94170 9159 -94154 9176
rect -93370 9176 -92962 9193
rect -92904 9193 -91304 9240
rect -92904 9176 -92496 9193
rect -93370 9159 -93354 9176
rect -94170 9143 -93354 9159
rect -92512 9159 -92496 9176
rect -91712 9176 -91304 9193
rect -91246 9193 -89646 9240
rect -91246 9176 -90838 9193
rect -91712 9159 -91696 9176
rect -92512 9143 -91696 9159
rect -90854 9159 -90838 9176
rect -90054 9176 -89646 9193
rect -89588 9193 -87988 9240
rect -89588 9176 -89180 9193
rect -90054 9159 -90038 9176
rect -90854 9143 -90038 9159
rect -89196 9159 -89180 9176
rect -88396 9176 -87988 9193
rect -87930 9193 -86330 9240
rect -87930 9176 -87522 9193
rect -88396 9159 -88380 9176
rect -89196 9143 -88380 9159
rect -87538 9159 -87522 9176
rect -86738 9176 -86330 9193
rect -86272 9193 -84672 9240
rect -86272 9176 -85864 9193
rect -86738 9159 -86722 9176
rect -87538 9143 -86722 9159
rect -85880 9159 -85864 9176
rect -85080 9176 -84672 9193
rect -84614 9193 -83014 9240
rect -84614 9176 -84206 9193
rect -85080 9159 -85064 9176
rect -85880 9143 -85064 9159
rect -84222 9159 -84206 9176
rect -83422 9176 -83014 9193
rect -82956 9193 -81356 9240
rect -82956 9176 -82548 9193
rect -83422 9159 -83406 9176
rect -84222 9143 -83406 9159
rect -82564 9159 -82548 9176
rect -81764 9176 -81356 9193
rect -81298 9193 -79698 9240
rect -81298 9176 -80890 9193
rect -81764 9159 -81748 9176
rect -82564 9143 -81748 9159
rect -80906 9159 -80890 9176
rect -80106 9176 -79698 9193
rect -79640 9193 -78040 9240
rect -79640 9176 -79232 9193
rect -80106 9159 -80090 9176
rect -80906 9143 -80090 9159
rect -79248 9159 -79232 9176
rect -78448 9176 -78040 9193
rect -77982 9193 -76382 9240
rect -77982 9176 -77574 9193
rect -78448 9159 -78432 9176
rect -79248 9143 -78432 9159
rect -77590 9159 -77574 9176
rect -76790 9176 -76382 9193
rect -76324 9193 -74724 9240
rect -76324 9176 -75916 9193
rect -76790 9159 -76774 9176
rect -77590 9143 -76774 9159
rect -75932 9159 -75916 9176
rect -75132 9176 -74724 9193
rect -74666 9193 -73066 9240
rect -74666 9176 -74258 9193
rect -75132 9159 -75116 9176
rect -75932 9143 -75116 9159
rect -74274 9159 -74258 9176
rect -73474 9176 -73066 9193
rect -73008 9193 -71408 9240
rect -73008 9176 -72600 9193
rect -73474 9159 -73458 9176
rect -74274 9143 -73458 9159
rect -72616 9159 -72600 9176
rect -71816 9176 -71408 9193
rect -71350 9193 -69750 9240
rect -71350 9176 -70942 9193
rect -71816 9159 -71800 9176
rect -72616 9143 -71800 9159
rect -70958 9159 -70942 9176
rect -70158 9176 -69750 9193
rect -69692 9193 -68092 9240
rect -69692 9176 -69284 9193
rect -70158 9159 -70142 9176
rect -70958 9143 -70142 9159
rect -69300 9159 -69284 9176
rect -68500 9176 -68092 9193
rect -68034 9193 -66434 9240
rect -68034 9176 -67626 9193
rect -68500 9159 -68484 9176
rect -69300 9143 -68484 9159
rect -67642 9159 -67626 9176
rect -66842 9176 -66434 9193
rect -66376 9193 -64776 9240
rect -66376 9176 -65968 9193
rect -66842 9159 -66826 9176
rect -67642 9143 -66826 9159
rect -65984 9159 -65968 9176
rect -65184 9176 -64776 9193
rect -64718 9193 -63118 9240
rect -64718 9176 -64310 9193
rect -65184 9159 -65168 9176
rect -65984 9143 -65168 9159
rect -64326 9159 -64310 9176
rect -63526 9176 -63118 9193
rect -63060 9193 -61460 9240
rect -63060 9176 -62652 9193
rect -63526 9159 -63510 9176
rect -64326 9143 -63510 9159
rect -62668 9159 -62652 9176
rect -61868 9176 -61460 9193
rect -61402 9193 -59802 9240
rect -61402 9176 -60994 9193
rect -61868 9159 -61852 9176
rect -62668 9143 -61852 9159
rect -61010 9159 -60994 9176
rect -60210 9176 -59802 9193
rect -59744 9193 -58144 9240
rect -59744 9176 -59336 9193
rect -60210 9159 -60194 9176
rect -61010 9143 -60194 9159
rect -59352 9159 -59336 9176
rect -58552 9176 -58144 9193
rect -58086 9193 -56486 9240
rect -58086 9176 -57678 9193
rect -58552 9159 -58536 9176
rect -59352 9143 -58536 9159
rect -57694 9159 -57678 9176
rect -56894 9176 -56486 9193
rect -56428 9193 -54828 9240
rect -56428 9176 -56020 9193
rect -56894 9159 -56878 9176
rect -57694 9143 -56878 9159
rect -56036 9159 -56020 9176
rect -55236 9176 -54828 9193
rect -54770 9193 -53170 9240
rect -54770 9176 -54362 9193
rect -55236 9159 -55220 9176
rect -56036 9143 -55220 9159
rect -54378 9159 -54362 9176
rect -53578 9176 -53170 9193
rect -53112 9193 -51512 9240
rect -53112 9176 -52704 9193
rect -53578 9159 -53562 9176
rect -54378 9143 -53562 9159
rect -52720 9159 -52704 9176
rect -51920 9176 -51512 9193
rect -51454 9193 -49854 9240
rect -51454 9176 -51046 9193
rect -51920 9159 -51904 9176
rect -52720 9143 -51904 9159
rect -51062 9159 -51046 9176
rect -50262 9176 -49854 9193
rect -49796 9193 -48196 9240
rect -49796 9176 -49388 9193
rect -50262 9159 -50246 9176
rect -51062 9143 -50246 9159
rect -49404 9159 -49388 9176
rect -48604 9176 -48196 9193
rect -48138 9193 -46538 9240
rect -48138 9176 -47730 9193
rect -48604 9159 -48588 9176
rect -49404 9143 -48588 9159
rect -47746 9159 -47730 9176
rect -46946 9176 -46538 9193
rect -46480 9193 -44880 9240
rect -46480 9176 -46072 9193
rect -46946 9159 -46930 9176
rect -47746 9143 -46930 9159
rect -46088 9159 -46072 9176
rect -45288 9176 -44880 9193
rect -44822 9193 -43222 9240
rect -44822 9176 -44414 9193
rect -45288 9159 -45272 9176
rect -46088 9143 -45272 9159
rect -44430 9159 -44414 9176
rect -43630 9176 -43222 9193
rect -43164 9193 -41564 9240
rect -43164 9176 -42756 9193
rect -43630 9159 -43614 9176
rect -44430 9143 -43614 9159
rect -42772 9159 -42756 9176
rect -41972 9176 -41564 9193
rect -41506 9193 -39906 9240
rect -41506 9176 -41098 9193
rect -41972 9159 -41956 9176
rect -42772 9143 -41956 9159
rect -41114 9159 -41098 9176
rect -40314 9176 -39906 9193
rect -39848 9193 -38248 9240
rect -39848 9176 -39440 9193
rect -40314 9159 -40298 9176
rect -41114 9143 -40298 9159
rect -39456 9159 -39440 9176
rect -38656 9176 -38248 9193
rect -38190 9193 -36590 9240
rect -38190 9176 -37782 9193
rect -38656 9159 -38640 9176
rect -39456 9143 -38640 9159
rect -37798 9159 -37782 9176
rect -36998 9176 -36590 9193
rect -36532 9193 -34932 9240
rect -36532 9176 -36124 9193
rect -36998 9159 -36982 9176
rect -37798 9143 -36982 9159
rect -36140 9159 -36124 9176
rect -35340 9176 -34932 9193
rect -34874 9193 -33274 9240
rect -34874 9176 -34466 9193
rect -35340 9159 -35324 9176
rect -36140 9143 -35324 9159
rect -34482 9159 -34466 9176
rect -33682 9176 -33274 9193
rect -33216 9193 -31616 9240
rect -33216 9176 -32808 9193
rect -33682 9159 -33666 9176
rect -34482 9143 -33666 9159
rect -32824 9159 -32808 9176
rect -32024 9176 -31616 9193
rect -31558 9193 -29958 9240
rect -31558 9176 -31150 9193
rect -32024 9159 -32008 9176
rect -32824 9143 -32008 9159
rect -31166 9159 -31150 9176
rect -30366 9176 -29958 9193
rect -29900 9193 -28300 9240
rect -29900 9176 -29492 9193
rect -30366 9159 -30350 9176
rect -31166 9143 -30350 9159
rect -29508 9159 -29492 9176
rect -28708 9176 -28300 9193
rect -28708 9159 -28692 9176
rect -29508 9143 -28692 9159
rect -94170 9085 -93354 9101
rect -94170 9068 -94154 9085
rect -94562 9051 -94154 9068
rect -93370 9068 -93354 9085
rect -92512 9085 -91696 9101
rect -92512 9068 -92496 9085
rect -93370 9051 -92962 9068
rect -94562 9004 -92962 9051
rect -92904 9051 -92496 9068
rect -91712 9068 -91696 9085
rect -90854 9085 -90038 9101
rect -90854 9068 -90838 9085
rect -91712 9051 -91304 9068
rect -92904 9004 -91304 9051
rect -91246 9051 -90838 9068
rect -90054 9068 -90038 9085
rect -89196 9085 -88380 9101
rect -89196 9068 -89180 9085
rect -90054 9051 -89646 9068
rect -91246 9004 -89646 9051
rect -89588 9051 -89180 9068
rect -88396 9068 -88380 9085
rect -87538 9085 -86722 9101
rect -87538 9068 -87522 9085
rect -88396 9051 -87988 9068
rect -89588 9004 -87988 9051
rect -87930 9051 -87522 9068
rect -86738 9068 -86722 9085
rect -85880 9085 -85064 9101
rect -85880 9068 -85864 9085
rect -86738 9051 -86330 9068
rect -87930 9004 -86330 9051
rect -86272 9051 -85864 9068
rect -85080 9068 -85064 9085
rect -84222 9085 -83406 9101
rect -84222 9068 -84206 9085
rect -85080 9051 -84672 9068
rect -86272 9004 -84672 9051
rect -84614 9051 -84206 9068
rect -83422 9068 -83406 9085
rect -82564 9085 -81748 9101
rect -82564 9068 -82548 9085
rect -83422 9051 -83014 9068
rect -84614 9004 -83014 9051
rect -82956 9051 -82548 9068
rect -81764 9068 -81748 9085
rect -80906 9085 -80090 9101
rect -80906 9068 -80890 9085
rect -81764 9051 -81356 9068
rect -82956 9004 -81356 9051
rect -81298 9051 -80890 9068
rect -80106 9068 -80090 9085
rect -79248 9085 -78432 9101
rect -79248 9068 -79232 9085
rect -80106 9051 -79698 9068
rect -81298 9004 -79698 9051
rect -79640 9051 -79232 9068
rect -78448 9068 -78432 9085
rect -77590 9085 -76774 9101
rect -77590 9068 -77574 9085
rect -78448 9051 -78040 9068
rect -79640 9004 -78040 9051
rect -77982 9051 -77574 9068
rect -76790 9068 -76774 9085
rect -75932 9085 -75116 9101
rect -75932 9068 -75916 9085
rect -76790 9051 -76382 9068
rect -77982 9004 -76382 9051
rect -76324 9051 -75916 9068
rect -75132 9068 -75116 9085
rect -74274 9085 -73458 9101
rect -74274 9068 -74258 9085
rect -75132 9051 -74724 9068
rect -76324 9004 -74724 9051
rect -74666 9051 -74258 9068
rect -73474 9068 -73458 9085
rect -72616 9085 -71800 9101
rect -72616 9068 -72600 9085
rect -73474 9051 -73066 9068
rect -74666 9004 -73066 9051
rect -73008 9051 -72600 9068
rect -71816 9068 -71800 9085
rect -70958 9085 -70142 9101
rect -70958 9068 -70942 9085
rect -71816 9051 -71408 9068
rect -73008 9004 -71408 9051
rect -71350 9051 -70942 9068
rect -70158 9068 -70142 9085
rect -69300 9085 -68484 9101
rect -69300 9068 -69284 9085
rect -70158 9051 -69750 9068
rect -71350 9004 -69750 9051
rect -69692 9051 -69284 9068
rect -68500 9068 -68484 9085
rect -67642 9085 -66826 9101
rect -67642 9068 -67626 9085
rect -68500 9051 -68092 9068
rect -69692 9004 -68092 9051
rect -68034 9051 -67626 9068
rect -66842 9068 -66826 9085
rect -65984 9085 -65168 9101
rect -65984 9068 -65968 9085
rect -66842 9051 -66434 9068
rect -68034 9004 -66434 9051
rect -66376 9051 -65968 9068
rect -65184 9068 -65168 9085
rect -64326 9085 -63510 9101
rect -64326 9068 -64310 9085
rect -65184 9051 -64776 9068
rect -66376 9004 -64776 9051
rect -64718 9051 -64310 9068
rect -63526 9068 -63510 9085
rect -62668 9085 -61852 9101
rect -62668 9068 -62652 9085
rect -63526 9051 -63118 9068
rect -64718 9004 -63118 9051
rect -63060 9051 -62652 9068
rect -61868 9068 -61852 9085
rect -61010 9085 -60194 9101
rect -61010 9068 -60994 9085
rect -61868 9051 -61460 9068
rect -63060 9004 -61460 9051
rect -61402 9051 -60994 9068
rect -60210 9068 -60194 9085
rect -59352 9085 -58536 9101
rect -59352 9068 -59336 9085
rect -60210 9051 -59802 9068
rect -61402 9004 -59802 9051
rect -59744 9051 -59336 9068
rect -58552 9068 -58536 9085
rect -57694 9085 -56878 9101
rect -57694 9068 -57678 9085
rect -58552 9051 -58144 9068
rect -59744 9004 -58144 9051
rect -58086 9051 -57678 9068
rect -56894 9068 -56878 9085
rect -56036 9085 -55220 9101
rect -56036 9068 -56020 9085
rect -56894 9051 -56486 9068
rect -58086 9004 -56486 9051
rect -56428 9051 -56020 9068
rect -55236 9068 -55220 9085
rect -54378 9085 -53562 9101
rect -54378 9068 -54362 9085
rect -55236 9051 -54828 9068
rect -56428 9004 -54828 9051
rect -54770 9051 -54362 9068
rect -53578 9068 -53562 9085
rect -52720 9085 -51904 9101
rect -52720 9068 -52704 9085
rect -53578 9051 -53170 9068
rect -54770 9004 -53170 9051
rect -53112 9051 -52704 9068
rect -51920 9068 -51904 9085
rect -51062 9085 -50246 9101
rect -51062 9068 -51046 9085
rect -51920 9051 -51512 9068
rect -53112 9004 -51512 9051
rect -51454 9051 -51046 9068
rect -50262 9068 -50246 9085
rect -49404 9085 -48588 9101
rect -49404 9068 -49388 9085
rect -50262 9051 -49854 9068
rect -51454 9004 -49854 9051
rect -49796 9051 -49388 9068
rect -48604 9068 -48588 9085
rect -47746 9085 -46930 9101
rect -47746 9068 -47730 9085
rect -48604 9051 -48196 9068
rect -49796 9004 -48196 9051
rect -48138 9051 -47730 9068
rect -46946 9068 -46930 9085
rect -46088 9085 -45272 9101
rect -46088 9068 -46072 9085
rect -46946 9051 -46538 9068
rect -48138 9004 -46538 9051
rect -46480 9051 -46072 9068
rect -45288 9068 -45272 9085
rect -44430 9085 -43614 9101
rect -44430 9068 -44414 9085
rect -45288 9051 -44880 9068
rect -46480 9004 -44880 9051
rect -44822 9051 -44414 9068
rect -43630 9068 -43614 9085
rect -42772 9085 -41956 9101
rect -42772 9068 -42756 9085
rect -43630 9051 -43222 9068
rect -44822 9004 -43222 9051
rect -43164 9051 -42756 9068
rect -41972 9068 -41956 9085
rect -41114 9085 -40298 9101
rect -41114 9068 -41098 9085
rect -41972 9051 -41564 9068
rect -43164 9004 -41564 9051
rect -41506 9051 -41098 9068
rect -40314 9068 -40298 9085
rect -39456 9085 -38640 9101
rect -39456 9068 -39440 9085
rect -40314 9051 -39906 9068
rect -41506 9004 -39906 9051
rect -39848 9051 -39440 9068
rect -38656 9068 -38640 9085
rect -37798 9085 -36982 9101
rect -37798 9068 -37782 9085
rect -38656 9051 -38248 9068
rect -39848 9004 -38248 9051
rect -38190 9051 -37782 9068
rect -36998 9068 -36982 9085
rect -36140 9085 -35324 9101
rect -36140 9068 -36124 9085
rect -36998 9051 -36590 9068
rect -38190 9004 -36590 9051
rect -36532 9051 -36124 9068
rect -35340 9068 -35324 9085
rect -34482 9085 -33666 9101
rect -34482 9068 -34466 9085
rect -35340 9051 -34932 9068
rect -36532 9004 -34932 9051
rect -34874 9051 -34466 9068
rect -33682 9068 -33666 9085
rect -32824 9085 -32008 9101
rect -32824 9068 -32808 9085
rect -33682 9051 -33274 9068
rect -34874 9004 -33274 9051
rect -33216 9051 -32808 9068
rect -32024 9068 -32008 9085
rect -31166 9085 -30350 9101
rect -31166 9068 -31150 9085
rect -32024 9051 -31616 9068
rect -33216 9004 -31616 9051
rect -31558 9051 -31150 9068
rect -30366 9068 -30350 9085
rect -29508 9085 -28692 9101
rect -29508 9068 -29492 9085
rect -30366 9051 -29958 9068
rect -31558 9004 -29958 9051
rect -29900 9051 -29492 9068
rect -28708 9068 -28692 9085
rect -28708 9051 -28300 9068
rect -29900 9004 -28300 9051
rect -94562 7557 -92962 7604
rect -94562 7540 -94154 7557
rect -94170 7523 -94154 7540
rect -93370 7540 -92962 7557
rect -92904 7557 -91304 7604
rect -92904 7540 -92496 7557
rect -93370 7523 -93354 7540
rect -94170 7507 -93354 7523
rect -92512 7523 -92496 7540
rect -91712 7540 -91304 7557
rect -91246 7557 -89646 7604
rect -91246 7540 -90838 7557
rect -91712 7523 -91696 7540
rect -92512 7507 -91696 7523
rect -90854 7523 -90838 7540
rect -90054 7540 -89646 7557
rect -89588 7557 -87988 7604
rect -89588 7540 -89180 7557
rect -90054 7523 -90038 7540
rect -90854 7507 -90038 7523
rect -89196 7523 -89180 7540
rect -88396 7540 -87988 7557
rect -87930 7557 -86330 7604
rect -87930 7540 -87522 7557
rect -88396 7523 -88380 7540
rect -89196 7507 -88380 7523
rect -87538 7523 -87522 7540
rect -86738 7540 -86330 7557
rect -86272 7557 -84672 7604
rect -86272 7540 -85864 7557
rect -86738 7523 -86722 7540
rect -87538 7507 -86722 7523
rect -85880 7523 -85864 7540
rect -85080 7540 -84672 7557
rect -84614 7557 -83014 7604
rect -84614 7540 -84206 7557
rect -85080 7523 -85064 7540
rect -85880 7507 -85064 7523
rect -84222 7523 -84206 7540
rect -83422 7540 -83014 7557
rect -82956 7557 -81356 7604
rect -82956 7540 -82548 7557
rect -83422 7523 -83406 7540
rect -84222 7507 -83406 7523
rect -82564 7523 -82548 7540
rect -81764 7540 -81356 7557
rect -81298 7557 -79698 7604
rect -81298 7540 -80890 7557
rect -81764 7523 -81748 7540
rect -82564 7507 -81748 7523
rect -80906 7523 -80890 7540
rect -80106 7540 -79698 7557
rect -79640 7557 -78040 7604
rect -79640 7540 -79232 7557
rect -80106 7523 -80090 7540
rect -80906 7507 -80090 7523
rect -79248 7523 -79232 7540
rect -78448 7540 -78040 7557
rect -77982 7557 -76382 7604
rect -77982 7540 -77574 7557
rect -78448 7523 -78432 7540
rect -79248 7507 -78432 7523
rect -77590 7523 -77574 7540
rect -76790 7540 -76382 7557
rect -76324 7557 -74724 7604
rect -76324 7540 -75916 7557
rect -76790 7523 -76774 7540
rect -77590 7507 -76774 7523
rect -75932 7523 -75916 7540
rect -75132 7540 -74724 7557
rect -74666 7557 -73066 7604
rect -74666 7540 -74258 7557
rect -75132 7523 -75116 7540
rect -75932 7507 -75116 7523
rect -74274 7523 -74258 7540
rect -73474 7540 -73066 7557
rect -73008 7557 -71408 7604
rect -73008 7540 -72600 7557
rect -73474 7523 -73458 7540
rect -74274 7507 -73458 7523
rect -72616 7523 -72600 7540
rect -71816 7540 -71408 7557
rect -71350 7557 -69750 7604
rect -71350 7540 -70942 7557
rect -71816 7523 -71800 7540
rect -72616 7507 -71800 7523
rect -70958 7523 -70942 7540
rect -70158 7540 -69750 7557
rect -69692 7557 -68092 7604
rect -69692 7540 -69284 7557
rect -70158 7523 -70142 7540
rect -70958 7507 -70142 7523
rect -69300 7523 -69284 7540
rect -68500 7540 -68092 7557
rect -68034 7557 -66434 7604
rect -68034 7540 -67626 7557
rect -68500 7523 -68484 7540
rect -69300 7507 -68484 7523
rect -67642 7523 -67626 7540
rect -66842 7540 -66434 7557
rect -66376 7557 -64776 7604
rect -66376 7540 -65968 7557
rect -66842 7523 -66826 7540
rect -67642 7507 -66826 7523
rect -65984 7523 -65968 7540
rect -65184 7540 -64776 7557
rect -64718 7557 -63118 7604
rect -64718 7540 -64310 7557
rect -65184 7523 -65168 7540
rect -65984 7507 -65168 7523
rect -64326 7523 -64310 7540
rect -63526 7540 -63118 7557
rect -63060 7557 -61460 7604
rect -63060 7540 -62652 7557
rect -63526 7523 -63510 7540
rect -64326 7507 -63510 7523
rect -62668 7523 -62652 7540
rect -61868 7540 -61460 7557
rect -61402 7557 -59802 7604
rect -61402 7540 -60994 7557
rect -61868 7523 -61852 7540
rect -62668 7507 -61852 7523
rect -61010 7523 -60994 7540
rect -60210 7540 -59802 7557
rect -59744 7557 -58144 7604
rect -59744 7540 -59336 7557
rect -60210 7523 -60194 7540
rect -61010 7507 -60194 7523
rect -59352 7523 -59336 7540
rect -58552 7540 -58144 7557
rect -58086 7557 -56486 7604
rect -58086 7540 -57678 7557
rect -58552 7523 -58536 7540
rect -59352 7507 -58536 7523
rect -57694 7523 -57678 7540
rect -56894 7540 -56486 7557
rect -56428 7557 -54828 7604
rect -56428 7540 -56020 7557
rect -56894 7523 -56878 7540
rect -57694 7507 -56878 7523
rect -56036 7523 -56020 7540
rect -55236 7540 -54828 7557
rect -54770 7557 -53170 7604
rect -54770 7540 -54362 7557
rect -55236 7523 -55220 7540
rect -56036 7507 -55220 7523
rect -54378 7523 -54362 7540
rect -53578 7540 -53170 7557
rect -53112 7557 -51512 7604
rect -53112 7540 -52704 7557
rect -53578 7523 -53562 7540
rect -54378 7507 -53562 7523
rect -52720 7523 -52704 7540
rect -51920 7540 -51512 7557
rect -51454 7557 -49854 7604
rect -51454 7540 -51046 7557
rect -51920 7523 -51904 7540
rect -52720 7507 -51904 7523
rect -51062 7523 -51046 7540
rect -50262 7540 -49854 7557
rect -49796 7557 -48196 7604
rect -49796 7540 -49388 7557
rect -50262 7523 -50246 7540
rect -51062 7507 -50246 7523
rect -49404 7523 -49388 7540
rect -48604 7540 -48196 7557
rect -48138 7557 -46538 7604
rect -48138 7540 -47730 7557
rect -48604 7523 -48588 7540
rect -49404 7507 -48588 7523
rect -47746 7523 -47730 7540
rect -46946 7540 -46538 7557
rect -46480 7557 -44880 7604
rect -46480 7540 -46072 7557
rect -46946 7523 -46930 7540
rect -47746 7507 -46930 7523
rect -46088 7523 -46072 7540
rect -45288 7540 -44880 7557
rect -44822 7557 -43222 7604
rect -44822 7540 -44414 7557
rect -45288 7523 -45272 7540
rect -46088 7507 -45272 7523
rect -44430 7523 -44414 7540
rect -43630 7540 -43222 7557
rect -43164 7557 -41564 7604
rect -43164 7540 -42756 7557
rect -43630 7523 -43614 7540
rect -44430 7507 -43614 7523
rect -42772 7523 -42756 7540
rect -41972 7540 -41564 7557
rect -41506 7557 -39906 7604
rect -41506 7540 -41098 7557
rect -41972 7523 -41956 7540
rect -42772 7507 -41956 7523
rect -41114 7523 -41098 7540
rect -40314 7540 -39906 7557
rect -39848 7557 -38248 7604
rect -39848 7540 -39440 7557
rect -40314 7523 -40298 7540
rect -41114 7507 -40298 7523
rect -39456 7523 -39440 7540
rect -38656 7540 -38248 7557
rect -38190 7557 -36590 7604
rect -38190 7540 -37782 7557
rect -38656 7523 -38640 7540
rect -39456 7507 -38640 7523
rect -37798 7523 -37782 7540
rect -36998 7540 -36590 7557
rect -36532 7557 -34932 7604
rect -36532 7540 -36124 7557
rect -36998 7523 -36982 7540
rect -37798 7507 -36982 7523
rect -36140 7523 -36124 7540
rect -35340 7540 -34932 7557
rect -34874 7557 -33274 7604
rect -34874 7540 -34466 7557
rect -35340 7523 -35324 7540
rect -36140 7507 -35324 7523
rect -34482 7523 -34466 7540
rect -33682 7540 -33274 7557
rect -33216 7557 -31616 7604
rect -33216 7540 -32808 7557
rect -33682 7523 -33666 7540
rect -34482 7507 -33666 7523
rect -32824 7523 -32808 7540
rect -32024 7540 -31616 7557
rect -31558 7557 -29958 7604
rect -31558 7540 -31150 7557
rect -32024 7523 -32008 7540
rect -32824 7507 -32008 7523
rect -31166 7523 -31150 7540
rect -30366 7540 -29958 7557
rect -29900 7557 -28300 7604
rect -29900 7540 -29492 7557
rect -30366 7523 -30350 7540
rect -31166 7507 -30350 7523
rect -29508 7523 -29492 7540
rect -28708 7540 -28300 7557
rect -28708 7523 -28692 7540
rect -29508 7507 -28692 7523
rect -94170 7449 -93354 7465
rect -94170 7432 -94154 7449
rect -94562 7415 -94154 7432
rect -93370 7432 -93354 7449
rect -92512 7449 -91696 7465
rect -92512 7432 -92496 7449
rect -93370 7415 -92962 7432
rect -94562 7368 -92962 7415
rect -92904 7415 -92496 7432
rect -91712 7432 -91696 7449
rect -90854 7449 -90038 7465
rect -90854 7432 -90838 7449
rect -91712 7415 -91304 7432
rect -92904 7368 -91304 7415
rect -91246 7415 -90838 7432
rect -90054 7432 -90038 7449
rect -89196 7449 -88380 7465
rect -89196 7432 -89180 7449
rect -90054 7415 -89646 7432
rect -91246 7368 -89646 7415
rect -89588 7415 -89180 7432
rect -88396 7432 -88380 7449
rect -87538 7449 -86722 7465
rect -87538 7432 -87522 7449
rect -88396 7415 -87988 7432
rect -89588 7368 -87988 7415
rect -87930 7415 -87522 7432
rect -86738 7432 -86722 7449
rect -85880 7449 -85064 7465
rect -85880 7432 -85864 7449
rect -86738 7415 -86330 7432
rect -87930 7368 -86330 7415
rect -86272 7415 -85864 7432
rect -85080 7432 -85064 7449
rect -84222 7449 -83406 7465
rect -84222 7432 -84206 7449
rect -85080 7415 -84672 7432
rect -86272 7368 -84672 7415
rect -84614 7415 -84206 7432
rect -83422 7432 -83406 7449
rect -82564 7449 -81748 7465
rect -82564 7432 -82548 7449
rect -83422 7415 -83014 7432
rect -84614 7368 -83014 7415
rect -82956 7415 -82548 7432
rect -81764 7432 -81748 7449
rect -80906 7449 -80090 7465
rect -80906 7432 -80890 7449
rect -81764 7415 -81356 7432
rect -82956 7368 -81356 7415
rect -81298 7415 -80890 7432
rect -80106 7432 -80090 7449
rect -79248 7449 -78432 7465
rect -79248 7432 -79232 7449
rect -80106 7415 -79698 7432
rect -81298 7368 -79698 7415
rect -79640 7415 -79232 7432
rect -78448 7432 -78432 7449
rect -77590 7449 -76774 7465
rect -77590 7432 -77574 7449
rect -78448 7415 -78040 7432
rect -79640 7368 -78040 7415
rect -77982 7415 -77574 7432
rect -76790 7432 -76774 7449
rect -75932 7449 -75116 7465
rect -75932 7432 -75916 7449
rect -76790 7415 -76382 7432
rect -77982 7368 -76382 7415
rect -76324 7415 -75916 7432
rect -75132 7432 -75116 7449
rect -74274 7449 -73458 7465
rect -74274 7432 -74258 7449
rect -75132 7415 -74724 7432
rect -76324 7368 -74724 7415
rect -74666 7415 -74258 7432
rect -73474 7432 -73458 7449
rect -72616 7449 -71800 7465
rect -72616 7432 -72600 7449
rect -73474 7415 -73066 7432
rect -74666 7368 -73066 7415
rect -73008 7415 -72600 7432
rect -71816 7432 -71800 7449
rect -70958 7449 -70142 7465
rect -70958 7432 -70942 7449
rect -71816 7415 -71408 7432
rect -73008 7368 -71408 7415
rect -71350 7415 -70942 7432
rect -70158 7432 -70142 7449
rect -69300 7449 -68484 7465
rect -69300 7432 -69284 7449
rect -70158 7415 -69750 7432
rect -71350 7368 -69750 7415
rect -69692 7415 -69284 7432
rect -68500 7432 -68484 7449
rect -67642 7449 -66826 7465
rect -67642 7432 -67626 7449
rect -68500 7415 -68092 7432
rect -69692 7368 -68092 7415
rect -68034 7415 -67626 7432
rect -66842 7432 -66826 7449
rect -65984 7449 -65168 7465
rect -65984 7432 -65968 7449
rect -66842 7415 -66434 7432
rect -68034 7368 -66434 7415
rect -66376 7415 -65968 7432
rect -65184 7432 -65168 7449
rect -64326 7449 -63510 7465
rect -64326 7432 -64310 7449
rect -65184 7415 -64776 7432
rect -66376 7368 -64776 7415
rect -64718 7415 -64310 7432
rect -63526 7432 -63510 7449
rect -62668 7449 -61852 7465
rect -62668 7432 -62652 7449
rect -63526 7415 -63118 7432
rect -64718 7368 -63118 7415
rect -63060 7415 -62652 7432
rect -61868 7432 -61852 7449
rect -61010 7449 -60194 7465
rect -61010 7432 -60994 7449
rect -61868 7415 -61460 7432
rect -63060 7368 -61460 7415
rect -61402 7415 -60994 7432
rect -60210 7432 -60194 7449
rect -59352 7449 -58536 7465
rect -59352 7432 -59336 7449
rect -60210 7415 -59802 7432
rect -61402 7368 -59802 7415
rect -59744 7415 -59336 7432
rect -58552 7432 -58536 7449
rect -57694 7449 -56878 7465
rect -57694 7432 -57678 7449
rect -58552 7415 -58144 7432
rect -59744 7368 -58144 7415
rect -58086 7415 -57678 7432
rect -56894 7432 -56878 7449
rect -56036 7449 -55220 7465
rect -56036 7432 -56020 7449
rect -56894 7415 -56486 7432
rect -58086 7368 -56486 7415
rect -56428 7415 -56020 7432
rect -55236 7432 -55220 7449
rect -54378 7449 -53562 7465
rect -54378 7432 -54362 7449
rect -55236 7415 -54828 7432
rect -56428 7368 -54828 7415
rect -54770 7415 -54362 7432
rect -53578 7432 -53562 7449
rect -52720 7449 -51904 7465
rect -52720 7432 -52704 7449
rect -53578 7415 -53170 7432
rect -54770 7368 -53170 7415
rect -53112 7415 -52704 7432
rect -51920 7432 -51904 7449
rect -51062 7449 -50246 7465
rect -51062 7432 -51046 7449
rect -51920 7415 -51512 7432
rect -53112 7368 -51512 7415
rect -51454 7415 -51046 7432
rect -50262 7432 -50246 7449
rect -49404 7449 -48588 7465
rect -49404 7432 -49388 7449
rect -50262 7415 -49854 7432
rect -51454 7368 -49854 7415
rect -49796 7415 -49388 7432
rect -48604 7432 -48588 7449
rect -47746 7449 -46930 7465
rect -47746 7432 -47730 7449
rect -48604 7415 -48196 7432
rect -49796 7368 -48196 7415
rect -48138 7415 -47730 7432
rect -46946 7432 -46930 7449
rect -46088 7449 -45272 7465
rect -46088 7432 -46072 7449
rect -46946 7415 -46538 7432
rect -48138 7368 -46538 7415
rect -46480 7415 -46072 7432
rect -45288 7432 -45272 7449
rect -44430 7449 -43614 7465
rect -44430 7432 -44414 7449
rect -45288 7415 -44880 7432
rect -46480 7368 -44880 7415
rect -44822 7415 -44414 7432
rect -43630 7432 -43614 7449
rect -42772 7449 -41956 7465
rect -42772 7432 -42756 7449
rect -43630 7415 -43222 7432
rect -44822 7368 -43222 7415
rect -43164 7415 -42756 7432
rect -41972 7432 -41956 7449
rect -41114 7449 -40298 7465
rect -41114 7432 -41098 7449
rect -41972 7415 -41564 7432
rect -43164 7368 -41564 7415
rect -41506 7415 -41098 7432
rect -40314 7432 -40298 7449
rect -39456 7449 -38640 7465
rect -39456 7432 -39440 7449
rect -40314 7415 -39906 7432
rect -41506 7368 -39906 7415
rect -39848 7415 -39440 7432
rect -38656 7432 -38640 7449
rect -37798 7449 -36982 7465
rect -37798 7432 -37782 7449
rect -38656 7415 -38248 7432
rect -39848 7368 -38248 7415
rect -38190 7415 -37782 7432
rect -36998 7432 -36982 7449
rect -36140 7449 -35324 7465
rect -36140 7432 -36124 7449
rect -36998 7415 -36590 7432
rect -38190 7368 -36590 7415
rect -36532 7415 -36124 7432
rect -35340 7432 -35324 7449
rect -34482 7449 -33666 7465
rect -34482 7432 -34466 7449
rect -35340 7415 -34932 7432
rect -36532 7368 -34932 7415
rect -34874 7415 -34466 7432
rect -33682 7432 -33666 7449
rect -32824 7449 -32008 7465
rect -32824 7432 -32808 7449
rect -33682 7415 -33274 7432
rect -34874 7368 -33274 7415
rect -33216 7415 -32808 7432
rect -32024 7432 -32008 7449
rect -31166 7449 -30350 7465
rect -31166 7432 -31150 7449
rect -32024 7415 -31616 7432
rect -33216 7368 -31616 7415
rect -31558 7415 -31150 7432
rect -30366 7432 -30350 7449
rect -29508 7449 -28692 7465
rect -29508 7432 -29492 7449
rect -30366 7415 -29958 7432
rect -31558 7368 -29958 7415
rect -29900 7415 -29492 7432
rect -28708 7432 -28692 7449
rect -28708 7415 -28300 7432
rect -29900 7368 -28300 7415
rect -94562 5921 -92962 5968
rect -94562 5904 -94154 5921
rect -94170 5887 -94154 5904
rect -93370 5904 -92962 5921
rect -92904 5921 -91304 5968
rect -92904 5904 -92496 5921
rect -93370 5887 -93354 5904
rect -94170 5871 -93354 5887
rect -92512 5887 -92496 5904
rect -91712 5904 -91304 5921
rect -91246 5921 -89646 5968
rect -91246 5904 -90838 5921
rect -91712 5887 -91696 5904
rect -92512 5871 -91696 5887
rect -90854 5887 -90838 5904
rect -90054 5904 -89646 5921
rect -89588 5921 -87988 5968
rect -89588 5904 -89180 5921
rect -90054 5887 -90038 5904
rect -90854 5871 -90038 5887
rect -89196 5887 -89180 5904
rect -88396 5904 -87988 5921
rect -87930 5921 -86330 5968
rect -87930 5904 -87522 5921
rect -88396 5887 -88380 5904
rect -89196 5871 -88380 5887
rect -87538 5887 -87522 5904
rect -86738 5904 -86330 5921
rect -86272 5921 -84672 5968
rect -86272 5904 -85864 5921
rect -86738 5887 -86722 5904
rect -87538 5871 -86722 5887
rect -85880 5887 -85864 5904
rect -85080 5904 -84672 5921
rect -84614 5921 -83014 5968
rect -84614 5904 -84206 5921
rect -85080 5887 -85064 5904
rect -85880 5871 -85064 5887
rect -84222 5887 -84206 5904
rect -83422 5904 -83014 5921
rect -82956 5921 -81356 5968
rect -82956 5904 -82548 5921
rect -83422 5887 -83406 5904
rect -84222 5871 -83406 5887
rect -82564 5887 -82548 5904
rect -81764 5904 -81356 5921
rect -81298 5921 -79698 5968
rect -81298 5904 -80890 5921
rect -81764 5887 -81748 5904
rect -82564 5871 -81748 5887
rect -80906 5887 -80890 5904
rect -80106 5904 -79698 5921
rect -79640 5921 -78040 5968
rect -79640 5904 -79232 5921
rect -80106 5887 -80090 5904
rect -80906 5871 -80090 5887
rect -79248 5887 -79232 5904
rect -78448 5904 -78040 5921
rect -77982 5921 -76382 5968
rect -77982 5904 -77574 5921
rect -78448 5887 -78432 5904
rect -79248 5871 -78432 5887
rect -77590 5887 -77574 5904
rect -76790 5904 -76382 5921
rect -76324 5921 -74724 5968
rect -76324 5904 -75916 5921
rect -76790 5887 -76774 5904
rect -77590 5871 -76774 5887
rect -75932 5887 -75916 5904
rect -75132 5904 -74724 5921
rect -74666 5921 -73066 5968
rect -74666 5904 -74258 5921
rect -75132 5887 -75116 5904
rect -75932 5871 -75116 5887
rect -74274 5887 -74258 5904
rect -73474 5904 -73066 5921
rect -73008 5921 -71408 5968
rect -73008 5904 -72600 5921
rect -73474 5887 -73458 5904
rect -74274 5871 -73458 5887
rect -72616 5887 -72600 5904
rect -71816 5904 -71408 5921
rect -71350 5921 -69750 5968
rect -71350 5904 -70942 5921
rect -71816 5887 -71800 5904
rect -72616 5871 -71800 5887
rect -70958 5887 -70942 5904
rect -70158 5904 -69750 5921
rect -69692 5921 -68092 5968
rect -69692 5904 -69284 5921
rect -70158 5887 -70142 5904
rect -70958 5871 -70142 5887
rect -69300 5887 -69284 5904
rect -68500 5904 -68092 5921
rect -68034 5921 -66434 5968
rect -68034 5904 -67626 5921
rect -68500 5887 -68484 5904
rect -69300 5871 -68484 5887
rect -67642 5887 -67626 5904
rect -66842 5904 -66434 5921
rect -66376 5921 -64776 5968
rect -66376 5904 -65968 5921
rect -66842 5887 -66826 5904
rect -67642 5871 -66826 5887
rect -65984 5887 -65968 5904
rect -65184 5904 -64776 5921
rect -64718 5921 -63118 5968
rect -64718 5904 -64310 5921
rect -65184 5887 -65168 5904
rect -65984 5871 -65168 5887
rect -64326 5887 -64310 5904
rect -63526 5904 -63118 5921
rect -63060 5921 -61460 5968
rect -63060 5904 -62652 5921
rect -63526 5887 -63510 5904
rect -64326 5871 -63510 5887
rect -62668 5887 -62652 5904
rect -61868 5904 -61460 5921
rect -61402 5921 -59802 5968
rect -61402 5904 -60994 5921
rect -61868 5887 -61852 5904
rect -62668 5871 -61852 5887
rect -61010 5887 -60994 5904
rect -60210 5904 -59802 5921
rect -59744 5921 -58144 5968
rect -59744 5904 -59336 5921
rect -60210 5887 -60194 5904
rect -61010 5871 -60194 5887
rect -59352 5887 -59336 5904
rect -58552 5904 -58144 5921
rect -58086 5921 -56486 5968
rect -58086 5904 -57678 5921
rect -58552 5887 -58536 5904
rect -59352 5871 -58536 5887
rect -57694 5887 -57678 5904
rect -56894 5904 -56486 5921
rect -56428 5921 -54828 5968
rect -56428 5904 -56020 5921
rect -56894 5887 -56878 5904
rect -57694 5871 -56878 5887
rect -56036 5887 -56020 5904
rect -55236 5904 -54828 5921
rect -54770 5921 -53170 5968
rect -54770 5904 -54362 5921
rect -55236 5887 -55220 5904
rect -56036 5871 -55220 5887
rect -54378 5887 -54362 5904
rect -53578 5904 -53170 5921
rect -53112 5921 -51512 5968
rect -53112 5904 -52704 5921
rect -53578 5887 -53562 5904
rect -54378 5871 -53562 5887
rect -52720 5887 -52704 5904
rect -51920 5904 -51512 5921
rect -51454 5921 -49854 5968
rect -51454 5904 -51046 5921
rect -51920 5887 -51904 5904
rect -52720 5871 -51904 5887
rect -51062 5887 -51046 5904
rect -50262 5904 -49854 5921
rect -49796 5921 -48196 5968
rect -49796 5904 -49388 5921
rect -50262 5887 -50246 5904
rect -51062 5871 -50246 5887
rect -49404 5887 -49388 5904
rect -48604 5904 -48196 5921
rect -48138 5921 -46538 5968
rect -48138 5904 -47730 5921
rect -48604 5887 -48588 5904
rect -49404 5871 -48588 5887
rect -47746 5887 -47730 5904
rect -46946 5904 -46538 5921
rect -46480 5921 -44880 5968
rect -46480 5904 -46072 5921
rect -46946 5887 -46930 5904
rect -47746 5871 -46930 5887
rect -46088 5887 -46072 5904
rect -45288 5904 -44880 5921
rect -44822 5921 -43222 5968
rect -44822 5904 -44414 5921
rect -45288 5887 -45272 5904
rect -46088 5871 -45272 5887
rect -44430 5887 -44414 5904
rect -43630 5904 -43222 5921
rect -43164 5921 -41564 5968
rect -43164 5904 -42756 5921
rect -43630 5887 -43614 5904
rect -44430 5871 -43614 5887
rect -42772 5887 -42756 5904
rect -41972 5904 -41564 5921
rect -41506 5921 -39906 5968
rect -41506 5904 -41098 5921
rect -41972 5887 -41956 5904
rect -42772 5871 -41956 5887
rect -41114 5887 -41098 5904
rect -40314 5904 -39906 5921
rect -39848 5921 -38248 5968
rect -39848 5904 -39440 5921
rect -40314 5887 -40298 5904
rect -41114 5871 -40298 5887
rect -39456 5887 -39440 5904
rect -38656 5904 -38248 5921
rect -38190 5921 -36590 5968
rect -38190 5904 -37782 5921
rect -38656 5887 -38640 5904
rect -39456 5871 -38640 5887
rect -37798 5887 -37782 5904
rect -36998 5904 -36590 5921
rect -36532 5921 -34932 5968
rect -36532 5904 -36124 5921
rect -36998 5887 -36982 5904
rect -37798 5871 -36982 5887
rect -36140 5887 -36124 5904
rect -35340 5904 -34932 5921
rect -34874 5921 -33274 5968
rect -34874 5904 -34466 5921
rect -35340 5887 -35324 5904
rect -36140 5871 -35324 5887
rect -34482 5887 -34466 5904
rect -33682 5904 -33274 5921
rect -33216 5921 -31616 5968
rect -33216 5904 -32808 5921
rect -33682 5887 -33666 5904
rect -34482 5871 -33666 5887
rect -32824 5887 -32808 5904
rect -32024 5904 -31616 5921
rect -31558 5921 -29958 5968
rect -31558 5904 -31150 5921
rect -32024 5887 -32008 5904
rect -32824 5871 -32008 5887
rect -31166 5887 -31150 5904
rect -30366 5904 -29958 5921
rect -29900 5921 -28300 5968
rect -29900 5904 -29492 5921
rect -30366 5887 -30350 5904
rect -31166 5871 -30350 5887
rect -29508 5887 -29492 5904
rect -28708 5904 -28300 5921
rect -28708 5887 -28692 5904
rect -29508 5871 -28692 5887
rect -94170 5813 -93354 5829
rect -94170 5796 -94154 5813
rect -94562 5779 -94154 5796
rect -93370 5796 -93354 5813
rect -92512 5813 -91696 5829
rect -92512 5796 -92496 5813
rect -93370 5779 -92962 5796
rect -94562 5732 -92962 5779
rect -92904 5779 -92496 5796
rect -91712 5796 -91696 5813
rect -90854 5813 -90038 5829
rect -90854 5796 -90838 5813
rect -91712 5779 -91304 5796
rect -92904 5732 -91304 5779
rect -91246 5779 -90838 5796
rect -90054 5796 -90038 5813
rect -89196 5813 -88380 5829
rect -89196 5796 -89180 5813
rect -90054 5779 -89646 5796
rect -91246 5732 -89646 5779
rect -89588 5779 -89180 5796
rect -88396 5796 -88380 5813
rect -87538 5813 -86722 5829
rect -87538 5796 -87522 5813
rect -88396 5779 -87988 5796
rect -89588 5732 -87988 5779
rect -87930 5779 -87522 5796
rect -86738 5796 -86722 5813
rect -85880 5813 -85064 5829
rect -85880 5796 -85864 5813
rect -86738 5779 -86330 5796
rect -87930 5732 -86330 5779
rect -86272 5779 -85864 5796
rect -85080 5796 -85064 5813
rect -84222 5813 -83406 5829
rect -84222 5796 -84206 5813
rect -85080 5779 -84672 5796
rect -86272 5732 -84672 5779
rect -84614 5779 -84206 5796
rect -83422 5796 -83406 5813
rect -82564 5813 -81748 5829
rect -82564 5796 -82548 5813
rect -83422 5779 -83014 5796
rect -84614 5732 -83014 5779
rect -82956 5779 -82548 5796
rect -81764 5796 -81748 5813
rect -80906 5813 -80090 5829
rect -80906 5796 -80890 5813
rect -81764 5779 -81356 5796
rect -82956 5732 -81356 5779
rect -81298 5779 -80890 5796
rect -80106 5796 -80090 5813
rect -79248 5813 -78432 5829
rect -79248 5796 -79232 5813
rect -80106 5779 -79698 5796
rect -81298 5732 -79698 5779
rect -79640 5779 -79232 5796
rect -78448 5796 -78432 5813
rect -77590 5813 -76774 5829
rect -77590 5796 -77574 5813
rect -78448 5779 -78040 5796
rect -79640 5732 -78040 5779
rect -77982 5779 -77574 5796
rect -76790 5796 -76774 5813
rect -75932 5813 -75116 5829
rect -75932 5796 -75916 5813
rect -76790 5779 -76382 5796
rect -77982 5732 -76382 5779
rect -76324 5779 -75916 5796
rect -75132 5796 -75116 5813
rect -74274 5813 -73458 5829
rect -74274 5796 -74258 5813
rect -75132 5779 -74724 5796
rect -76324 5732 -74724 5779
rect -74666 5779 -74258 5796
rect -73474 5796 -73458 5813
rect -72616 5813 -71800 5829
rect -72616 5796 -72600 5813
rect -73474 5779 -73066 5796
rect -74666 5732 -73066 5779
rect -73008 5779 -72600 5796
rect -71816 5796 -71800 5813
rect -70958 5813 -70142 5829
rect -70958 5796 -70942 5813
rect -71816 5779 -71408 5796
rect -73008 5732 -71408 5779
rect -71350 5779 -70942 5796
rect -70158 5796 -70142 5813
rect -69300 5813 -68484 5829
rect -69300 5796 -69284 5813
rect -70158 5779 -69750 5796
rect -71350 5732 -69750 5779
rect -69692 5779 -69284 5796
rect -68500 5796 -68484 5813
rect -67642 5813 -66826 5829
rect -67642 5796 -67626 5813
rect -68500 5779 -68092 5796
rect -69692 5732 -68092 5779
rect -68034 5779 -67626 5796
rect -66842 5796 -66826 5813
rect -65984 5813 -65168 5829
rect -65984 5796 -65968 5813
rect -66842 5779 -66434 5796
rect -68034 5732 -66434 5779
rect -66376 5779 -65968 5796
rect -65184 5796 -65168 5813
rect -64326 5813 -63510 5829
rect -64326 5796 -64310 5813
rect -65184 5779 -64776 5796
rect -66376 5732 -64776 5779
rect -64718 5779 -64310 5796
rect -63526 5796 -63510 5813
rect -62668 5813 -61852 5829
rect -62668 5796 -62652 5813
rect -63526 5779 -63118 5796
rect -64718 5732 -63118 5779
rect -63060 5779 -62652 5796
rect -61868 5796 -61852 5813
rect -61010 5813 -60194 5829
rect -61010 5796 -60994 5813
rect -61868 5779 -61460 5796
rect -63060 5732 -61460 5779
rect -61402 5779 -60994 5796
rect -60210 5796 -60194 5813
rect -59352 5813 -58536 5829
rect -59352 5796 -59336 5813
rect -60210 5779 -59802 5796
rect -61402 5732 -59802 5779
rect -59744 5779 -59336 5796
rect -58552 5796 -58536 5813
rect -57694 5813 -56878 5829
rect -57694 5796 -57678 5813
rect -58552 5779 -58144 5796
rect -59744 5732 -58144 5779
rect -58086 5779 -57678 5796
rect -56894 5796 -56878 5813
rect -56036 5813 -55220 5829
rect -56036 5796 -56020 5813
rect -56894 5779 -56486 5796
rect -58086 5732 -56486 5779
rect -56428 5779 -56020 5796
rect -55236 5796 -55220 5813
rect -54378 5813 -53562 5829
rect -54378 5796 -54362 5813
rect -55236 5779 -54828 5796
rect -56428 5732 -54828 5779
rect -54770 5779 -54362 5796
rect -53578 5796 -53562 5813
rect -52720 5813 -51904 5829
rect -52720 5796 -52704 5813
rect -53578 5779 -53170 5796
rect -54770 5732 -53170 5779
rect -53112 5779 -52704 5796
rect -51920 5796 -51904 5813
rect -51062 5813 -50246 5829
rect -51062 5796 -51046 5813
rect -51920 5779 -51512 5796
rect -53112 5732 -51512 5779
rect -51454 5779 -51046 5796
rect -50262 5796 -50246 5813
rect -49404 5813 -48588 5829
rect -49404 5796 -49388 5813
rect -50262 5779 -49854 5796
rect -51454 5732 -49854 5779
rect -49796 5779 -49388 5796
rect -48604 5796 -48588 5813
rect -47746 5813 -46930 5829
rect -47746 5796 -47730 5813
rect -48604 5779 -48196 5796
rect -49796 5732 -48196 5779
rect -48138 5779 -47730 5796
rect -46946 5796 -46930 5813
rect -46088 5813 -45272 5829
rect -46088 5796 -46072 5813
rect -46946 5779 -46538 5796
rect -48138 5732 -46538 5779
rect -46480 5779 -46072 5796
rect -45288 5796 -45272 5813
rect -44430 5813 -43614 5829
rect -44430 5796 -44414 5813
rect -45288 5779 -44880 5796
rect -46480 5732 -44880 5779
rect -44822 5779 -44414 5796
rect -43630 5796 -43614 5813
rect -42772 5813 -41956 5829
rect -42772 5796 -42756 5813
rect -43630 5779 -43222 5796
rect -44822 5732 -43222 5779
rect -43164 5779 -42756 5796
rect -41972 5796 -41956 5813
rect -41114 5813 -40298 5829
rect -41114 5796 -41098 5813
rect -41972 5779 -41564 5796
rect -43164 5732 -41564 5779
rect -41506 5779 -41098 5796
rect -40314 5796 -40298 5813
rect -39456 5813 -38640 5829
rect -39456 5796 -39440 5813
rect -40314 5779 -39906 5796
rect -41506 5732 -39906 5779
rect -39848 5779 -39440 5796
rect -38656 5796 -38640 5813
rect -37798 5813 -36982 5829
rect -37798 5796 -37782 5813
rect -38656 5779 -38248 5796
rect -39848 5732 -38248 5779
rect -38190 5779 -37782 5796
rect -36998 5796 -36982 5813
rect -36140 5813 -35324 5829
rect -36140 5796 -36124 5813
rect -36998 5779 -36590 5796
rect -38190 5732 -36590 5779
rect -36532 5779 -36124 5796
rect -35340 5796 -35324 5813
rect -34482 5813 -33666 5829
rect -34482 5796 -34466 5813
rect -35340 5779 -34932 5796
rect -36532 5732 -34932 5779
rect -34874 5779 -34466 5796
rect -33682 5796 -33666 5813
rect -32824 5813 -32008 5829
rect -32824 5796 -32808 5813
rect -33682 5779 -33274 5796
rect -34874 5732 -33274 5779
rect -33216 5779 -32808 5796
rect -32024 5796 -32008 5813
rect -31166 5813 -30350 5829
rect -31166 5796 -31150 5813
rect -32024 5779 -31616 5796
rect -33216 5732 -31616 5779
rect -31558 5779 -31150 5796
rect -30366 5796 -30350 5813
rect -29508 5813 -28692 5829
rect -29508 5796 -29492 5813
rect -30366 5779 -29958 5796
rect -31558 5732 -29958 5779
rect -29900 5779 -29492 5796
rect -28708 5796 -28692 5813
rect -28708 5779 -28300 5796
rect -29900 5732 -28300 5779
rect 2708 5997 2824 6013
rect 2708 5980 2724 5997
rect 2666 5963 2724 5980
rect 2808 5980 2824 5997
rect 3364 6005 3480 6021
rect 3364 5988 3380 6005
rect 2808 5963 2866 5980
rect 2666 5916 2866 5963
rect 3322 5971 3380 5988
rect 3464 5988 3480 6005
rect 3622 6005 3738 6021
rect 3622 5988 3638 6005
rect 3464 5971 3522 5988
rect 3322 5924 3522 5971
rect 3580 5971 3638 5988
rect 3722 5988 3738 6005
rect 4364 6005 4480 6021
rect 4364 5988 4380 6005
rect 3722 5971 3780 5988
rect 3580 5924 3780 5971
rect 4322 5971 4380 5988
rect 4464 5988 4480 6005
rect 4622 6005 4738 6021
rect 4622 5988 4638 6005
rect 4464 5971 4522 5988
rect 4322 5924 4522 5971
rect 4580 5971 4638 5988
rect 4722 5988 4738 6005
rect 5270 6009 5386 6025
rect 5270 5992 5286 6009
rect 4722 5971 4780 5988
rect 4580 5924 4780 5971
rect 5228 5975 5286 5992
rect 5370 5992 5386 6009
rect 5370 5975 5428 5992
rect 5228 5928 5428 5975
rect -94562 4285 -92962 4332
rect -94562 4268 -94154 4285
rect -94170 4251 -94154 4268
rect -93370 4268 -92962 4285
rect -92904 4285 -91304 4332
rect -92904 4268 -92496 4285
rect -93370 4251 -93354 4268
rect -94170 4235 -93354 4251
rect -92512 4251 -92496 4268
rect -91712 4268 -91304 4285
rect -91246 4285 -89646 4332
rect -91246 4268 -90838 4285
rect -91712 4251 -91696 4268
rect -92512 4235 -91696 4251
rect -90854 4251 -90838 4268
rect -90054 4268 -89646 4285
rect -89588 4285 -87988 4332
rect -89588 4268 -89180 4285
rect -90054 4251 -90038 4268
rect -90854 4235 -90038 4251
rect -89196 4251 -89180 4268
rect -88396 4268 -87988 4285
rect -87930 4285 -86330 4332
rect -87930 4268 -87522 4285
rect -88396 4251 -88380 4268
rect -89196 4235 -88380 4251
rect -87538 4251 -87522 4268
rect -86738 4268 -86330 4285
rect -86272 4285 -84672 4332
rect -86272 4268 -85864 4285
rect -86738 4251 -86722 4268
rect -87538 4235 -86722 4251
rect -85880 4251 -85864 4268
rect -85080 4268 -84672 4285
rect -84614 4285 -83014 4332
rect -84614 4268 -84206 4285
rect -85080 4251 -85064 4268
rect -85880 4235 -85064 4251
rect -84222 4251 -84206 4268
rect -83422 4268 -83014 4285
rect -82956 4285 -81356 4332
rect -82956 4268 -82548 4285
rect -83422 4251 -83406 4268
rect -84222 4235 -83406 4251
rect -82564 4251 -82548 4268
rect -81764 4268 -81356 4285
rect -81298 4285 -79698 4332
rect -81298 4268 -80890 4285
rect -81764 4251 -81748 4268
rect -82564 4235 -81748 4251
rect -80906 4251 -80890 4268
rect -80106 4268 -79698 4285
rect -79640 4285 -78040 4332
rect -79640 4268 -79232 4285
rect -80106 4251 -80090 4268
rect -80906 4235 -80090 4251
rect -79248 4251 -79232 4268
rect -78448 4268 -78040 4285
rect -77982 4285 -76382 4332
rect -77982 4268 -77574 4285
rect -78448 4251 -78432 4268
rect -79248 4235 -78432 4251
rect -77590 4251 -77574 4268
rect -76790 4268 -76382 4285
rect -76324 4285 -74724 4332
rect -76324 4268 -75916 4285
rect -76790 4251 -76774 4268
rect -77590 4235 -76774 4251
rect -75932 4251 -75916 4268
rect -75132 4268 -74724 4285
rect -74666 4285 -73066 4332
rect -74666 4268 -74258 4285
rect -75132 4251 -75116 4268
rect -75932 4235 -75116 4251
rect -74274 4251 -74258 4268
rect -73474 4268 -73066 4285
rect -73008 4285 -71408 4332
rect -73008 4268 -72600 4285
rect -73474 4251 -73458 4268
rect -74274 4235 -73458 4251
rect -72616 4251 -72600 4268
rect -71816 4268 -71408 4285
rect -71350 4285 -69750 4332
rect -71350 4268 -70942 4285
rect -71816 4251 -71800 4268
rect -72616 4235 -71800 4251
rect -70958 4251 -70942 4268
rect -70158 4268 -69750 4285
rect -69692 4285 -68092 4332
rect -69692 4268 -69284 4285
rect -70158 4251 -70142 4268
rect -70958 4235 -70142 4251
rect -69300 4251 -69284 4268
rect -68500 4268 -68092 4285
rect -68034 4285 -66434 4332
rect -68034 4268 -67626 4285
rect -68500 4251 -68484 4268
rect -69300 4235 -68484 4251
rect -67642 4251 -67626 4268
rect -66842 4268 -66434 4285
rect -66376 4285 -64776 4332
rect -66376 4268 -65968 4285
rect -66842 4251 -66826 4268
rect -67642 4235 -66826 4251
rect -65984 4251 -65968 4268
rect -65184 4268 -64776 4285
rect -64718 4285 -63118 4332
rect -64718 4268 -64310 4285
rect -65184 4251 -65168 4268
rect -65984 4235 -65168 4251
rect -64326 4251 -64310 4268
rect -63526 4268 -63118 4285
rect -63060 4285 -61460 4332
rect -63060 4268 -62652 4285
rect -63526 4251 -63510 4268
rect -64326 4235 -63510 4251
rect -62668 4251 -62652 4268
rect -61868 4268 -61460 4285
rect -61402 4285 -59802 4332
rect -61402 4268 -60994 4285
rect -61868 4251 -61852 4268
rect -62668 4235 -61852 4251
rect -61010 4251 -60994 4268
rect -60210 4268 -59802 4285
rect -59744 4285 -58144 4332
rect -59744 4268 -59336 4285
rect -60210 4251 -60194 4268
rect -61010 4235 -60194 4251
rect -59352 4251 -59336 4268
rect -58552 4268 -58144 4285
rect -58086 4285 -56486 4332
rect -58086 4268 -57678 4285
rect -58552 4251 -58536 4268
rect -59352 4235 -58536 4251
rect -57694 4251 -57678 4268
rect -56894 4268 -56486 4285
rect -56428 4285 -54828 4332
rect -56428 4268 -56020 4285
rect -56894 4251 -56878 4268
rect -57694 4235 -56878 4251
rect -56036 4251 -56020 4268
rect -55236 4268 -54828 4285
rect -54770 4285 -53170 4332
rect -54770 4268 -54362 4285
rect -55236 4251 -55220 4268
rect -56036 4235 -55220 4251
rect -54378 4251 -54362 4268
rect -53578 4268 -53170 4285
rect -53112 4285 -51512 4332
rect -53112 4268 -52704 4285
rect -53578 4251 -53562 4268
rect -54378 4235 -53562 4251
rect -52720 4251 -52704 4268
rect -51920 4268 -51512 4285
rect -51454 4285 -49854 4332
rect -51454 4268 -51046 4285
rect -51920 4251 -51904 4268
rect -52720 4235 -51904 4251
rect -51062 4251 -51046 4268
rect -50262 4268 -49854 4285
rect -49796 4285 -48196 4332
rect -49796 4268 -49388 4285
rect -50262 4251 -50246 4268
rect -51062 4235 -50246 4251
rect -49404 4251 -49388 4268
rect -48604 4268 -48196 4285
rect -48138 4285 -46538 4332
rect -48138 4268 -47730 4285
rect -48604 4251 -48588 4268
rect -49404 4235 -48588 4251
rect -47746 4251 -47730 4268
rect -46946 4268 -46538 4285
rect -46480 4285 -44880 4332
rect -46480 4268 -46072 4285
rect -46946 4251 -46930 4268
rect -47746 4235 -46930 4251
rect -46088 4251 -46072 4268
rect -45288 4268 -44880 4285
rect -44822 4285 -43222 4332
rect -44822 4268 -44414 4285
rect -45288 4251 -45272 4268
rect -46088 4235 -45272 4251
rect -44430 4251 -44414 4268
rect -43630 4268 -43222 4285
rect -43164 4285 -41564 4332
rect -43164 4268 -42756 4285
rect -43630 4251 -43614 4268
rect -44430 4235 -43614 4251
rect -42772 4251 -42756 4268
rect -41972 4268 -41564 4285
rect -41506 4285 -39906 4332
rect -41506 4268 -41098 4285
rect -41972 4251 -41956 4268
rect -42772 4235 -41956 4251
rect -41114 4251 -41098 4268
rect -40314 4268 -39906 4285
rect -39848 4285 -38248 4332
rect -39848 4268 -39440 4285
rect -40314 4251 -40298 4268
rect -41114 4235 -40298 4251
rect -39456 4251 -39440 4268
rect -38656 4268 -38248 4285
rect -38190 4285 -36590 4332
rect -38190 4268 -37782 4285
rect -38656 4251 -38640 4268
rect -39456 4235 -38640 4251
rect -37798 4251 -37782 4268
rect -36998 4268 -36590 4285
rect -36532 4285 -34932 4332
rect -36532 4268 -36124 4285
rect -36998 4251 -36982 4268
rect -37798 4235 -36982 4251
rect -36140 4251 -36124 4268
rect -35340 4268 -34932 4285
rect -34874 4285 -33274 4332
rect -34874 4268 -34466 4285
rect -35340 4251 -35324 4268
rect -36140 4235 -35324 4251
rect -34482 4251 -34466 4268
rect -33682 4268 -33274 4285
rect -33216 4285 -31616 4332
rect -33216 4268 -32808 4285
rect -33682 4251 -33666 4268
rect -34482 4235 -33666 4251
rect -32824 4251 -32808 4268
rect -32024 4268 -31616 4285
rect -31558 4285 -29958 4332
rect -31558 4268 -31150 4285
rect -32024 4251 -32008 4268
rect -32824 4235 -32008 4251
rect -31166 4251 -31150 4268
rect -30366 4268 -29958 4285
rect -29900 4285 -28300 4332
rect -29900 4268 -29492 4285
rect -30366 4251 -30350 4268
rect -31166 4235 -30350 4251
rect -29508 4251 -29492 4268
rect -28708 4268 -28300 4285
rect -28708 4251 -28692 4268
rect -29508 4235 -28692 4251
rect -61642 3971 -61576 3987
rect -61642 3937 -61626 3971
rect -61592 3937 -61576 3971
rect -61642 3921 -61576 3937
rect -61450 3971 -61384 3987
rect -61450 3937 -61434 3971
rect -61400 3937 -61384 3971
rect -61450 3921 -61384 3937
rect -61720 3890 -61690 3916
rect -61624 3890 -61594 3921
rect -61528 3890 -61498 3916
rect -61432 3890 -61402 3921
rect 1102 5119 1168 5135
rect 1102 5085 1118 5119
rect 1152 5085 1168 5119
rect 1102 5069 1168 5085
rect 1334 5117 1400 5133
rect 1334 5083 1350 5117
rect 1384 5083 1400 5117
rect 1120 5038 1150 5069
rect 1334 5067 1400 5083
rect 1562 5115 1628 5131
rect 1562 5081 1578 5115
rect 1612 5081 1628 5115
rect 1352 5036 1382 5067
rect 1562 5065 1628 5081
rect 1780 5117 1846 5133
rect 1780 5083 1796 5117
rect 1830 5083 1846 5117
rect 1780 5067 1846 5083
rect 1120 4607 1150 4638
rect 1580 5034 1610 5065
rect 1798 5036 1828 5067
rect 1102 4591 1168 4607
rect 1352 4605 1382 4636
rect 8644 5737 8760 5753
rect 8644 5720 8660 5737
rect 8602 5703 8660 5720
rect 8744 5720 8760 5737
rect 9123 5729 9239 5745
rect 8744 5703 8802 5720
rect 9123 5712 9139 5729
rect 8602 5656 8802 5703
rect 9081 5695 9139 5712
rect 9223 5712 9239 5729
rect 9381 5729 9497 5745
rect 9381 5712 9397 5729
rect 9223 5695 9281 5712
rect 6288 5137 6354 5153
rect 6288 5103 6304 5137
rect 6338 5103 6354 5137
rect 6288 5087 6354 5103
rect 6520 5135 6586 5151
rect 6520 5101 6536 5135
rect 6570 5101 6586 5135
rect 6306 5056 6336 5087
rect 6520 5085 6586 5101
rect 6748 5133 6814 5149
rect 6748 5099 6764 5133
rect 6798 5099 6814 5133
rect 2666 4890 2866 4916
rect 3322 4898 3522 4924
rect 3580 4898 3780 4924
rect 4322 4898 4522 4924
rect 4580 4898 4780 4924
rect 5228 4902 5428 4928
rect 6538 5054 6568 5085
rect 6748 5083 6814 5099
rect 6966 5135 7032 5151
rect 6966 5101 6982 5135
rect 7016 5101 7032 5135
rect 6966 5085 7032 5101
rect 1102 4557 1118 4591
rect 1152 4557 1168 4591
rect 1102 4541 1168 4557
rect 1334 4589 1400 4605
rect 1580 4603 1610 4634
rect 1798 4605 1828 4636
rect 6306 4625 6336 4656
rect 6766 5052 6796 5083
rect 6984 5054 7014 5085
rect 6288 4609 6354 4625
rect 6538 4623 6568 4654
rect 9081 5648 9281 5695
rect 9339 5695 9397 5712
rect 9481 5712 9497 5729
rect 9781 5731 9897 5747
rect 9781 5714 9797 5731
rect 9481 5695 9539 5712
rect 9339 5648 9539 5695
rect 9741 5697 9797 5714
rect 9881 5714 9897 5731
rect 10039 5731 10155 5747
rect 10039 5714 10055 5731
rect 9881 5697 9939 5714
rect 9741 5676 9939 5697
rect 9739 5650 9939 5676
rect 9997 5697 10055 5714
rect 10139 5714 10155 5731
rect 10139 5697 10197 5714
rect 9997 5650 10197 5697
rect 10438 5711 10554 5727
rect 10438 5694 10454 5711
rect 10396 5677 10454 5694
rect 10538 5694 10554 5711
rect 10538 5677 10596 5694
rect 1334 4555 1350 4589
rect 1384 4555 1400 4589
rect 1334 4539 1400 4555
rect 1562 4587 1628 4603
rect 1562 4553 1578 4587
rect 1612 4553 1628 4587
rect 1562 4537 1628 4553
rect 1780 4589 1846 4605
rect 1780 4555 1796 4589
rect 1830 4555 1846 4589
rect 6288 4575 6304 4609
rect 6338 4575 6354 4609
rect 6288 4559 6354 4575
rect 6520 4607 6586 4623
rect 6766 4621 6796 4652
rect 6984 4623 7014 4654
rect 8602 4630 8802 4656
rect 10396 5630 10596 5677
rect 6520 4573 6536 4607
rect 6570 4573 6586 4607
rect 6520 4557 6586 4573
rect 6748 4605 6814 4621
rect 6748 4571 6764 4605
rect 6798 4571 6814 4605
rect 6748 4555 6814 4571
rect 6966 4607 7032 4623
rect 9081 4622 9281 4648
rect 9339 4622 9539 4648
rect 9739 4624 9939 4650
rect 9997 4624 10197 4650
rect 13918 5609 14034 5625
rect 13918 5592 13934 5609
rect 13876 5575 13934 5592
rect 14018 5592 14034 5609
rect 15506 5621 15622 5637
rect 14018 5575 14076 5592
rect 13876 5528 14076 5575
rect 14362 5591 14578 5607
rect 14362 5574 14378 5591
rect 14270 5557 14378 5574
rect 14562 5574 14578 5591
rect 14934 5591 15150 5607
rect 15506 5604 15522 5621
rect 14934 5574 14950 5591
rect 14562 5557 14670 5574
rect 11464 5149 11530 5165
rect 11464 5115 11480 5149
rect 11514 5115 11530 5149
rect 11464 5099 11530 5115
rect 11696 5147 11762 5163
rect 11696 5113 11712 5147
rect 11746 5113 11762 5147
rect 11482 5068 11512 5099
rect 11696 5097 11762 5113
rect 11924 5145 11990 5161
rect 11924 5111 11940 5145
rect 11974 5111 11990 5145
rect 11714 5066 11744 5097
rect 11924 5095 11990 5111
rect 12142 5147 12208 5163
rect 12142 5113 12158 5147
rect 12192 5113 12208 5147
rect 12142 5097 12208 5113
rect 11482 4637 11512 4668
rect 11942 5064 11972 5095
rect 12160 5066 12190 5097
rect 6966 4573 6982 4607
rect 7016 4573 7032 4607
rect 10396 4604 10596 4630
rect 11464 4621 11530 4637
rect 11714 4635 11744 4666
rect 6966 4557 7032 4573
rect 11464 4587 11480 4621
rect 11514 4587 11530 4621
rect 11464 4571 11530 4587
rect 11696 4619 11762 4635
rect 11942 4633 11972 4664
rect 12160 4635 12190 4666
rect 11696 4585 11712 4619
rect 11746 4585 11762 4619
rect 11696 4569 11762 4585
rect 11924 4617 11990 4633
rect 11924 4583 11940 4617
rect 11974 4583 11990 4617
rect 11924 4567 11990 4583
rect 12142 4619 12208 4635
rect 12142 4585 12158 4619
rect 12192 4585 12208 4619
rect 12142 4569 12208 4585
rect 1780 4539 1846 4555
rect 14270 5510 14670 5557
rect 14842 5557 14950 5574
rect 15134 5574 15150 5591
rect 15464 5587 15522 5604
rect 15606 5604 15622 5621
rect 15606 5587 15664 5604
rect 15134 5557 15242 5574
rect 14842 5510 15242 5557
rect 15464 5540 15664 5587
rect 6312 4490 6378 4506
rect 1126 4472 1192 4488
rect 1126 4438 1142 4472
rect 1176 4438 1192 4472
rect 1126 4422 1192 4438
rect 1342 4474 1408 4490
rect 1342 4440 1358 4474
rect 1392 4440 1408 4474
rect 1342 4424 1408 4440
rect 1560 4474 1626 4490
rect 1560 4440 1576 4474
rect 1610 4440 1626 4474
rect 1560 4424 1626 4440
rect 1782 4472 1848 4488
rect 1782 4438 1798 4472
rect 1832 4438 1848 4472
rect 6312 4456 6328 4490
rect 6362 4456 6378 4490
rect 6312 4440 6378 4456
rect 6528 4492 6594 4508
rect 6528 4458 6544 4492
rect 6578 4458 6594 4492
rect 6528 4442 6594 4458
rect 6746 4492 6812 4508
rect 6746 4458 6762 4492
rect 6796 4458 6812 4492
rect 6746 4442 6812 4458
rect 6968 4490 7034 4506
rect 6968 4456 6984 4490
rect 7018 4456 7034 4490
rect 1144 4400 1174 4422
rect 1360 4402 1390 4424
rect 1578 4402 1608 4424
rect 1782 4422 1848 4438
rect 1800 4400 1830 4422
rect 6330 4418 6360 4440
rect 6546 4420 6576 4442
rect 6764 4420 6794 4442
rect 6968 4440 7034 4456
rect 11488 4502 11554 4518
rect 11488 4468 11504 4502
rect 11538 4468 11554 4502
rect 11488 4452 11554 4468
rect 11704 4504 11770 4520
rect 11704 4470 11720 4504
rect 11754 4470 11770 4504
rect 11704 4454 11770 4470
rect 11922 4504 11988 4520
rect 11922 4470 11938 4504
rect 11972 4470 11988 4504
rect 11922 4454 11988 4470
rect 12144 4502 12210 4518
rect 13876 4502 14076 4528
rect 17120 4941 17186 4957
rect 17120 4907 17136 4941
rect 17170 4907 17186 4941
rect 17120 4891 17186 4907
rect 17352 4939 17418 4955
rect 17352 4905 17368 4939
rect 17402 4905 17418 4939
rect 17138 4860 17168 4891
rect 17352 4889 17418 4905
rect 17580 4937 17646 4953
rect 17580 4903 17596 4937
rect 17630 4903 17646 4937
rect 15464 4514 15664 4540
rect 12144 4468 12160 4502
rect 12194 4468 12210 4502
rect 14270 4484 14670 4510
rect 14842 4484 15242 4510
rect 1144 4178 1174 4200
rect 1360 4180 1390 4202
rect 1578 4180 1608 4202
rect 6986 4418 7016 4440
rect 11506 4430 11536 4452
rect 11722 4432 11752 4454
rect 11940 4432 11970 4454
rect 12144 4452 12210 4468
rect 17370 4858 17400 4889
rect 17580 4887 17646 4903
rect 17798 4939 17864 4955
rect 17798 4905 17814 4939
rect 17848 4905 17864 4939
rect 17798 4889 17864 4905
rect 1126 4162 1192 4178
rect 1126 4128 1142 4162
rect 1176 4128 1192 4162
rect 1126 4112 1192 4128
rect 1342 4164 1408 4180
rect 1342 4130 1358 4164
rect 1392 4130 1408 4164
rect 1342 4114 1408 4130
rect 1560 4164 1626 4180
rect 1800 4178 1830 4200
rect 6330 4196 6360 4218
rect 6546 4198 6576 4220
rect 6764 4198 6794 4220
rect 12162 4430 12192 4452
rect 6312 4180 6378 4196
rect 1560 4130 1576 4164
rect 1610 4130 1626 4164
rect 1560 4114 1626 4130
rect 1782 4162 1848 4178
rect 1782 4128 1798 4162
rect 1832 4128 1848 4162
rect 6312 4146 6328 4180
rect 6362 4146 6378 4180
rect 6312 4130 6378 4146
rect 6528 4182 6594 4198
rect 6528 4148 6544 4182
rect 6578 4148 6594 4182
rect 6528 4132 6594 4148
rect 6746 4182 6812 4198
rect 6986 4196 7016 4218
rect 11506 4208 11536 4230
rect 11722 4210 11752 4232
rect 11940 4210 11970 4232
rect 17138 4429 17168 4460
rect 17598 4856 17628 4887
rect 17816 4858 17846 4889
rect 17120 4413 17186 4429
rect 17370 4427 17400 4458
rect 17120 4379 17136 4413
rect 17170 4379 17186 4413
rect 17120 4363 17186 4379
rect 17352 4411 17418 4427
rect 17598 4425 17628 4456
rect 17816 4427 17846 4458
rect 17352 4377 17368 4411
rect 17402 4377 17418 4411
rect 17352 4361 17418 4377
rect 17580 4409 17646 4425
rect 17580 4375 17596 4409
rect 17630 4375 17646 4409
rect 17580 4359 17646 4375
rect 17798 4411 17864 4427
rect 17798 4377 17814 4411
rect 17848 4377 17864 4411
rect 17798 4361 17864 4377
rect 17144 4294 17210 4310
rect 17144 4260 17160 4294
rect 17194 4260 17210 4294
rect 17144 4244 17210 4260
rect 17360 4296 17426 4312
rect 17360 4262 17376 4296
rect 17410 4262 17426 4296
rect 17360 4246 17426 4262
rect 17578 4296 17644 4312
rect 17578 4262 17594 4296
rect 17628 4262 17644 4296
rect 17578 4246 17644 4262
rect 17800 4294 17866 4310
rect 17800 4260 17816 4294
rect 17850 4260 17866 4294
rect 6746 4148 6762 4182
rect 6796 4148 6812 4182
rect 6746 4132 6812 4148
rect 6968 4180 7034 4196
rect 6968 4146 6984 4180
rect 7018 4146 7034 4180
rect 6968 4130 7034 4146
rect 11488 4192 11554 4208
rect 11488 4158 11504 4192
rect 11538 4158 11554 4192
rect 11488 4142 11554 4158
rect 11704 4194 11770 4210
rect 11704 4160 11720 4194
rect 11754 4160 11770 4194
rect 11704 4144 11770 4160
rect 11922 4194 11988 4210
rect 12162 4208 12192 4230
rect 17162 4222 17192 4244
rect 17378 4224 17408 4246
rect 17596 4224 17626 4246
rect 17800 4244 17866 4260
rect 11922 4160 11938 4194
rect 11972 4160 11988 4194
rect 11922 4144 11988 4160
rect 12144 4192 12210 4208
rect 12144 4158 12160 4192
rect 12194 4158 12210 4192
rect 12144 4142 12210 4158
rect 1782 4112 1848 4128
rect 17818 4222 17848 4244
rect 17162 4000 17192 4022
rect 17378 4002 17408 4024
rect 17596 4002 17626 4024
rect 17144 3984 17210 4000
rect 17144 3950 17160 3984
rect 17194 3950 17210 3984
rect 17144 3934 17210 3950
rect 17360 3986 17426 4002
rect 17360 3952 17376 3986
rect 17410 3952 17426 3986
rect 17360 3936 17426 3952
rect 17578 3986 17644 4002
rect 17818 4000 17848 4022
rect 17578 3952 17594 3986
rect 17628 3952 17644 3986
rect 17578 3936 17644 3952
rect 17800 3984 17866 4000
rect 17800 3950 17816 3984
rect 17850 3950 17866 3984
rect 17800 3934 17866 3950
rect -61720 3459 -61690 3490
rect -61624 3464 -61594 3490
rect -61528 3459 -61498 3490
rect -61432 3464 -61402 3490
rect -61738 3443 -61672 3459
rect -61738 3409 -61722 3443
rect -61688 3409 -61672 3443
rect -61738 3393 -61672 3409
rect -61546 3443 -61480 3459
rect -61546 3409 -61530 3443
rect -61496 3409 -61480 3443
rect -61546 3393 -61480 3409
rect -61690 3318 -61624 3334
rect -61690 3284 -61674 3318
rect -61640 3284 -61624 3318
rect -61768 3246 -61738 3272
rect -61690 3268 -61624 3284
rect -61498 3318 -61432 3334
rect -61498 3284 -61482 3318
rect -61448 3284 -61432 3318
rect -61672 3246 -61642 3268
rect -61576 3246 -61546 3272
rect -61498 3268 -61432 3284
rect 8882 3756 8982 3772
rect 8882 3739 8898 3756
rect 8832 3722 8898 3739
rect 8966 3739 8982 3756
rect 9140 3756 9240 3772
rect 9140 3739 9156 3756
rect 8966 3722 9032 3739
rect 8832 3684 9032 3722
rect 9090 3722 9156 3739
rect 9224 3739 9240 3756
rect 9398 3756 9498 3772
rect 9398 3739 9414 3756
rect 9224 3722 9290 3739
rect 9090 3684 9290 3722
rect 9348 3722 9414 3739
rect 9482 3739 9498 3756
rect 9896 3756 9996 3772
rect 9896 3739 9912 3756
rect 9482 3722 9548 3739
rect 9348 3684 9548 3722
rect 9846 3722 9912 3739
rect 9980 3739 9996 3756
rect 10154 3756 10254 3772
rect 10154 3739 10170 3756
rect 9980 3722 10046 3739
rect 9846 3684 10046 3722
rect 10104 3722 10170 3739
rect 10238 3739 10254 3756
rect 10412 3756 10512 3772
rect 10412 3739 10428 3756
rect 10238 3722 10304 3739
rect 10104 3684 10304 3722
rect 10362 3722 10428 3739
rect 10496 3739 10512 3756
rect 10496 3722 10562 3739
rect 10362 3684 10562 3722
rect -61480 3246 -61450 3268
rect 8832 3258 9032 3284
rect 9090 3258 9290 3284
rect 9348 3258 9548 3284
rect 9846 3258 10046 3284
rect 10104 3258 10304 3284
rect 10362 3258 10562 3284
rect 8882 3200 8982 3216
rect 8882 3183 8898 3200
rect 8832 3166 8898 3183
rect 8966 3183 8982 3200
rect 9140 3200 9240 3216
rect 9140 3183 9156 3200
rect 8966 3166 9032 3183
rect 8832 3128 9032 3166
rect 9090 3166 9156 3183
rect 9224 3183 9240 3200
rect 9398 3200 9498 3216
rect 9398 3183 9414 3200
rect 9224 3166 9290 3183
rect 9090 3128 9290 3166
rect 9348 3166 9414 3183
rect 9482 3183 9498 3200
rect 9896 3200 9996 3216
rect 9896 3183 9912 3200
rect 9482 3166 9548 3183
rect 9348 3128 9548 3166
rect 9846 3166 9912 3183
rect 9980 3183 9996 3200
rect 10154 3200 10254 3216
rect 10154 3183 10170 3200
rect 9980 3166 10046 3183
rect 9846 3128 10046 3166
rect 10104 3166 10170 3183
rect 10238 3183 10254 3200
rect 10412 3200 10512 3216
rect 10412 3183 10428 3200
rect 10238 3166 10304 3183
rect 10104 3128 10304 3166
rect 10362 3166 10428 3183
rect 10496 3183 10512 3200
rect 13406 3186 13522 3202
rect 10496 3166 10562 3183
rect 13406 3169 13422 3186
rect 10362 3128 10562 3166
rect 13364 3152 13422 3169
rect 13506 3169 13522 3186
rect 13506 3152 13564 3169
rect -61768 3024 -61738 3046
rect -61786 3008 -61720 3024
rect -61672 3020 -61642 3046
rect -61576 3024 -61546 3046
rect -61786 2974 -61770 3008
rect -61736 2974 -61720 3008
rect -61786 2958 -61720 2974
rect -61594 3008 -61528 3024
rect -61480 3020 -61450 3046
rect -61594 2974 -61578 3008
rect -61544 2974 -61528 3008
rect -61594 2958 -61528 2974
rect 13364 3114 13564 3152
rect 16004 3136 16120 3152
rect 16004 3119 16020 3136
rect 8832 2702 9032 2728
rect 9090 2702 9290 2728
rect 9348 2702 9548 2728
rect 9846 2702 10046 2728
rect 10104 2702 10304 2728
rect 10362 2702 10562 2728
rect 2714 2604 2830 2620
rect 2714 2587 2730 2604
rect 2672 2570 2730 2587
rect 2814 2587 2830 2604
rect 3340 2606 3756 2622
rect 3340 2589 3356 2606
rect 2814 2570 2872 2587
rect 2672 2532 2872 2570
rect 3148 2572 3356 2589
rect 3740 2589 3756 2606
rect 4312 2606 4728 2622
rect 4312 2589 4328 2606
rect 3740 2572 3948 2589
rect 3148 2534 3948 2572
rect 4120 2572 4328 2589
rect 4712 2589 4728 2606
rect 5248 2604 5364 2620
rect 4712 2572 4920 2589
rect 5248 2587 5264 2604
rect 4120 2534 4920 2572
rect 5206 2570 5264 2587
rect 5348 2587 5364 2604
rect 5348 2570 5406 2587
rect 5206 2532 5406 2570
rect 2672 2306 2872 2332
rect 3148 2308 3948 2334
rect 4120 2308 4920 2334
rect 5206 2306 5406 2332
rect 9245 1956 9461 1972
rect 9245 1939 9261 1956
rect 9153 1922 9261 1939
rect 9445 1939 9461 1956
rect 9840 1956 10056 1972
rect 9840 1939 9856 1956
rect 9445 1922 9553 1939
rect 9153 1884 9553 1922
rect 9748 1922 9856 1939
rect 10040 1939 10056 1956
rect 10040 1922 10148 1939
rect 9748 1884 10148 1922
rect 9153 1658 9553 1684
rect 9748 1658 10148 1684
rect 15962 3102 16020 3119
rect 16104 3119 16120 3136
rect 16104 3102 16162 3119
rect 13956 3052 14072 3068
rect 13956 3035 13972 3052
rect 13914 3018 13972 3035
rect 14056 3035 14072 3052
rect 14214 3052 14330 3068
rect 14214 3035 14230 3052
rect 14056 3018 14114 3035
rect 13914 2980 14114 3018
rect 14172 3018 14230 3035
rect 14314 3035 14330 3052
rect 14472 3052 14588 3068
rect 14472 3035 14488 3052
rect 14314 3018 14372 3035
rect 14172 2980 14372 3018
rect 14430 3018 14488 3035
rect 14572 3035 14588 3052
rect 14956 3052 15072 3068
rect 14956 3035 14972 3052
rect 14572 3018 14630 3035
rect 14430 2980 14630 3018
rect 14914 3018 14972 3035
rect 15056 3035 15072 3052
rect 15214 3052 15330 3068
rect 15214 3035 15230 3052
rect 15056 3018 15114 3035
rect 14914 2980 15114 3018
rect 15172 3018 15230 3035
rect 15314 3035 15330 3052
rect 15472 3052 15588 3068
rect 15962 3064 16162 3102
rect 15472 3035 15488 3052
rect 15314 3018 15372 3035
rect 15172 2980 15372 3018
rect 15430 3018 15488 3035
rect 15572 3035 15588 3052
rect 15572 3018 15630 3035
rect 15430 2980 15630 3018
rect 13914 2154 14114 2180
rect 14172 2154 14372 2180
rect 14430 2154 14630 2180
rect 14914 2154 15114 2180
rect 15172 2154 15372 2180
rect 15430 2154 15630 2180
rect 13956 2096 14072 2112
rect 13956 2079 13972 2096
rect 13914 2062 13972 2079
rect 14056 2079 14072 2096
rect 14214 2096 14330 2112
rect 14214 2079 14230 2096
rect 14056 2062 14114 2079
rect 13914 2024 14114 2062
rect 14172 2062 14230 2079
rect 14314 2079 14330 2096
rect 14472 2096 14588 2112
rect 14472 2079 14488 2096
rect 14314 2062 14372 2079
rect 14172 2024 14372 2062
rect 14430 2062 14488 2079
rect 14572 2079 14588 2096
rect 14956 2096 15072 2112
rect 14956 2079 14972 2096
rect 14572 2062 14630 2079
rect 14430 2024 14630 2062
rect 14914 2062 14972 2079
rect 15056 2079 15072 2096
rect 15214 2096 15330 2112
rect 15214 2079 15230 2096
rect 15056 2062 15114 2079
rect 14914 2024 15114 2062
rect 15172 2062 15230 2079
rect 15314 2079 15330 2096
rect 15472 2096 15588 2112
rect 15472 2079 15488 2096
rect 15314 2062 15372 2079
rect 15172 2024 15372 2062
rect 15430 2062 15488 2079
rect 15572 2079 15588 2096
rect 15572 2062 15630 2079
rect 15430 2024 15630 2062
rect 13914 1198 14114 1224
rect 14172 1198 14372 1224
rect 14430 1198 14630 1224
rect 14914 1198 15114 1224
rect 15172 1198 15372 1224
rect 15430 1198 15630 1224
rect 13956 1140 14072 1156
rect 13956 1123 13972 1140
rect 13914 1106 13972 1123
rect 14056 1123 14072 1140
rect 14214 1140 14330 1156
rect 14214 1123 14230 1140
rect 14056 1106 14114 1123
rect 13914 1068 14114 1106
rect 14172 1106 14230 1123
rect 14314 1123 14330 1140
rect 14472 1140 14588 1156
rect 14472 1123 14488 1140
rect 14314 1106 14372 1123
rect 14172 1068 14372 1106
rect 14430 1106 14488 1123
rect 14572 1123 14588 1140
rect 14956 1140 15072 1156
rect 14956 1123 14972 1140
rect 14572 1106 14630 1123
rect 14430 1068 14630 1106
rect 14914 1106 14972 1123
rect 15056 1123 15072 1140
rect 15214 1140 15330 1156
rect 15214 1123 15230 1140
rect 15056 1106 15114 1123
rect 14914 1068 15114 1106
rect 15172 1106 15230 1123
rect 15314 1123 15330 1140
rect 15472 1140 15588 1156
rect 15472 1123 15488 1140
rect 15314 1106 15372 1123
rect 15172 1068 15372 1106
rect 15430 1106 15488 1123
rect 15572 1123 15588 1140
rect 15572 1106 15630 1123
rect 15430 1068 15630 1106
rect 13364 288 13564 314
rect 13914 242 14114 268
rect 14172 242 14372 268
rect 14430 242 14630 268
rect 14914 242 15114 268
rect 15172 242 15372 268
rect 15430 242 15630 268
rect 26914 2887 26980 2903
rect 26914 2853 26930 2887
rect 26964 2853 26980 2887
rect 27526 2895 27592 2911
rect 26914 2837 26980 2853
rect 27136 2844 27166 2870
rect 27526 2861 27542 2895
rect 27576 2861 27592 2895
rect 28104 2891 28170 2907
rect 27526 2845 27592 2861
rect 27748 2852 27778 2878
rect 28104 2857 28120 2891
rect 28154 2857 28170 2891
rect 28678 2899 28744 2915
rect 26932 2806 26962 2837
rect 27544 2814 27574 2845
rect 27136 2477 27166 2508
rect 28104 2841 28170 2857
rect 28326 2848 28356 2874
rect 28678 2865 28694 2899
rect 28728 2865 28744 2899
rect 29256 2899 29322 2915
rect 28678 2849 28744 2865
rect 28900 2856 28930 2882
rect 29256 2865 29272 2899
rect 29306 2865 29322 2899
rect 29834 2899 29900 2915
rect 28122 2810 28152 2841
rect 27748 2485 27778 2516
rect 26932 2444 26962 2470
rect 27118 2461 27184 2477
rect 27118 2427 27134 2461
rect 27168 2427 27184 2461
rect 27544 2452 27574 2478
rect 27730 2469 27796 2485
rect 28696 2818 28726 2849
rect 28326 2481 28356 2512
rect 29256 2849 29322 2865
rect 29478 2856 29508 2882
rect 29834 2865 29850 2899
rect 29884 2865 29900 2899
rect 30416 2903 30482 2919
rect 29274 2818 29304 2849
rect 28900 2489 28930 2520
rect 27118 2411 27184 2427
rect 27730 2435 27746 2469
rect 27780 2435 27796 2469
rect 28122 2448 28152 2474
rect 28308 2465 28374 2481
rect 27730 2419 27796 2435
rect 28308 2431 28324 2465
rect 28358 2431 28374 2465
rect 28696 2456 28726 2482
rect 28882 2473 28948 2489
rect 29834 2849 29900 2865
rect 30056 2856 30086 2882
rect 30416 2869 30432 2903
rect 30466 2869 30482 2903
rect 30992 2899 31058 2915
rect 29852 2818 29882 2849
rect 29478 2489 29508 2520
rect 28308 2415 28374 2431
rect 28882 2439 28898 2473
rect 28932 2439 28948 2473
rect 29274 2456 29304 2482
rect 29460 2473 29526 2489
rect 30416 2853 30482 2869
rect 30638 2860 30668 2886
rect 30992 2865 31008 2899
rect 31042 2865 31058 2899
rect 31562 2895 31628 2911
rect 30434 2822 30464 2853
rect 30056 2489 30086 2520
rect 28882 2423 28948 2439
rect 29460 2439 29476 2473
rect 29510 2439 29526 2473
rect 29852 2456 29882 2482
rect 30038 2473 30104 2489
rect 30992 2849 31058 2865
rect 31214 2856 31244 2882
rect 31562 2861 31578 2895
rect 31612 2861 31628 2895
rect 31010 2818 31040 2849
rect 30638 2493 30668 2524
rect 29460 2423 29526 2439
rect 30038 2439 30054 2473
rect 30088 2439 30104 2473
rect 30434 2460 30464 2486
rect 30620 2477 30686 2493
rect 31562 2845 31628 2861
rect 31784 2852 31814 2878
rect 31580 2814 31610 2845
rect 31214 2489 31244 2520
rect 30038 2423 30104 2439
rect 30620 2443 30636 2477
rect 30670 2443 30686 2477
rect 31010 2456 31040 2482
rect 31196 2473 31262 2489
rect 31784 2485 31814 2516
rect 30620 2427 30686 2443
rect 31196 2439 31212 2473
rect 31246 2439 31262 2473
rect 31580 2452 31610 2478
rect 31766 2469 31832 2485
rect 31196 2423 31262 2439
rect 31766 2435 31782 2469
rect 31816 2435 31832 2469
rect 31766 2419 31832 2435
rect 27014 2280 27080 2296
rect 27014 2246 27030 2280
rect 27064 2246 27080 2280
rect 26936 2208 26966 2234
rect 27014 2230 27080 2246
rect 27626 2288 27692 2304
rect 27626 2254 27642 2288
rect 27676 2254 27692 2288
rect 27032 2208 27062 2230
rect 27548 2216 27578 2242
rect 27626 2238 27692 2254
rect 28204 2284 28270 2300
rect 28204 2250 28220 2284
rect 28254 2250 28270 2284
rect 27644 2216 27674 2238
rect 28126 2212 28156 2238
rect 28204 2234 28270 2250
rect 28778 2292 28844 2308
rect 28778 2258 28794 2292
rect 28828 2258 28844 2292
rect 28222 2212 28252 2234
rect 28700 2220 28730 2246
rect 28778 2242 28844 2258
rect 29356 2292 29422 2308
rect 29356 2258 29372 2292
rect 29406 2258 29422 2292
rect 28796 2220 28826 2242
rect 29278 2220 29308 2246
rect 29356 2242 29422 2258
rect 29934 2292 30000 2308
rect 29934 2258 29950 2292
rect 29984 2258 30000 2292
rect 29374 2220 29404 2242
rect 29856 2220 29886 2246
rect 29934 2242 30000 2258
rect 30516 2296 30582 2312
rect 30516 2262 30532 2296
rect 30566 2262 30582 2296
rect 29952 2220 29982 2242
rect 30438 2224 30468 2250
rect 30516 2246 30582 2262
rect 31092 2292 31158 2308
rect 31092 2258 31108 2292
rect 31142 2258 31158 2292
rect 30534 2224 30564 2246
rect 26936 2038 26966 2060
rect 26918 2022 26984 2038
rect 27032 2034 27062 2060
rect 27548 2046 27578 2068
rect 26918 1988 26934 2022
rect 26968 1988 26984 2022
rect 26918 1972 26984 1988
rect 27530 2030 27596 2046
rect 27644 2042 27674 2068
rect 31014 2220 31044 2246
rect 31092 2242 31158 2258
rect 31662 2288 31728 2304
rect 31662 2254 31678 2288
rect 31712 2254 31728 2288
rect 31110 2220 31140 2242
rect 28126 2042 28156 2064
rect 27530 1996 27546 2030
rect 27580 1996 27596 2030
rect 27530 1980 27596 1996
rect 28108 2026 28174 2042
rect 28222 2038 28252 2064
rect 28700 2050 28730 2072
rect 28108 1992 28124 2026
rect 28158 1992 28174 2026
rect 28108 1976 28174 1992
rect 28682 2034 28748 2050
rect 28796 2046 28826 2072
rect 29278 2050 29308 2072
rect 28682 2000 28698 2034
rect 28732 2000 28748 2034
rect 28682 1984 28748 2000
rect 29260 2034 29326 2050
rect 29374 2046 29404 2072
rect 29856 2050 29886 2072
rect 29260 2000 29276 2034
rect 29310 2000 29326 2034
rect 29260 1984 29326 2000
rect 29838 2034 29904 2050
rect 29952 2046 29982 2072
rect 30438 2054 30468 2076
rect 29838 2000 29854 2034
rect 29888 2000 29904 2034
rect 29838 1984 29904 2000
rect 30420 2038 30486 2054
rect 30534 2050 30564 2076
rect 31584 2216 31614 2242
rect 31662 2238 31728 2254
rect 31680 2216 31710 2238
rect 31014 2050 31044 2072
rect 30420 2004 30436 2038
rect 30470 2004 30486 2038
rect 30420 1988 30486 2004
rect 30996 2034 31062 2050
rect 31110 2046 31140 2072
rect 31584 2046 31614 2068
rect 30996 2000 31012 2034
rect 31046 2000 31062 2034
rect 30996 1984 31062 2000
rect 31566 2030 31632 2046
rect 31680 2042 31710 2068
rect 31566 1996 31582 2030
rect 31616 1996 31632 2030
rect 31566 1980 31632 1996
rect 28308 833 28374 849
rect 28308 799 28324 833
rect 28358 799 28374 833
rect 28710 831 28776 847
rect 28308 783 28374 799
rect 28526 790 28556 816
rect 28710 797 28726 831
rect 28760 797 28776 831
rect 28326 752 28356 783
rect 28710 781 28776 797
rect 28728 750 28758 781
rect 28526 423 28556 454
rect 28326 390 28356 416
rect 28508 407 28574 423
rect 29072 442 29138 458
rect 15962 238 16162 264
rect 28508 373 28524 407
rect 28558 373 28574 407
rect 28728 388 28758 414
rect 29072 408 29088 442
rect 29122 408 29138 442
rect 28508 357 28574 373
rect 28994 370 29024 396
rect 29072 392 29138 408
rect 29264 442 29330 458
rect 29264 408 29280 442
rect 29314 408 29330 442
rect 29090 370 29120 392
rect 29186 370 29216 396
rect 29264 392 29330 408
rect 29456 442 29522 458
rect 29456 408 29472 442
rect 29506 408 29522 442
rect 29282 370 29312 392
rect 29378 370 29408 396
rect 29456 392 29522 408
rect 29648 442 29714 458
rect 29648 408 29664 442
rect 29698 408 29714 442
rect 29474 370 29504 392
rect 29570 370 29600 396
rect 29648 392 29714 408
rect 29666 370 29696 392
rect 29762 370 29792 396
rect 28308 327 28374 343
rect 28308 293 28324 327
rect 28358 293 28374 327
rect 28708 327 28774 343
rect 28308 277 28374 293
rect 28526 284 28556 310
rect 28708 293 28724 327
rect 28758 293 28774 327
rect 28326 246 28356 277
rect 28708 277 28774 293
rect 28726 246 28756 277
rect 28526 -83 28556 -52
rect 28326 -116 28356 -90
rect 28508 -99 28574 -83
rect 28508 -133 28524 -99
rect 28558 -133 28574 -99
rect 28726 -116 28756 -90
rect 28508 -149 28574 -133
rect 28308 -181 28374 -165
rect 28308 -215 28324 -181
rect 28358 -215 28374 -181
rect 28708 -181 28774 -165
rect 28308 -231 28374 -215
rect 28526 -224 28556 -198
rect 28708 -215 28724 -181
rect 28758 -215 28774 -181
rect 28326 -262 28356 -231
rect 28708 -231 28774 -215
rect 28726 -262 28756 -231
rect 28526 -591 28556 -560
rect 28326 -624 28356 -598
rect 28508 -607 28574 -591
rect 28994 -300 29024 -278
rect 28976 -316 29042 -300
rect 29090 -304 29120 -278
rect 29186 -300 29216 -278
rect 28976 -350 28992 -316
rect 29026 -350 29042 -316
rect 28976 -366 29042 -350
rect 29168 -316 29234 -300
rect 29282 -304 29312 -278
rect 29378 -300 29408 -278
rect 29168 -350 29184 -316
rect 29218 -350 29234 -316
rect 29168 -366 29234 -350
rect 29360 -316 29426 -300
rect 29474 -304 29504 -278
rect 29570 -300 29600 -278
rect 29360 -350 29376 -316
rect 29410 -350 29426 -316
rect 29360 -366 29426 -350
rect 29552 -316 29618 -300
rect 29666 -304 29696 -278
rect 29762 -300 29792 -278
rect 29552 -350 29568 -316
rect 29602 -350 29618 -316
rect 29552 -366 29618 -350
rect 29744 -316 29810 -300
rect 29744 -350 29760 -316
rect 29794 -350 29810 -316
rect 29744 -366 29810 -350
rect 28508 -641 28524 -607
rect 28558 -641 28574 -607
rect 28726 -624 28756 -598
rect 28508 -657 28574 -641
rect 8813 -1028 8843 -1002
rect 8897 -1028 8927 -1002
rect 9164 -1022 9194 -996
rect 9256 -1022 9286 -996
rect 9355 -1022 9385 -996
rect 9495 -1022 9525 -996
rect 9592 -1022 9622 -996
rect 9789 -1022 9819 -996
rect 9888 -1022 9918 -996
rect 9974 -1022 10004 -996
rect 10058 -1022 10088 -996
rect 10166 -1022 10196 -996
rect 10250 -1022 10280 -996
rect 10414 -1022 10444 -996
rect 10633 -1022 10663 -996
rect 10730 -1022 10760 -996
rect 8813 -1171 8843 -1156
rect 8780 -1201 8843 -1171
rect 8780 -1254 8810 -1201
rect 8897 -1245 8927 -1156
rect 9164 -1193 9194 -1106
rect 9256 -1144 9286 -1106
rect 8756 -1270 8810 -1254
rect 8756 -1304 8766 -1270
rect 8800 -1304 8810 -1270
rect 8852 -1255 8927 -1245
rect 8852 -1289 8868 -1255
rect 8902 -1289 8927 -1255
rect 9065 -1209 9194 -1193
rect 9240 -1154 9306 -1144
rect 9240 -1188 9256 -1154
rect 9290 -1188 9306 -1154
rect 9240 -1198 9306 -1188
rect 9065 -1243 9075 -1209
rect 9109 -1223 9194 -1209
rect 9109 -1243 9182 -1223
rect 9355 -1240 9385 -1106
rect 9495 -1164 9525 -1106
rect 9495 -1180 9550 -1164
rect 9495 -1214 9505 -1180
rect 9539 -1214 9550 -1180
rect 9495 -1230 9550 -1214
rect 9065 -1259 9182 -1243
rect 8852 -1299 8927 -1289
rect 8756 -1320 8810 -1304
rect 8780 -1343 8810 -1320
rect 8780 -1373 8843 -1343
rect 8813 -1388 8843 -1373
rect 8897 -1388 8927 -1299
rect 9152 -1388 9182 -1259
rect 9247 -1270 9385 -1240
rect 9247 -1300 9278 -1270
rect 9224 -1316 9278 -1300
rect 9224 -1350 9234 -1316
rect 9268 -1350 9278 -1316
rect 9224 -1366 9278 -1350
rect 9320 -1322 9386 -1312
rect 9320 -1356 9336 -1322
rect 9370 -1356 9386 -1322
rect 9320 -1366 9386 -1356
rect 9247 -1400 9277 -1366
rect 9343 -1400 9373 -1366
rect 9509 -1388 9539 -1230
rect 9592 -1300 9622 -1106
rect 9789 -1205 9819 -1190
rect 9713 -1235 9819 -1205
rect 9713 -1252 9743 -1235
rect 9677 -1268 9743 -1252
rect 9581 -1316 9635 -1300
rect 9581 -1350 9591 -1316
rect 9625 -1350 9635 -1316
rect 9677 -1302 9687 -1268
rect 9721 -1302 9743 -1268
rect 9888 -1240 9918 -1106
rect 9974 -1138 10004 -1106
rect 9960 -1154 10014 -1138
rect 9960 -1188 9970 -1154
rect 10004 -1188 10014 -1154
rect 9960 -1204 10014 -1188
rect 9888 -1252 9938 -1240
rect 9888 -1264 9951 -1252
rect 9888 -1270 9975 -1264
rect 9909 -1280 9975 -1270
rect 9909 -1282 9931 -1280
rect 9677 -1318 9743 -1302
rect 9713 -1344 9743 -1318
rect 9812 -1328 9879 -1312
rect 9581 -1366 9635 -1350
rect 9581 -1388 9611 -1366
rect 9812 -1362 9835 -1328
rect 9869 -1362 9879 -1328
rect 9812 -1378 9879 -1362
rect 9921 -1314 9931 -1282
rect 9965 -1314 9975 -1280
rect 9921 -1330 9975 -1314
rect 10058 -1290 10088 -1106
rect 10166 -1262 10196 -1106
rect 10250 -1154 10280 -1106
rect 10238 -1170 10292 -1154
rect 10238 -1204 10248 -1170
rect 10282 -1204 10292 -1170
rect 10238 -1220 10292 -1204
rect 10161 -1278 10215 -1262
rect 10058 -1306 10119 -1290
rect 10058 -1326 10075 -1306
rect 9812 -1400 9842 -1378
rect 9921 -1400 9951 -1330
rect 10017 -1340 10075 -1326
rect 10109 -1340 10119 -1306
rect 10161 -1312 10171 -1278
rect 10205 -1312 10215 -1278
rect 10161 -1328 10215 -1312
rect 10017 -1356 10119 -1340
rect 10017 -1388 10047 -1356
rect 10166 -1388 10196 -1328
rect 10257 -1388 10287 -1220
rect 10633 -1186 10663 -1150
rect 10622 -1216 10663 -1186
rect 10414 -1254 10444 -1222
rect 10622 -1254 10652 -1216
rect 11279 -1028 11309 -1002
rect 11363 -1028 11393 -1002
rect 11630 -1022 11660 -996
rect 11722 -1022 11752 -996
rect 11821 -1022 11851 -996
rect 11961 -1022 11991 -996
rect 12058 -1022 12088 -996
rect 12255 -1022 12285 -996
rect 12354 -1022 12384 -996
rect 12440 -1022 12470 -996
rect 12524 -1022 12554 -996
rect 12632 -1022 12662 -996
rect 12716 -1022 12746 -996
rect 12880 -1022 12910 -996
rect 13099 -1022 13129 -996
rect 13196 -1022 13226 -996
rect 11279 -1171 11309 -1156
rect 11246 -1201 11309 -1171
rect 10730 -1254 10760 -1222
rect 11246 -1254 11276 -1201
rect 11363 -1245 11393 -1156
rect 11630 -1193 11660 -1106
rect 11722 -1144 11752 -1106
rect 10343 -1270 10652 -1254
rect 10343 -1304 10371 -1270
rect 10405 -1304 10652 -1270
rect 10343 -1320 10652 -1304
rect 10701 -1270 10760 -1254
rect 10701 -1304 10711 -1270
rect 10745 -1304 10760 -1270
rect 10701 -1320 10760 -1304
rect 11222 -1270 11276 -1254
rect 11222 -1304 11232 -1270
rect 11266 -1304 11276 -1270
rect 11318 -1255 11393 -1245
rect 11318 -1289 11334 -1255
rect 11368 -1289 11393 -1255
rect 11531 -1209 11660 -1193
rect 11706 -1154 11772 -1144
rect 11706 -1188 11722 -1154
rect 11756 -1188 11772 -1154
rect 11706 -1198 11772 -1188
rect 11531 -1243 11541 -1209
rect 11575 -1223 11660 -1209
rect 11575 -1243 11648 -1223
rect 11821 -1240 11851 -1106
rect 11961 -1164 11991 -1106
rect 11961 -1180 12016 -1164
rect 11961 -1214 11971 -1180
rect 12005 -1214 12016 -1180
rect 11961 -1230 12016 -1214
rect 11531 -1259 11648 -1243
rect 11318 -1299 11393 -1289
rect 11222 -1320 11276 -1304
rect 10445 -1342 10475 -1320
rect 10622 -1343 10652 -1320
rect 10730 -1342 10760 -1320
rect 10622 -1373 10663 -1343
rect 10633 -1388 10663 -1373
rect 11246 -1343 11276 -1320
rect 11246 -1373 11309 -1343
rect 11279 -1388 11309 -1373
rect 11363 -1388 11393 -1299
rect 11618 -1388 11648 -1259
rect 11713 -1270 11851 -1240
rect 11713 -1300 11744 -1270
rect 11690 -1316 11744 -1300
rect 11690 -1350 11700 -1316
rect 11734 -1350 11744 -1316
rect 11690 -1366 11744 -1350
rect 11786 -1322 11852 -1312
rect 11786 -1356 11802 -1322
rect 11836 -1356 11852 -1322
rect 11786 -1366 11852 -1356
rect 11713 -1400 11743 -1366
rect 11809 -1400 11839 -1366
rect 11975 -1388 12005 -1230
rect 12058 -1300 12088 -1106
rect 12255 -1205 12285 -1190
rect 12179 -1235 12285 -1205
rect 12179 -1252 12209 -1235
rect 12143 -1268 12209 -1252
rect 12047 -1316 12101 -1300
rect 12047 -1350 12057 -1316
rect 12091 -1350 12101 -1316
rect 12143 -1302 12153 -1268
rect 12187 -1302 12209 -1268
rect 12354 -1240 12384 -1106
rect 12440 -1138 12470 -1106
rect 12426 -1154 12480 -1138
rect 12426 -1188 12436 -1154
rect 12470 -1188 12480 -1154
rect 12426 -1204 12480 -1188
rect 12354 -1252 12404 -1240
rect 12354 -1264 12417 -1252
rect 12354 -1270 12441 -1264
rect 12375 -1280 12441 -1270
rect 12375 -1282 12397 -1280
rect 12143 -1318 12209 -1302
rect 12179 -1344 12209 -1318
rect 12278 -1328 12345 -1312
rect 12047 -1366 12101 -1350
rect 12047 -1388 12077 -1366
rect 12278 -1362 12301 -1328
rect 12335 -1362 12345 -1328
rect 12278 -1378 12345 -1362
rect 12387 -1314 12397 -1282
rect 12431 -1314 12441 -1280
rect 12387 -1330 12441 -1314
rect 12524 -1290 12554 -1106
rect 12632 -1262 12662 -1106
rect 12716 -1154 12746 -1106
rect 12704 -1170 12758 -1154
rect 12704 -1204 12714 -1170
rect 12748 -1204 12758 -1170
rect 12704 -1220 12758 -1204
rect 12627 -1278 12681 -1262
rect 12524 -1306 12585 -1290
rect 12524 -1326 12541 -1306
rect 12278 -1400 12308 -1378
rect 12387 -1400 12417 -1330
rect 12483 -1340 12541 -1326
rect 12575 -1340 12585 -1306
rect 12627 -1312 12637 -1278
rect 12671 -1312 12681 -1278
rect 12627 -1328 12681 -1312
rect 12483 -1356 12585 -1340
rect 12483 -1388 12513 -1356
rect 12632 -1388 12662 -1328
rect 12723 -1388 12753 -1220
rect 13099 -1186 13129 -1150
rect 13088 -1216 13129 -1186
rect 12880 -1254 12910 -1222
rect 13088 -1254 13118 -1216
rect 13196 -1254 13226 -1222
rect 12809 -1270 13118 -1254
rect 12809 -1304 12837 -1270
rect 12871 -1304 13118 -1270
rect 12809 -1320 13118 -1304
rect 13167 -1270 13226 -1254
rect 13167 -1304 13177 -1270
rect 13211 -1304 13226 -1270
rect 13167 -1320 13226 -1304
rect 12911 -1342 12941 -1320
rect 13088 -1343 13118 -1320
rect 13196 -1342 13226 -1320
rect 13088 -1373 13129 -1343
rect 13099 -1388 13129 -1373
rect 8813 -1498 8843 -1472
rect 8897 -1498 8927 -1472
rect 9152 -1498 9182 -1472
rect 9247 -1498 9277 -1472
rect 9343 -1498 9373 -1472
rect 9509 -1498 9539 -1472
rect 9581 -1498 9611 -1472
rect 9713 -1498 9743 -1472
rect 9812 -1498 9842 -1472
rect 9921 -1498 9951 -1472
rect 10017 -1498 10047 -1472
rect 10166 -1498 10196 -1472
rect 10257 -1498 10287 -1472
rect 10445 -1498 10475 -1472
rect 10633 -1498 10663 -1472
rect 10730 -1498 10760 -1472
rect 11279 -1498 11309 -1472
rect 11363 -1498 11393 -1472
rect 11618 -1498 11648 -1472
rect 11713 -1498 11743 -1472
rect 11809 -1498 11839 -1472
rect 11975 -1498 12005 -1472
rect 12047 -1498 12077 -1472
rect 12179 -1498 12209 -1472
rect 12278 -1498 12308 -1472
rect 12387 -1498 12417 -1472
rect 12483 -1498 12513 -1472
rect 12632 -1498 12662 -1472
rect 12723 -1498 12753 -1472
rect 12911 -1498 12941 -1472
rect 13099 -1498 13129 -1472
rect 13196 -1498 13226 -1472
rect 10233 -1824 10263 -1798
rect 10317 -1824 10347 -1798
rect 11279 -1830 11309 -1804
rect 11363 -1830 11393 -1804
rect 11630 -1824 11660 -1798
rect 11722 -1824 11752 -1798
rect 11821 -1824 11851 -1798
rect 11961 -1824 11991 -1798
rect 12058 -1824 12088 -1798
rect 12255 -1824 12285 -1798
rect 12354 -1824 12384 -1798
rect 12440 -1824 12470 -1798
rect 12524 -1824 12554 -1798
rect 12632 -1824 12662 -1798
rect 12716 -1824 12746 -1798
rect 12880 -1824 12910 -1798
rect 13099 -1824 13129 -1798
rect 13196 -1824 13226 -1798
rect 11279 -1973 11309 -1958
rect 11246 -2003 11309 -1973
rect 10233 -2056 10263 -2024
rect 10317 -2056 10347 -2024
rect 11246 -2056 11276 -2003
rect 11363 -2047 11393 -1958
rect 11630 -1995 11660 -1908
rect 11722 -1946 11752 -1908
rect 10173 -2072 10347 -2056
rect 10173 -2106 10189 -2072
rect 10223 -2106 10347 -2072
rect 10173 -2122 10347 -2106
rect 11222 -2072 11276 -2056
rect 11222 -2106 11232 -2072
rect 11266 -2106 11276 -2072
rect 11318 -2057 11393 -2047
rect 11318 -2091 11334 -2057
rect 11368 -2091 11393 -2057
rect 11531 -2011 11660 -1995
rect 11706 -1956 11772 -1946
rect 11706 -1990 11722 -1956
rect 11756 -1990 11772 -1956
rect 11706 -2000 11772 -1990
rect 11531 -2045 11541 -2011
rect 11575 -2025 11660 -2011
rect 11575 -2045 11648 -2025
rect 11821 -2042 11851 -1908
rect 11961 -1966 11991 -1908
rect 11961 -1982 12016 -1966
rect 11961 -2016 11971 -1982
rect 12005 -2016 12016 -1982
rect 11961 -2032 12016 -2016
rect 11531 -2061 11648 -2045
rect 11318 -2101 11393 -2091
rect 11222 -2122 11276 -2106
rect 10233 -2144 10263 -2122
rect 10317 -2144 10347 -2122
rect 11246 -2145 11276 -2122
rect 11246 -2175 11309 -2145
rect 11279 -2190 11309 -2175
rect 11363 -2190 11393 -2101
rect 11618 -2190 11648 -2061
rect 11713 -2072 11851 -2042
rect 11713 -2102 11744 -2072
rect 11690 -2118 11744 -2102
rect 11690 -2152 11700 -2118
rect 11734 -2152 11744 -2118
rect 11690 -2168 11744 -2152
rect 11786 -2124 11852 -2114
rect 11786 -2158 11802 -2124
rect 11836 -2158 11852 -2124
rect 11786 -2168 11852 -2158
rect 11713 -2202 11743 -2168
rect 11809 -2202 11839 -2168
rect 11975 -2190 12005 -2032
rect 12058 -2102 12088 -1908
rect 12255 -2007 12285 -1992
rect 12179 -2037 12285 -2007
rect 12179 -2054 12209 -2037
rect 12143 -2070 12209 -2054
rect 12047 -2118 12101 -2102
rect 12047 -2152 12057 -2118
rect 12091 -2152 12101 -2118
rect 12143 -2104 12153 -2070
rect 12187 -2104 12209 -2070
rect 12354 -2042 12384 -1908
rect 12440 -1940 12470 -1908
rect 12426 -1956 12480 -1940
rect 12426 -1990 12436 -1956
rect 12470 -1990 12480 -1956
rect 12426 -2006 12480 -1990
rect 12354 -2054 12404 -2042
rect 12354 -2066 12417 -2054
rect 12354 -2072 12441 -2066
rect 12375 -2082 12441 -2072
rect 12375 -2084 12397 -2082
rect 12143 -2120 12209 -2104
rect 12179 -2146 12209 -2120
rect 12278 -2130 12345 -2114
rect 12047 -2168 12101 -2152
rect 12047 -2190 12077 -2168
rect 12278 -2164 12301 -2130
rect 12335 -2164 12345 -2130
rect 12278 -2180 12345 -2164
rect 12387 -2116 12397 -2084
rect 12431 -2116 12441 -2082
rect 12387 -2132 12441 -2116
rect 12524 -2092 12554 -1908
rect 12632 -2064 12662 -1908
rect 12716 -1956 12746 -1908
rect 12704 -1972 12758 -1956
rect 12704 -2006 12714 -1972
rect 12748 -2006 12758 -1972
rect 12704 -2022 12758 -2006
rect 12627 -2080 12681 -2064
rect 12524 -2108 12585 -2092
rect 12524 -2128 12541 -2108
rect 12278 -2202 12308 -2180
rect 12387 -2202 12417 -2132
rect 12483 -2142 12541 -2128
rect 12575 -2142 12585 -2108
rect 12627 -2114 12637 -2080
rect 12671 -2114 12681 -2080
rect 12627 -2130 12681 -2114
rect 12483 -2158 12585 -2142
rect 12483 -2190 12513 -2158
rect 12632 -2190 12662 -2130
rect 12723 -2190 12753 -2022
rect 13099 -1988 13129 -1952
rect 13088 -2018 13129 -1988
rect 12880 -2056 12910 -2024
rect 13088 -2056 13118 -2018
rect 13196 -2056 13226 -2024
rect 12809 -2072 13118 -2056
rect 12809 -2106 12837 -2072
rect 12871 -2106 13118 -2072
rect 12809 -2122 13118 -2106
rect 13167 -2072 13226 -2056
rect 13167 -2106 13177 -2072
rect 13211 -2106 13226 -2072
rect 13167 -2122 13226 -2106
rect 12911 -2144 12941 -2122
rect 13088 -2145 13118 -2122
rect 13196 -2144 13226 -2122
rect 13088 -2175 13129 -2145
rect 13099 -2190 13129 -2175
rect 10233 -2300 10263 -2274
rect 10317 -2300 10347 -2274
rect 11279 -2300 11309 -2274
rect 11363 -2300 11393 -2274
rect 11618 -2300 11648 -2274
rect 11713 -2300 11743 -2274
rect 11809 -2300 11839 -2274
rect 11975 -2300 12005 -2274
rect 12047 -2300 12077 -2274
rect 12179 -2300 12209 -2274
rect 12278 -2300 12308 -2274
rect 12387 -2300 12417 -2274
rect 12483 -2300 12513 -2274
rect 12632 -2300 12662 -2274
rect 12723 -2300 12753 -2274
rect 12911 -2300 12941 -2274
rect 13099 -2300 13129 -2274
rect 13196 -2300 13226 -2274
rect -9079 -4298 -9049 -4272
rect -8995 -4298 -8965 -4272
rect -8728 -4292 -8698 -4266
rect -8636 -4292 -8606 -4266
rect -8537 -4292 -8507 -4266
rect -8397 -4292 -8367 -4266
rect -8300 -4292 -8270 -4266
rect -8103 -4292 -8073 -4266
rect -8004 -4292 -7974 -4266
rect -7918 -4292 -7888 -4266
rect -7834 -4292 -7804 -4266
rect -7726 -4292 -7696 -4266
rect -7642 -4292 -7612 -4266
rect -7478 -4292 -7448 -4266
rect -7259 -4292 -7229 -4266
rect -7162 -4292 -7132 -4266
rect -9079 -4441 -9049 -4426
rect -9112 -4471 -9049 -4441
rect -9112 -4524 -9082 -4471
rect -8995 -4515 -8965 -4426
rect -8728 -4463 -8698 -4376
rect -8636 -4414 -8606 -4376
rect -9136 -4540 -9082 -4524
rect -9136 -4574 -9126 -4540
rect -9092 -4574 -9082 -4540
rect -9040 -4525 -8965 -4515
rect -9040 -4559 -9024 -4525
rect -8990 -4559 -8965 -4525
rect -8827 -4479 -8698 -4463
rect -8652 -4424 -8586 -4414
rect -8652 -4458 -8636 -4424
rect -8602 -4458 -8586 -4424
rect -8652 -4468 -8586 -4458
rect -8827 -4513 -8817 -4479
rect -8783 -4493 -8698 -4479
rect -8783 -4513 -8710 -4493
rect -8537 -4510 -8507 -4376
rect -8397 -4434 -8367 -4376
rect -8397 -4450 -8342 -4434
rect -8397 -4484 -8387 -4450
rect -8353 -4484 -8342 -4450
rect -8397 -4500 -8342 -4484
rect -8827 -4529 -8710 -4513
rect -9040 -4569 -8965 -4559
rect -9136 -4590 -9082 -4574
rect -9112 -4613 -9082 -4590
rect -9112 -4643 -9049 -4613
rect -9079 -4658 -9049 -4643
rect -8995 -4658 -8965 -4569
rect -8740 -4658 -8710 -4529
rect -8645 -4540 -8507 -4510
rect -8645 -4570 -8614 -4540
rect -8668 -4586 -8614 -4570
rect -8668 -4620 -8658 -4586
rect -8624 -4620 -8614 -4586
rect -8668 -4636 -8614 -4620
rect -8572 -4592 -8506 -4582
rect -8572 -4626 -8556 -4592
rect -8522 -4626 -8506 -4592
rect -8572 -4636 -8506 -4626
rect -8645 -4670 -8615 -4636
rect -8549 -4670 -8519 -4636
rect -8383 -4658 -8353 -4500
rect -8300 -4570 -8270 -4376
rect -8103 -4475 -8073 -4460
rect -8179 -4505 -8073 -4475
rect -8179 -4522 -8149 -4505
rect -8215 -4538 -8149 -4522
rect -8311 -4586 -8257 -4570
rect -8311 -4620 -8301 -4586
rect -8267 -4620 -8257 -4586
rect -8215 -4572 -8205 -4538
rect -8171 -4572 -8149 -4538
rect -8004 -4510 -7974 -4376
rect -7918 -4408 -7888 -4376
rect -7932 -4424 -7878 -4408
rect -7932 -4458 -7922 -4424
rect -7888 -4458 -7878 -4424
rect -7932 -4474 -7878 -4458
rect -8004 -4522 -7954 -4510
rect -8004 -4534 -7941 -4522
rect -8004 -4540 -7917 -4534
rect -7983 -4550 -7917 -4540
rect -7983 -4552 -7961 -4550
rect -8215 -4588 -8149 -4572
rect -8179 -4614 -8149 -4588
rect -8080 -4598 -8013 -4582
rect -8311 -4636 -8257 -4620
rect -8311 -4658 -8281 -4636
rect -8080 -4632 -8057 -4598
rect -8023 -4632 -8013 -4598
rect -8080 -4648 -8013 -4632
rect -7971 -4584 -7961 -4552
rect -7927 -4584 -7917 -4550
rect -7971 -4600 -7917 -4584
rect -7834 -4560 -7804 -4376
rect -7726 -4532 -7696 -4376
rect -7642 -4424 -7612 -4376
rect -7654 -4440 -7600 -4424
rect -7654 -4474 -7644 -4440
rect -7610 -4474 -7600 -4440
rect -7654 -4490 -7600 -4474
rect -7731 -4548 -7677 -4532
rect -7834 -4576 -7773 -4560
rect -7834 -4596 -7817 -4576
rect -8080 -4670 -8050 -4648
rect -7971 -4670 -7941 -4600
rect -7875 -4610 -7817 -4596
rect -7783 -4610 -7773 -4576
rect -7731 -4582 -7721 -4548
rect -7687 -4582 -7677 -4548
rect -7731 -4598 -7677 -4582
rect -7875 -4626 -7773 -4610
rect -7875 -4658 -7845 -4626
rect -7726 -4658 -7696 -4598
rect -7635 -4658 -7605 -4490
rect -7259 -4456 -7229 -4420
rect -7270 -4486 -7229 -4456
rect -7478 -4524 -7448 -4492
rect -7270 -4524 -7240 -4486
rect -6963 -4298 -6933 -4272
rect -6879 -4298 -6849 -4272
rect -6612 -4292 -6582 -4266
rect -6520 -4292 -6490 -4266
rect -6421 -4292 -6391 -4266
rect -6281 -4292 -6251 -4266
rect -6184 -4292 -6154 -4266
rect -5987 -4292 -5957 -4266
rect -5888 -4292 -5858 -4266
rect -5802 -4292 -5772 -4266
rect -5718 -4292 -5688 -4266
rect -5610 -4292 -5580 -4266
rect -5526 -4292 -5496 -4266
rect -5362 -4292 -5332 -4266
rect -5143 -4292 -5113 -4266
rect -5046 -4292 -5016 -4266
rect -6963 -4441 -6933 -4426
rect -6996 -4471 -6933 -4441
rect -7162 -4524 -7132 -4492
rect -6996 -4524 -6966 -4471
rect -6879 -4515 -6849 -4426
rect -6612 -4463 -6582 -4376
rect -6520 -4414 -6490 -4376
rect -7549 -4540 -7240 -4524
rect -7549 -4574 -7521 -4540
rect -7487 -4574 -7240 -4540
rect -7549 -4590 -7240 -4574
rect -7191 -4540 -7132 -4524
rect -7191 -4574 -7181 -4540
rect -7147 -4574 -7132 -4540
rect -7191 -4590 -7132 -4574
rect -7020 -4540 -6966 -4524
rect -7020 -4574 -7010 -4540
rect -6976 -4574 -6966 -4540
rect -6924 -4525 -6849 -4515
rect -6924 -4559 -6908 -4525
rect -6874 -4559 -6849 -4525
rect -6711 -4479 -6582 -4463
rect -6536 -4424 -6470 -4414
rect -6536 -4458 -6520 -4424
rect -6486 -4458 -6470 -4424
rect -6536 -4468 -6470 -4458
rect -6711 -4513 -6701 -4479
rect -6667 -4493 -6582 -4479
rect -6667 -4513 -6594 -4493
rect -6421 -4510 -6391 -4376
rect -6281 -4434 -6251 -4376
rect -6281 -4450 -6226 -4434
rect -6281 -4484 -6271 -4450
rect -6237 -4484 -6226 -4450
rect -6281 -4500 -6226 -4484
rect -6711 -4529 -6594 -4513
rect -6924 -4569 -6849 -4559
rect -7020 -4590 -6966 -4574
rect -7447 -4612 -7417 -4590
rect -7270 -4613 -7240 -4590
rect -7162 -4612 -7132 -4590
rect -7270 -4643 -7229 -4613
rect -7259 -4658 -7229 -4643
rect -6996 -4613 -6966 -4590
rect -6996 -4643 -6933 -4613
rect -6963 -4658 -6933 -4643
rect -6879 -4658 -6849 -4569
rect -6624 -4658 -6594 -4529
rect -6529 -4540 -6391 -4510
rect -6529 -4570 -6498 -4540
rect -6552 -4586 -6498 -4570
rect -6552 -4620 -6542 -4586
rect -6508 -4620 -6498 -4586
rect -6552 -4636 -6498 -4620
rect -6456 -4592 -6390 -4582
rect -6456 -4626 -6440 -4592
rect -6406 -4626 -6390 -4592
rect -6456 -4636 -6390 -4626
rect -6529 -4670 -6499 -4636
rect -6433 -4670 -6403 -4636
rect -6267 -4658 -6237 -4500
rect -6184 -4570 -6154 -4376
rect -5987 -4475 -5957 -4460
rect -6063 -4505 -5957 -4475
rect -6063 -4522 -6033 -4505
rect -6099 -4538 -6033 -4522
rect -6195 -4586 -6141 -4570
rect -6195 -4620 -6185 -4586
rect -6151 -4620 -6141 -4586
rect -6099 -4572 -6089 -4538
rect -6055 -4572 -6033 -4538
rect -5888 -4510 -5858 -4376
rect -5802 -4408 -5772 -4376
rect -5816 -4424 -5762 -4408
rect -5816 -4458 -5806 -4424
rect -5772 -4458 -5762 -4424
rect -5816 -4474 -5762 -4458
rect -5888 -4522 -5838 -4510
rect -5888 -4534 -5825 -4522
rect -5888 -4540 -5801 -4534
rect -5867 -4550 -5801 -4540
rect -5867 -4552 -5845 -4550
rect -6099 -4588 -6033 -4572
rect -6063 -4614 -6033 -4588
rect -5964 -4598 -5897 -4582
rect -6195 -4636 -6141 -4620
rect -6195 -4658 -6165 -4636
rect -5964 -4632 -5941 -4598
rect -5907 -4632 -5897 -4598
rect -5964 -4648 -5897 -4632
rect -5855 -4584 -5845 -4552
rect -5811 -4584 -5801 -4550
rect -5855 -4600 -5801 -4584
rect -5718 -4560 -5688 -4376
rect -5610 -4532 -5580 -4376
rect -5526 -4424 -5496 -4376
rect -5538 -4440 -5484 -4424
rect -5538 -4474 -5528 -4440
rect -5494 -4474 -5484 -4440
rect -5538 -4490 -5484 -4474
rect -5615 -4548 -5561 -4532
rect -5718 -4576 -5657 -4560
rect -5718 -4596 -5701 -4576
rect -5964 -4670 -5934 -4648
rect -5855 -4670 -5825 -4600
rect -5759 -4610 -5701 -4596
rect -5667 -4610 -5657 -4576
rect -5615 -4582 -5605 -4548
rect -5571 -4582 -5561 -4548
rect -5615 -4598 -5561 -4582
rect -5759 -4626 -5657 -4610
rect -5759 -4658 -5729 -4626
rect -5610 -4658 -5580 -4598
rect -5519 -4658 -5489 -4490
rect -5143 -4456 -5113 -4420
rect -5154 -4486 -5113 -4456
rect -5362 -4524 -5332 -4492
rect -5154 -4524 -5124 -4486
rect -4847 -4298 -4817 -4272
rect -4763 -4298 -4733 -4272
rect -4496 -4292 -4466 -4266
rect -4404 -4292 -4374 -4266
rect -4305 -4292 -4275 -4266
rect -4165 -4292 -4135 -4266
rect -4068 -4292 -4038 -4266
rect -3871 -4292 -3841 -4266
rect -3772 -4292 -3742 -4266
rect -3686 -4292 -3656 -4266
rect -3602 -4292 -3572 -4266
rect -3494 -4292 -3464 -4266
rect -3410 -4292 -3380 -4266
rect -3246 -4292 -3216 -4266
rect -3027 -4292 -2997 -4266
rect -2930 -4292 -2900 -4266
rect -4847 -4441 -4817 -4426
rect -4880 -4471 -4817 -4441
rect -5046 -4524 -5016 -4492
rect -4880 -4524 -4850 -4471
rect -4763 -4515 -4733 -4426
rect -4496 -4463 -4466 -4376
rect -4404 -4414 -4374 -4376
rect -5433 -4540 -5124 -4524
rect -5433 -4574 -5405 -4540
rect -5371 -4574 -5124 -4540
rect -5433 -4590 -5124 -4574
rect -5075 -4540 -5016 -4524
rect -5075 -4574 -5065 -4540
rect -5031 -4574 -5016 -4540
rect -5075 -4590 -5016 -4574
rect -4904 -4540 -4850 -4524
rect -4904 -4574 -4894 -4540
rect -4860 -4574 -4850 -4540
rect -4808 -4525 -4733 -4515
rect -4808 -4559 -4792 -4525
rect -4758 -4559 -4733 -4525
rect -4595 -4479 -4466 -4463
rect -4420 -4424 -4354 -4414
rect -4420 -4458 -4404 -4424
rect -4370 -4458 -4354 -4424
rect -4420 -4468 -4354 -4458
rect -4595 -4513 -4585 -4479
rect -4551 -4493 -4466 -4479
rect -4551 -4513 -4478 -4493
rect -4305 -4510 -4275 -4376
rect -4165 -4434 -4135 -4376
rect -4165 -4450 -4110 -4434
rect -4165 -4484 -4155 -4450
rect -4121 -4484 -4110 -4450
rect -4165 -4500 -4110 -4484
rect -4595 -4529 -4478 -4513
rect -4808 -4569 -4733 -4559
rect -4904 -4590 -4850 -4574
rect -5331 -4612 -5301 -4590
rect -5154 -4613 -5124 -4590
rect -5046 -4612 -5016 -4590
rect -5154 -4643 -5113 -4613
rect -5143 -4658 -5113 -4643
rect -4880 -4613 -4850 -4590
rect -4880 -4643 -4817 -4613
rect -4847 -4658 -4817 -4643
rect -4763 -4658 -4733 -4569
rect -4508 -4658 -4478 -4529
rect -4413 -4540 -4275 -4510
rect -4413 -4570 -4382 -4540
rect -4436 -4586 -4382 -4570
rect -4436 -4620 -4426 -4586
rect -4392 -4620 -4382 -4586
rect -4436 -4636 -4382 -4620
rect -4340 -4592 -4274 -4582
rect -4340 -4626 -4324 -4592
rect -4290 -4626 -4274 -4592
rect -4340 -4636 -4274 -4626
rect -4413 -4670 -4383 -4636
rect -4317 -4670 -4287 -4636
rect -4151 -4658 -4121 -4500
rect -4068 -4570 -4038 -4376
rect -3871 -4475 -3841 -4460
rect -3947 -4505 -3841 -4475
rect -3947 -4522 -3917 -4505
rect -3983 -4538 -3917 -4522
rect -4079 -4586 -4025 -4570
rect -4079 -4620 -4069 -4586
rect -4035 -4620 -4025 -4586
rect -3983 -4572 -3973 -4538
rect -3939 -4572 -3917 -4538
rect -3772 -4510 -3742 -4376
rect -3686 -4408 -3656 -4376
rect -3700 -4424 -3646 -4408
rect -3700 -4458 -3690 -4424
rect -3656 -4458 -3646 -4424
rect -3700 -4474 -3646 -4458
rect -3772 -4522 -3722 -4510
rect -3772 -4534 -3709 -4522
rect -3772 -4540 -3685 -4534
rect -3751 -4550 -3685 -4540
rect -3751 -4552 -3729 -4550
rect -3983 -4588 -3917 -4572
rect -3947 -4614 -3917 -4588
rect -3848 -4598 -3781 -4582
rect -4079 -4636 -4025 -4620
rect -4079 -4658 -4049 -4636
rect -3848 -4632 -3825 -4598
rect -3791 -4632 -3781 -4598
rect -3848 -4648 -3781 -4632
rect -3739 -4584 -3729 -4552
rect -3695 -4584 -3685 -4550
rect -3739 -4600 -3685 -4584
rect -3602 -4560 -3572 -4376
rect -3494 -4532 -3464 -4376
rect -3410 -4424 -3380 -4376
rect -3422 -4440 -3368 -4424
rect -3422 -4474 -3412 -4440
rect -3378 -4474 -3368 -4440
rect -3422 -4490 -3368 -4474
rect -3499 -4548 -3445 -4532
rect -3602 -4576 -3541 -4560
rect -3602 -4596 -3585 -4576
rect -3848 -4670 -3818 -4648
rect -3739 -4670 -3709 -4600
rect -3643 -4610 -3585 -4596
rect -3551 -4610 -3541 -4576
rect -3499 -4582 -3489 -4548
rect -3455 -4582 -3445 -4548
rect -3499 -4598 -3445 -4582
rect -3643 -4626 -3541 -4610
rect -3643 -4658 -3613 -4626
rect -3494 -4658 -3464 -4598
rect -3403 -4658 -3373 -4490
rect -3027 -4456 -2997 -4420
rect -3038 -4486 -2997 -4456
rect -3246 -4524 -3216 -4492
rect -3038 -4524 -3008 -4486
rect -2731 -4298 -2701 -4272
rect -2647 -4298 -2617 -4272
rect -2380 -4292 -2350 -4266
rect -2288 -4292 -2258 -4266
rect -2189 -4292 -2159 -4266
rect -2049 -4292 -2019 -4266
rect -1952 -4292 -1922 -4266
rect -1755 -4292 -1725 -4266
rect -1656 -4292 -1626 -4266
rect -1570 -4292 -1540 -4266
rect -1486 -4292 -1456 -4266
rect -1378 -4292 -1348 -4266
rect -1294 -4292 -1264 -4266
rect -1130 -4292 -1100 -4266
rect -911 -4292 -881 -4266
rect -814 -4292 -784 -4266
rect -2731 -4441 -2701 -4426
rect -2764 -4471 -2701 -4441
rect -2930 -4524 -2900 -4492
rect -2764 -4524 -2734 -4471
rect -2647 -4515 -2617 -4426
rect -2380 -4463 -2350 -4376
rect -2288 -4414 -2258 -4376
rect -3317 -4540 -3008 -4524
rect -3317 -4574 -3289 -4540
rect -3255 -4574 -3008 -4540
rect -3317 -4590 -3008 -4574
rect -2959 -4540 -2900 -4524
rect -2959 -4574 -2949 -4540
rect -2915 -4574 -2900 -4540
rect -2959 -4590 -2900 -4574
rect -2788 -4540 -2734 -4524
rect -2788 -4574 -2778 -4540
rect -2744 -4574 -2734 -4540
rect -2692 -4525 -2617 -4515
rect -2692 -4559 -2676 -4525
rect -2642 -4559 -2617 -4525
rect -2479 -4479 -2350 -4463
rect -2304 -4424 -2238 -4414
rect -2304 -4458 -2288 -4424
rect -2254 -4458 -2238 -4424
rect -2304 -4468 -2238 -4458
rect -2479 -4513 -2469 -4479
rect -2435 -4493 -2350 -4479
rect -2435 -4513 -2362 -4493
rect -2189 -4510 -2159 -4376
rect -2049 -4434 -2019 -4376
rect -2049 -4450 -1994 -4434
rect -2049 -4484 -2039 -4450
rect -2005 -4484 -1994 -4450
rect -2049 -4500 -1994 -4484
rect -2479 -4529 -2362 -4513
rect -2692 -4569 -2617 -4559
rect -2788 -4590 -2734 -4574
rect -3215 -4612 -3185 -4590
rect -3038 -4613 -3008 -4590
rect -2930 -4612 -2900 -4590
rect -3038 -4643 -2997 -4613
rect -3027 -4658 -2997 -4643
rect -2764 -4613 -2734 -4590
rect -2764 -4643 -2701 -4613
rect -2731 -4658 -2701 -4643
rect -2647 -4658 -2617 -4569
rect -2392 -4658 -2362 -4529
rect -2297 -4540 -2159 -4510
rect -2297 -4570 -2266 -4540
rect -2320 -4586 -2266 -4570
rect -2320 -4620 -2310 -4586
rect -2276 -4620 -2266 -4586
rect -2320 -4636 -2266 -4620
rect -2224 -4592 -2158 -4582
rect -2224 -4626 -2208 -4592
rect -2174 -4626 -2158 -4592
rect -2224 -4636 -2158 -4626
rect -2297 -4670 -2267 -4636
rect -2201 -4670 -2171 -4636
rect -2035 -4658 -2005 -4500
rect -1952 -4570 -1922 -4376
rect -1755 -4475 -1725 -4460
rect -1831 -4505 -1725 -4475
rect -1831 -4522 -1801 -4505
rect -1867 -4538 -1801 -4522
rect -1963 -4586 -1909 -4570
rect -1963 -4620 -1953 -4586
rect -1919 -4620 -1909 -4586
rect -1867 -4572 -1857 -4538
rect -1823 -4572 -1801 -4538
rect -1656 -4510 -1626 -4376
rect -1570 -4408 -1540 -4376
rect -1584 -4424 -1530 -4408
rect -1584 -4458 -1574 -4424
rect -1540 -4458 -1530 -4424
rect -1584 -4474 -1530 -4458
rect -1656 -4522 -1606 -4510
rect -1656 -4534 -1593 -4522
rect -1656 -4540 -1569 -4534
rect -1635 -4550 -1569 -4540
rect -1635 -4552 -1613 -4550
rect -1867 -4588 -1801 -4572
rect -1831 -4614 -1801 -4588
rect -1732 -4598 -1665 -4582
rect -1963 -4636 -1909 -4620
rect -1963 -4658 -1933 -4636
rect -1732 -4632 -1709 -4598
rect -1675 -4632 -1665 -4598
rect -1732 -4648 -1665 -4632
rect -1623 -4584 -1613 -4552
rect -1579 -4584 -1569 -4550
rect -1623 -4600 -1569 -4584
rect -1486 -4560 -1456 -4376
rect -1378 -4532 -1348 -4376
rect -1294 -4424 -1264 -4376
rect -1306 -4440 -1252 -4424
rect -1306 -4474 -1296 -4440
rect -1262 -4474 -1252 -4440
rect -1306 -4490 -1252 -4474
rect -1383 -4548 -1329 -4532
rect -1486 -4576 -1425 -4560
rect -1486 -4596 -1469 -4576
rect -1732 -4670 -1702 -4648
rect -1623 -4670 -1593 -4600
rect -1527 -4610 -1469 -4596
rect -1435 -4610 -1425 -4576
rect -1383 -4582 -1373 -4548
rect -1339 -4582 -1329 -4548
rect -1383 -4598 -1329 -4582
rect -1527 -4626 -1425 -4610
rect -1527 -4658 -1497 -4626
rect -1378 -4658 -1348 -4598
rect -1287 -4658 -1257 -4490
rect -911 -4456 -881 -4420
rect -922 -4486 -881 -4456
rect -1130 -4524 -1100 -4492
rect -922 -4524 -892 -4486
rect -615 -4298 -585 -4272
rect -531 -4298 -501 -4272
rect -264 -4292 -234 -4266
rect -172 -4292 -142 -4266
rect -73 -4292 -43 -4266
rect 67 -4292 97 -4266
rect 164 -4292 194 -4266
rect 361 -4292 391 -4266
rect 460 -4292 490 -4266
rect 546 -4292 576 -4266
rect 630 -4292 660 -4266
rect 738 -4292 768 -4266
rect 822 -4292 852 -4266
rect 986 -4292 1016 -4266
rect 1205 -4292 1235 -4266
rect 1302 -4292 1332 -4266
rect -615 -4441 -585 -4426
rect -648 -4471 -585 -4441
rect -814 -4524 -784 -4492
rect -648 -4524 -618 -4471
rect -531 -4515 -501 -4426
rect -264 -4463 -234 -4376
rect -172 -4414 -142 -4376
rect -1201 -4540 -892 -4524
rect -1201 -4574 -1173 -4540
rect -1139 -4574 -892 -4540
rect -1201 -4590 -892 -4574
rect -843 -4540 -784 -4524
rect -843 -4574 -833 -4540
rect -799 -4574 -784 -4540
rect -843 -4590 -784 -4574
rect -672 -4540 -618 -4524
rect -672 -4574 -662 -4540
rect -628 -4574 -618 -4540
rect -576 -4525 -501 -4515
rect -576 -4559 -560 -4525
rect -526 -4559 -501 -4525
rect -363 -4479 -234 -4463
rect -188 -4424 -122 -4414
rect -188 -4458 -172 -4424
rect -138 -4458 -122 -4424
rect -188 -4468 -122 -4458
rect -363 -4513 -353 -4479
rect -319 -4493 -234 -4479
rect -319 -4513 -246 -4493
rect -73 -4510 -43 -4376
rect 67 -4434 97 -4376
rect 67 -4450 122 -4434
rect 67 -4484 77 -4450
rect 111 -4484 122 -4450
rect 67 -4500 122 -4484
rect -363 -4529 -246 -4513
rect -576 -4569 -501 -4559
rect -672 -4590 -618 -4574
rect -1099 -4612 -1069 -4590
rect -922 -4613 -892 -4590
rect -814 -4612 -784 -4590
rect -922 -4643 -881 -4613
rect -911 -4658 -881 -4643
rect -648 -4613 -618 -4590
rect -648 -4643 -585 -4613
rect -615 -4658 -585 -4643
rect -531 -4658 -501 -4569
rect -276 -4658 -246 -4529
rect -181 -4540 -43 -4510
rect -181 -4570 -150 -4540
rect -204 -4586 -150 -4570
rect -204 -4620 -194 -4586
rect -160 -4620 -150 -4586
rect -204 -4636 -150 -4620
rect -108 -4592 -42 -4582
rect -108 -4626 -92 -4592
rect -58 -4626 -42 -4592
rect -108 -4636 -42 -4626
rect -181 -4670 -151 -4636
rect -85 -4670 -55 -4636
rect 81 -4658 111 -4500
rect 164 -4570 194 -4376
rect 361 -4475 391 -4460
rect 285 -4505 391 -4475
rect 285 -4522 315 -4505
rect 249 -4538 315 -4522
rect 153 -4586 207 -4570
rect 153 -4620 163 -4586
rect 197 -4620 207 -4586
rect 249 -4572 259 -4538
rect 293 -4572 315 -4538
rect 460 -4510 490 -4376
rect 546 -4408 576 -4376
rect 532 -4424 586 -4408
rect 532 -4458 542 -4424
rect 576 -4458 586 -4424
rect 532 -4474 586 -4458
rect 460 -4522 510 -4510
rect 460 -4534 523 -4522
rect 460 -4540 547 -4534
rect 481 -4550 547 -4540
rect 481 -4552 503 -4550
rect 249 -4588 315 -4572
rect 285 -4614 315 -4588
rect 384 -4598 451 -4582
rect 153 -4636 207 -4620
rect 153 -4658 183 -4636
rect 384 -4632 407 -4598
rect 441 -4632 451 -4598
rect 384 -4648 451 -4632
rect 493 -4584 503 -4552
rect 537 -4584 547 -4550
rect 493 -4600 547 -4584
rect 630 -4560 660 -4376
rect 738 -4532 768 -4376
rect 822 -4424 852 -4376
rect 810 -4440 864 -4424
rect 810 -4474 820 -4440
rect 854 -4474 864 -4440
rect 810 -4490 864 -4474
rect 733 -4548 787 -4532
rect 630 -4576 691 -4560
rect 630 -4596 647 -4576
rect 384 -4670 414 -4648
rect 493 -4670 523 -4600
rect 589 -4610 647 -4596
rect 681 -4610 691 -4576
rect 733 -4582 743 -4548
rect 777 -4582 787 -4548
rect 733 -4598 787 -4582
rect 589 -4626 691 -4610
rect 589 -4658 619 -4626
rect 738 -4658 768 -4598
rect 829 -4658 859 -4490
rect 1205 -4456 1235 -4420
rect 1194 -4486 1235 -4456
rect 986 -4524 1016 -4492
rect 1194 -4524 1224 -4486
rect 1501 -4298 1531 -4272
rect 1585 -4298 1615 -4272
rect 1852 -4292 1882 -4266
rect 1944 -4292 1974 -4266
rect 2043 -4292 2073 -4266
rect 2183 -4292 2213 -4266
rect 2280 -4292 2310 -4266
rect 2477 -4292 2507 -4266
rect 2576 -4292 2606 -4266
rect 2662 -4292 2692 -4266
rect 2746 -4292 2776 -4266
rect 2854 -4292 2884 -4266
rect 2938 -4292 2968 -4266
rect 3102 -4292 3132 -4266
rect 3321 -4292 3351 -4266
rect 3418 -4292 3448 -4266
rect 1501 -4441 1531 -4426
rect 1468 -4471 1531 -4441
rect 1302 -4524 1332 -4492
rect 1468 -4524 1498 -4471
rect 1585 -4515 1615 -4426
rect 1852 -4463 1882 -4376
rect 1944 -4414 1974 -4376
rect 915 -4540 1224 -4524
rect 915 -4574 943 -4540
rect 977 -4574 1224 -4540
rect 915 -4590 1224 -4574
rect 1273 -4540 1332 -4524
rect 1273 -4574 1283 -4540
rect 1317 -4574 1332 -4540
rect 1273 -4590 1332 -4574
rect 1444 -4540 1498 -4524
rect 1444 -4574 1454 -4540
rect 1488 -4574 1498 -4540
rect 1540 -4525 1615 -4515
rect 1540 -4559 1556 -4525
rect 1590 -4559 1615 -4525
rect 1753 -4479 1882 -4463
rect 1928 -4424 1994 -4414
rect 1928 -4458 1944 -4424
rect 1978 -4458 1994 -4424
rect 1928 -4468 1994 -4458
rect 1753 -4513 1763 -4479
rect 1797 -4493 1882 -4479
rect 1797 -4513 1870 -4493
rect 2043 -4510 2073 -4376
rect 2183 -4434 2213 -4376
rect 2183 -4450 2238 -4434
rect 2183 -4484 2193 -4450
rect 2227 -4484 2238 -4450
rect 2183 -4500 2238 -4484
rect 1753 -4529 1870 -4513
rect 1540 -4569 1615 -4559
rect 1444 -4590 1498 -4574
rect 1017 -4612 1047 -4590
rect 1194 -4613 1224 -4590
rect 1302 -4612 1332 -4590
rect 1194 -4643 1235 -4613
rect 1205 -4658 1235 -4643
rect 1468 -4613 1498 -4590
rect 1468 -4643 1531 -4613
rect 1501 -4658 1531 -4643
rect 1585 -4658 1615 -4569
rect 1840 -4658 1870 -4529
rect 1935 -4540 2073 -4510
rect 1935 -4570 1966 -4540
rect 1912 -4586 1966 -4570
rect 1912 -4620 1922 -4586
rect 1956 -4620 1966 -4586
rect 1912 -4636 1966 -4620
rect 2008 -4592 2074 -4582
rect 2008 -4626 2024 -4592
rect 2058 -4626 2074 -4592
rect 2008 -4636 2074 -4626
rect 1935 -4670 1965 -4636
rect 2031 -4670 2061 -4636
rect 2197 -4658 2227 -4500
rect 2280 -4570 2310 -4376
rect 2477 -4475 2507 -4460
rect 2401 -4505 2507 -4475
rect 2401 -4522 2431 -4505
rect 2365 -4538 2431 -4522
rect 2269 -4586 2323 -4570
rect 2269 -4620 2279 -4586
rect 2313 -4620 2323 -4586
rect 2365 -4572 2375 -4538
rect 2409 -4572 2431 -4538
rect 2576 -4510 2606 -4376
rect 2662 -4408 2692 -4376
rect 2648 -4424 2702 -4408
rect 2648 -4458 2658 -4424
rect 2692 -4458 2702 -4424
rect 2648 -4474 2702 -4458
rect 2576 -4522 2626 -4510
rect 2576 -4534 2639 -4522
rect 2576 -4540 2663 -4534
rect 2597 -4550 2663 -4540
rect 2597 -4552 2619 -4550
rect 2365 -4588 2431 -4572
rect 2401 -4614 2431 -4588
rect 2500 -4598 2567 -4582
rect 2269 -4636 2323 -4620
rect 2269 -4658 2299 -4636
rect 2500 -4632 2523 -4598
rect 2557 -4632 2567 -4598
rect 2500 -4648 2567 -4632
rect 2609 -4584 2619 -4552
rect 2653 -4584 2663 -4550
rect 2609 -4600 2663 -4584
rect 2746 -4560 2776 -4376
rect 2854 -4532 2884 -4376
rect 2938 -4424 2968 -4376
rect 2926 -4440 2980 -4424
rect 2926 -4474 2936 -4440
rect 2970 -4474 2980 -4440
rect 2926 -4490 2980 -4474
rect 2849 -4548 2903 -4532
rect 2746 -4576 2807 -4560
rect 2746 -4596 2763 -4576
rect 2500 -4670 2530 -4648
rect 2609 -4670 2639 -4600
rect 2705 -4610 2763 -4596
rect 2797 -4610 2807 -4576
rect 2849 -4582 2859 -4548
rect 2893 -4582 2903 -4548
rect 2849 -4598 2903 -4582
rect 2705 -4626 2807 -4610
rect 2705 -4658 2735 -4626
rect 2854 -4658 2884 -4598
rect 2945 -4658 2975 -4490
rect 3321 -4456 3351 -4420
rect 3310 -4486 3351 -4456
rect 3102 -4524 3132 -4492
rect 3310 -4524 3340 -4486
rect 3617 -4298 3647 -4272
rect 3701 -4298 3731 -4272
rect 3968 -4292 3998 -4266
rect 4060 -4292 4090 -4266
rect 4159 -4292 4189 -4266
rect 4299 -4292 4329 -4266
rect 4396 -4292 4426 -4266
rect 4593 -4292 4623 -4266
rect 4692 -4292 4722 -4266
rect 4778 -4292 4808 -4266
rect 4862 -4292 4892 -4266
rect 4970 -4292 5000 -4266
rect 5054 -4292 5084 -4266
rect 5218 -4292 5248 -4266
rect 5437 -4292 5467 -4266
rect 5534 -4292 5564 -4266
rect 3617 -4441 3647 -4426
rect 3584 -4471 3647 -4441
rect 3418 -4524 3448 -4492
rect 3584 -4524 3614 -4471
rect 3701 -4515 3731 -4426
rect 3968 -4463 3998 -4376
rect 4060 -4414 4090 -4376
rect 3031 -4540 3340 -4524
rect 3031 -4574 3059 -4540
rect 3093 -4574 3340 -4540
rect 3031 -4590 3340 -4574
rect 3389 -4540 3448 -4524
rect 3389 -4574 3399 -4540
rect 3433 -4574 3448 -4540
rect 3389 -4590 3448 -4574
rect 3560 -4540 3614 -4524
rect 3560 -4574 3570 -4540
rect 3604 -4574 3614 -4540
rect 3656 -4525 3731 -4515
rect 3656 -4559 3672 -4525
rect 3706 -4559 3731 -4525
rect 3869 -4479 3998 -4463
rect 4044 -4424 4110 -4414
rect 4044 -4458 4060 -4424
rect 4094 -4458 4110 -4424
rect 4044 -4468 4110 -4458
rect 3869 -4513 3879 -4479
rect 3913 -4493 3998 -4479
rect 3913 -4513 3986 -4493
rect 4159 -4510 4189 -4376
rect 4299 -4434 4329 -4376
rect 4299 -4450 4354 -4434
rect 4299 -4484 4309 -4450
rect 4343 -4484 4354 -4450
rect 4299 -4500 4354 -4484
rect 3869 -4529 3986 -4513
rect 3656 -4569 3731 -4559
rect 3560 -4590 3614 -4574
rect 3133 -4612 3163 -4590
rect 3310 -4613 3340 -4590
rect 3418 -4612 3448 -4590
rect 3310 -4643 3351 -4613
rect 3321 -4658 3351 -4643
rect 3584 -4613 3614 -4590
rect 3584 -4643 3647 -4613
rect 3617 -4658 3647 -4643
rect 3701 -4658 3731 -4569
rect 3956 -4658 3986 -4529
rect 4051 -4540 4189 -4510
rect 4051 -4570 4082 -4540
rect 4028 -4586 4082 -4570
rect 4028 -4620 4038 -4586
rect 4072 -4620 4082 -4586
rect 4028 -4636 4082 -4620
rect 4124 -4592 4190 -4582
rect 4124 -4626 4140 -4592
rect 4174 -4626 4190 -4592
rect 4124 -4636 4190 -4626
rect 4051 -4670 4081 -4636
rect 4147 -4670 4177 -4636
rect 4313 -4658 4343 -4500
rect 4396 -4570 4426 -4376
rect 4593 -4475 4623 -4460
rect 4517 -4505 4623 -4475
rect 4517 -4522 4547 -4505
rect 4481 -4538 4547 -4522
rect 4385 -4586 4439 -4570
rect 4385 -4620 4395 -4586
rect 4429 -4620 4439 -4586
rect 4481 -4572 4491 -4538
rect 4525 -4572 4547 -4538
rect 4692 -4510 4722 -4376
rect 4778 -4408 4808 -4376
rect 4764 -4424 4818 -4408
rect 4764 -4458 4774 -4424
rect 4808 -4458 4818 -4424
rect 4764 -4474 4818 -4458
rect 4692 -4522 4742 -4510
rect 4692 -4534 4755 -4522
rect 4692 -4540 4779 -4534
rect 4713 -4550 4779 -4540
rect 4713 -4552 4735 -4550
rect 4481 -4588 4547 -4572
rect 4517 -4614 4547 -4588
rect 4616 -4598 4683 -4582
rect 4385 -4636 4439 -4620
rect 4385 -4658 4415 -4636
rect 4616 -4632 4639 -4598
rect 4673 -4632 4683 -4598
rect 4616 -4648 4683 -4632
rect 4725 -4584 4735 -4552
rect 4769 -4584 4779 -4550
rect 4725 -4600 4779 -4584
rect 4862 -4560 4892 -4376
rect 4970 -4532 5000 -4376
rect 5054 -4424 5084 -4376
rect 5042 -4440 5096 -4424
rect 5042 -4474 5052 -4440
rect 5086 -4474 5096 -4440
rect 5042 -4490 5096 -4474
rect 4965 -4548 5019 -4532
rect 4862 -4576 4923 -4560
rect 4862 -4596 4879 -4576
rect 4616 -4670 4646 -4648
rect 4725 -4670 4755 -4600
rect 4821 -4610 4879 -4596
rect 4913 -4610 4923 -4576
rect 4965 -4582 4975 -4548
rect 5009 -4582 5019 -4548
rect 4965 -4598 5019 -4582
rect 4821 -4626 4923 -4610
rect 4821 -4658 4851 -4626
rect 4970 -4658 5000 -4598
rect 5061 -4658 5091 -4490
rect 5437 -4456 5467 -4420
rect 5426 -4486 5467 -4456
rect 5218 -4524 5248 -4492
rect 5426 -4524 5456 -4486
rect 5733 -4298 5763 -4272
rect 5817 -4298 5847 -4272
rect 6084 -4292 6114 -4266
rect 6176 -4292 6206 -4266
rect 6275 -4292 6305 -4266
rect 6415 -4292 6445 -4266
rect 6512 -4292 6542 -4266
rect 6709 -4292 6739 -4266
rect 6808 -4292 6838 -4266
rect 6894 -4292 6924 -4266
rect 6978 -4292 7008 -4266
rect 7086 -4292 7116 -4266
rect 7170 -4292 7200 -4266
rect 7334 -4292 7364 -4266
rect 7553 -4292 7583 -4266
rect 7650 -4292 7680 -4266
rect 5733 -4441 5763 -4426
rect 5700 -4471 5763 -4441
rect 5534 -4524 5564 -4492
rect 5700 -4524 5730 -4471
rect 5817 -4515 5847 -4426
rect 6084 -4463 6114 -4376
rect 6176 -4414 6206 -4376
rect 5147 -4540 5456 -4524
rect 5147 -4574 5175 -4540
rect 5209 -4574 5456 -4540
rect 5147 -4590 5456 -4574
rect 5505 -4540 5564 -4524
rect 5505 -4574 5515 -4540
rect 5549 -4574 5564 -4540
rect 5505 -4590 5564 -4574
rect 5676 -4540 5730 -4524
rect 5676 -4574 5686 -4540
rect 5720 -4574 5730 -4540
rect 5772 -4525 5847 -4515
rect 5772 -4559 5788 -4525
rect 5822 -4559 5847 -4525
rect 5985 -4479 6114 -4463
rect 6160 -4424 6226 -4414
rect 6160 -4458 6176 -4424
rect 6210 -4458 6226 -4424
rect 6160 -4468 6226 -4458
rect 5985 -4513 5995 -4479
rect 6029 -4493 6114 -4479
rect 6029 -4513 6102 -4493
rect 6275 -4510 6305 -4376
rect 6415 -4434 6445 -4376
rect 6415 -4450 6470 -4434
rect 6415 -4484 6425 -4450
rect 6459 -4484 6470 -4450
rect 6415 -4500 6470 -4484
rect 5985 -4529 6102 -4513
rect 5772 -4569 5847 -4559
rect 5676 -4590 5730 -4574
rect 5249 -4612 5279 -4590
rect 5426 -4613 5456 -4590
rect 5534 -4612 5564 -4590
rect 5426 -4643 5467 -4613
rect 5437 -4658 5467 -4643
rect 5700 -4613 5730 -4590
rect 5700 -4643 5763 -4613
rect 5733 -4658 5763 -4643
rect 5817 -4658 5847 -4569
rect 6072 -4658 6102 -4529
rect 6167 -4540 6305 -4510
rect 6167 -4570 6198 -4540
rect 6144 -4586 6198 -4570
rect 6144 -4620 6154 -4586
rect 6188 -4620 6198 -4586
rect 6144 -4636 6198 -4620
rect 6240 -4592 6306 -4582
rect 6240 -4626 6256 -4592
rect 6290 -4626 6306 -4592
rect 6240 -4636 6306 -4626
rect 6167 -4670 6197 -4636
rect 6263 -4670 6293 -4636
rect 6429 -4658 6459 -4500
rect 6512 -4570 6542 -4376
rect 6709 -4475 6739 -4460
rect 6633 -4505 6739 -4475
rect 6633 -4522 6663 -4505
rect 6597 -4538 6663 -4522
rect 6501 -4586 6555 -4570
rect 6501 -4620 6511 -4586
rect 6545 -4620 6555 -4586
rect 6597 -4572 6607 -4538
rect 6641 -4572 6663 -4538
rect 6808 -4510 6838 -4376
rect 6894 -4408 6924 -4376
rect 6880 -4424 6934 -4408
rect 6880 -4458 6890 -4424
rect 6924 -4458 6934 -4424
rect 6880 -4474 6934 -4458
rect 6808 -4522 6858 -4510
rect 6808 -4534 6871 -4522
rect 6808 -4540 6895 -4534
rect 6829 -4550 6895 -4540
rect 6829 -4552 6851 -4550
rect 6597 -4588 6663 -4572
rect 6633 -4614 6663 -4588
rect 6732 -4598 6799 -4582
rect 6501 -4636 6555 -4620
rect 6501 -4658 6531 -4636
rect 6732 -4632 6755 -4598
rect 6789 -4632 6799 -4598
rect 6732 -4648 6799 -4632
rect 6841 -4584 6851 -4552
rect 6885 -4584 6895 -4550
rect 6841 -4600 6895 -4584
rect 6978 -4560 7008 -4376
rect 7086 -4532 7116 -4376
rect 7170 -4424 7200 -4376
rect 7158 -4440 7212 -4424
rect 7158 -4474 7168 -4440
rect 7202 -4474 7212 -4440
rect 7158 -4490 7212 -4474
rect 7081 -4548 7135 -4532
rect 6978 -4576 7039 -4560
rect 6978 -4596 6995 -4576
rect 6732 -4670 6762 -4648
rect 6841 -4670 6871 -4600
rect 6937 -4610 6995 -4596
rect 7029 -4610 7039 -4576
rect 7081 -4582 7091 -4548
rect 7125 -4582 7135 -4548
rect 7081 -4598 7135 -4582
rect 6937 -4626 7039 -4610
rect 6937 -4658 6967 -4626
rect 7086 -4658 7116 -4598
rect 7177 -4658 7207 -4490
rect 7553 -4456 7583 -4420
rect 7542 -4486 7583 -4456
rect 7334 -4524 7364 -4492
rect 7542 -4524 7572 -4486
rect 7849 -4298 7879 -4272
rect 7933 -4298 7963 -4272
rect 8200 -4292 8230 -4266
rect 8292 -4292 8322 -4266
rect 8391 -4292 8421 -4266
rect 8531 -4292 8561 -4266
rect 8628 -4292 8658 -4266
rect 8825 -4292 8855 -4266
rect 8924 -4292 8954 -4266
rect 9010 -4292 9040 -4266
rect 9094 -4292 9124 -4266
rect 9202 -4292 9232 -4266
rect 9286 -4292 9316 -4266
rect 9450 -4292 9480 -4266
rect 9669 -4292 9699 -4266
rect 9766 -4292 9796 -4266
rect 7849 -4441 7879 -4426
rect 7816 -4471 7879 -4441
rect 7650 -4524 7680 -4492
rect 7816 -4524 7846 -4471
rect 7933 -4515 7963 -4426
rect 8200 -4463 8230 -4376
rect 8292 -4414 8322 -4376
rect 7263 -4540 7572 -4524
rect 7263 -4574 7291 -4540
rect 7325 -4574 7572 -4540
rect 7263 -4590 7572 -4574
rect 7621 -4540 7680 -4524
rect 7621 -4574 7631 -4540
rect 7665 -4574 7680 -4540
rect 7621 -4590 7680 -4574
rect 7792 -4540 7846 -4524
rect 7792 -4574 7802 -4540
rect 7836 -4574 7846 -4540
rect 7888 -4525 7963 -4515
rect 7888 -4559 7904 -4525
rect 7938 -4559 7963 -4525
rect 8101 -4479 8230 -4463
rect 8276 -4424 8342 -4414
rect 8276 -4458 8292 -4424
rect 8326 -4458 8342 -4424
rect 8276 -4468 8342 -4458
rect 8101 -4513 8111 -4479
rect 8145 -4493 8230 -4479
rect 8145 -4513 8218 -4493
rect 8391 -4510 8421 -4376
rect 8531 -4434 8561 -4376
rect 8531 -4450 8586 -4434
rect 8531 -4484 8541 -4450
rect 8575 -4484 8586 -4450
rect 8531 -4500 8586 -4484
rect 8101 -4529 8218 -4513
rect 7888 -4569 7963 -4559
rect 7792 -4590 7846 -4574
rect 7365 -4612 7395 -4590
rect 7542 -4613 7572 -4590
rect 7650 -4612 7680 -4590
rect 7542 -4643 7583 -4613
rect 7553 -4658 7583 -4643
rect 7816 -4613 7846 -4590
rect 7816 -4643 7879 -4613
rect 7849 -4658 7879 -4643
rect 7933 -4658 7963 -4569
rect 8188 -4658 8218 -4529
rect 8283 -4540 8421 -4510
rect 8283 -4570 8314 -4540
rect 8260 -4586 8314 -4570
rect 8260 -4620 8270 -4586
rect 8304 -4620 8314 -4586
rect 8260 -4636 8314 -4620
rect 8356 -4592 8422 -4582
rect 8356 -4626 8372 -4592
rect 8406 -4626 8422 -4592
rect 8356 -4636 8422 -4626
rect 8283 -4670 8313 -4636
rect 8379 -4670 8409 -4636
rect 8545 -4658 8575 -4500
rect 8628 -4570 8658 -4376
rect 8825 -4475 8855 -4460
rect 8749 -4505 8855 -4475
rect 8749 -4522 8779 -4505
rect 8713 -4538 8779 -4522
rect 8617 -4586 8671 -4570
rect 8617 -4620 8627 -4586
rect 8661 -4620 8671 -4586
rect 8713 -4572 8723 -4538
rect 8757 -4572 8779 -4538
rect 8924 -4510 8954 -4376
rect 9010 -4408 9040 -4376
rect 8996 -4424 9050 -4408
rect 8996 -4458 9006 -4424
rect 9040 -4458 9050 -4424
rect 8996 -4474 9050 -4458
rect 8924 -4522 8974 -4510
rect 8924 -4534 8987 -4522
rect 8924 -4540 9011 -4534
rect 8945 -4550 9011 -4540
rect 8945 -4552 8967 -4550
rect 8713 -4588 8779 -4572
rect 8749 -4614 8779 -4588
rect 8848 -4598 8915 -4582
rect 8617 -4636 8671 -4620
rect 8617 -4658 8647 -4636
rect 8848 -4632 8871 -4598
rect 8905 -4632 8915 -4598
rect 8848 -4648 8915 -4632
rect 8957 -4584 8967 -4552
rect 9001 -4584 9011 -4550
rect 8957 -4600 9011 -4584
rect 9094 -4560 9124 -4376
rect 9202 -4532 9232 -4376
rect 9286 -4424 9316 -4376
rect 9274 -4440 9328 -4424
rect 9274 -4474 9284 -4440
rect 9318 -4474 9328 -4440
rect 9274 -4490 9328 -4474
rect 9197 -4548 9251 -4532
rect 9094 -4576 9155 -4560
rect 9094 -4596 9111 -4576
rect 8848 -4670 8878 -4648
rect 8957 -4670 8987 -4600
rect 9053 -4610 9111 -4596
rect 9145 -4610 9155 -4576
rect 9197 -4582 9207 -4548
rect 9241 -4582 9251 -4548
rect 9197 -4598 9251 -4582
rect 9053 -4626 9155 -4610
rect 9053 -4658 9083 -4626
rect 9202 -4658 9232 -4598
rect 9293 -4658 9323 -4490
rect 9669 -4456 9699 -4420
rect 9658 -4486 9699 -4456
rect 9450 -4524 9480 -4492
rect 9658 -4524 9688 -4486
rect 9965 -4298 9995 -4272
rect 10049 -4298 10079 -4272
rect 10316 -4292 10346 -4266
rect 10408 -4292 10438 -4266
rect 10507 -4292 10537 -4266
rect 10647 -4292 10677 -4266
rect 10744 -4292 10774 -4266
rect 10941 -4292 10971 -4266
rect 11040 -4292 11070 -4266
rect 11126 -4292 11156 -4266
rect 11210 -4292 11240 -4266
rect 11318 -4292 11348 -4266
rect 11402 -4292 11432 -4266
rect 11566 -4292 11596 -4266
rect 11785 -4292 11815 -4266
rect 11882 -4292 11912 -4266
rect 9965 -4441 9995 -4426
rect 9932 -4471 9995 -4441
rect 9766 -4524 9796 -4492
rect 9932 -4524 9962 -4471
rect 10049 -4515 10079 -4426
rect 10316 -4463 10346 -4376
rect 10408 -4414 10438 -4376
rect 9379 -4540 9688 -4524
rect 9379 -4574 9407 -4540
rect 9441 -4574 9688 -4540
rect 9379 -4590 9688 -4574
rect 9737 -4540 9796 -4524
rect 9737 -4574 9747 -4540
rect 9781 -4574 9796 -4540
rect 9737 -4590 9796 -4574
rect 9908 -4540 9962 -4524
rect 9908 -4574 9918 -4540
rect 9952 -4574 9962 -4540
rect 10004 -4525 10079 -4515
rect 10004 -4559 10020 -4525
rect 10054 -4559 10079 -4525
rect 10217 -4479 10346 -4463
rect 10392 -4424 10458 -4414
rect 10392 -4458 10408 -4424
rect 10442 -4458 10458 -4424
rect 10392 -4468 10458 -4458
rect 10217 -4513 10227 -4479
rect 10261 -4493 10346 -4479
rect 10261 -4513 10334 -4493
rect 10507 -4510 10537 -4376
rect 10647 -4434 10677 -4376
rect 10647 -4450 10702 -4434
rect 10647 -4484 10657 -4450
rect 10691 -4484 10702 -4450
rect 10647 -4500 10702 -4484
rect 10217 -4529 10334 -4513
rect 10004 -4569 10079 -4559
rect 9908 -4590 9962 -4574
rect 9481 -4612 9511 -4590
rect 9658 -4613 9688 -4590
rect 9766 -4612 9796 -4590
rect 9658 -4643 9699 -4613
rect 9669 -4658 9699 -4643
rect 9932 -4613 9962 -4590
rect 9932 -4643 9995 -4613
rect 9965 -4658 9995 -4643
rect 10049 -4658 10079 -4569
rect 10304 -4658 10334 -4529
rect 10399 -4540 10537 -4510
rect 10399 -4570 10430 -4540
rect 10376 -4586 10430 -4570
rect 10376 -4620 10386 -4586
rect 10420 -4620 10430 -4586
rect 10376 -4636 10430 -4620
rect 10472 -4592 10538 -4582
rect 10472 -4626 10488 -4592
rect 10522 -4626 10538 -4592
rect 10472 -4636 10538 -4626
rect 10399 -4670 10429 -4636
rect 10495 -4670 10525 -4636
rect 10661 -4658 10691 -4500
rect 10744 -4570 10774 -4376
rect 10941 -4475 10971 -4460
rect 10865 -4505 10971 -4475
rect 10865 -4522 10895 -4505
rect 10829 -4538 10895 -4522
rect 10733 -4586 10787 -4570
rect 10733 -4620 10743 -4586
rect 10777 -4620 10787 -4586
rect 10829 -4572 10839 -4538
rect 10873 -4572 10895 -4538
rect 11040 -4510 11070 -4376
rect 11126 -4408 11156 -4376
rect 11112 -4424 11166 -4408
rect 11112 -4458 11122 -4424
rect 11156 -4458 11166 -4424
rect 11112 -4474 11166 -4458
rect 11040 -4522 11090 -4510
rect 11040 -4534 11103 -4522
rect 11040 -4540 11127 -4534
rect 11061 -4550 11127 -4540
rect 11061 -4552 11083 -4550
rect 10829 -4588 10895 -4572
rect 10865 -4614 10895 -4588
rect 10964 -4598 11031 -4582
rect 10733 -4636 10787 -4620
rect 10733 -4658 10763 -4636
rect 10964 -4632 10987 -4598
rect 11021 -4632 11031 -4598
rect 10964 -4648 11031 -4632
rect 11073 -4584 11083 -4552
rect 11117 -4584 11127 -4550
rect 11073 -4600 11127 -4584
rect 11210 -4560 11240 -4376
rect 11318 -4532 11348 -4376
rect 11402 -4424 11432 -4376
rect 11390 -4440 11444 -4424
rect 11390 -4474 11400 -4440
rect 11434 -4474 11444 -4440
rect 11390 -4490 11444 -4474
rect 11313 -4548 11367 -4532
rect 11210 -4576 11271 -4560
rect 11210 -4596 11227 -4576
rect 10964 -4670 10994 -4648
rect 11073 -4670 11103 -4600
rect 11169 -4610 11227 -4596
rect 11261 -4610 11271 -4576
rect 11313 -4582 11323 -4548
rect 11357 -4582 11367 -4548
rect 11313 -4598 11367 -4582
rect 11169 -4626 11271 -4610
rect 11169 -4658 11199 -4626
rect 11318 -4658 11348 -4598
rect 11409 -4658 11439 -4490
rect 11785 -4456 11815 -4420
rect 11774 -4486 11815 -4456
rect 11566 -4524 11596 -4492
rect 11774 -4524 11804 -4486
rect 12081 -4298 12111 -4272
rect 12165 -4298 12195 -4272
rect 12432 -4292 12462 -4266
rect 12524 -4292 12554 -4266
rect 12623 -4292 12653 -4266
rect 12763 -4292 12793 -4266
rect 12860 -4292 12890 -4266
rect 13057 -4292 13087 -4266
rect 13156 -4292 13186 -4266
rect 13242 -4292 13272 -4266
rect 13326 -4292 13356 -4266
rect 13434 -4292 13464 -4266
rect 13518 -4292 13548 -4266
rect 13682 -4292 13712 -4266
rect 13901 -4292 13931 -4266
rect 13998 -4292 14028 -4266
rect 12081 -4441 12111 -4426
rect 12048 -4471 12111 -4441
rect 11882 -4524 11912 -4492
rect 12048 -4524 12078 -4471
rect 12165 -4515 12195 -4426
rect 12432 -4463 12462 -4376
rect 12524 -4414 12554 -4376
rect 11495 -4540 11804 -4524
rect 11495 -4574 11523 -4540
rect 11557 -4574 11804 -4540
rect 11495 -4590 11804 -4574
rect 11853 -4540 11912 -4524
rect 11853 -4574 11863 -4540
rect 11897 -4574 11912 -4540
rect 11853 -4590 11912 -4574
rect 12024 -4540 12078 -4524
rect 12024 -4574 12034 -4540
rect 12068 -4574 12078 -4540
rect 12120 -4525 12195 -4515
rect 12120 -4559 12136 -4525
rect 12170 -4559 12195 -4525
rect 12333 -4479 12462 -4463
rect 12508 -4424 12574 -4414
rect 12508 -4458 12524 -4424
rect 12558 -4458 12574 -4424
rect 12508 -4468 12574 -4458
rect 12333 -4513 12343 -4479
rect 12377 -4493 12462 -4479
rect 12377 -4513 12450 -4493
rect 12623 -4510 12653 -4376
rect 12763 -4434 12793 -4376
rect 12763 -4450 12818 -4434
rect 12763 -4484 12773 -4450
rect 12807 -4484 12818 -4450
rect 12763 -4500 12818 -4484
rect 12333 -4529 12450 -4513
rect 12120 -4569 12195 -4559
rect 12024 -4590 12078 -4574
rect 11597 -4612 11627 -4590
rect 11774 -4613 11804 -4590
rect 11882 -4612 11912 -4590
rect 11774 -4643 11815 -4613
rect 11785 -4658 11815 -4643
rect 12048 -4613 12078 -4590
rect 12048 -4643 12111 -4613
rect 12081 -4658 12111 -4643
rect 12165 -4658 12195 -4569
rect 12420 -4658 12450 -4529
rect 12515 -4540 12653 -4510
rect 12515 -4570 12546 -4540
rect 12492 -4586 12546 -4570
rect 12492 -4620 12502 -4586
rect 12536 -4620 12546 -4586
rect 12492 -4636 12546 -4620
rect 12588 -4592 12654 -4582
rect 12588 -4626 12604 -4592
rect 12638 -4626 12654 -4592
rect 12588 -4636 12654 -4626
rect 12515 -4670 12545 -4636
rect 12611 -4670 12641 -4636
rect 12777 -4658 12807 -4500
rect 12860 -4570 12890 -4376
rect 13057 -4475 13087 -4460
rect 12981 -4505 13087 -4475
rect 12981 -4522 13011 -4505
rect 12945 -4538 13011 -4522
rect 12849 -4586 12903 -4570
rect 12849 -4620 12859 -4586
rect 12893 -4620 12903 -4586
rect 12945 -4572 12955 -4538
rect 12989 -4572 13011 -4538
rect 13156 -4510 13186 -4376
rect 13242 -4408 13272 -4376
rect 13228 -4424 13282 -4408
rect 13228 -4458 13238 -4424
rect 13272 -4458 13282 -4424
rect 13228 -4474 13282 -4458
rect 13156 -4522 13206 -4510
rect 13156 -4534 13219 -4522
rect 13156 -4540 13243 -4534
rect 13177 -4550 13243 -4540
rect 13177 -4552 13199 -4550
rect 12945 -4588 13011 -4572
rect 12981 -4614 13011 -4588
rect 13080 -4598 13147 -4582
rect 12849 -4636 12903 -4620
rect 12849 -4658 12879 -4636
rect 13080 -4632 13103 -4598
rect 13137 -4632 13147 -4598
rect 13080 -4648 13147 -4632
rect 13189 -4584 13199 -4552
rect 13233 -4584 13243 -4550
rect 13189 -4600 13243 -4584
rect 13326 -4560 13356 -4376
rect 13434 -4532 13464 -4376
rect 13518 -4424 13548 -4376
rect 13506 -4440 13560 -4424
rect 13506 -4474 13516 -4440
rect 13550 -4474 13560 -4440
rect 13506 -4490 13560 -4474
rect 13429 -4548 13483 -4532
rect 13326 -4576 13387 -4560
rect 13326 -4596 13343 -4576
rect 13080 -4670 13110 -4648
rect 13189 -4670 13219 -4600
rect 13285 -4610 13343 -4596
rect 13377 -4610 13387 -4576
rect 13429 -4582 13439 -4548
rect 13473 -4582 13483 -4548
rect 13429 -4598 13483 -4582
rect 13285 -4626 13387 -4610
rect 13285 -4658 13315 -4626
rect 13434 -4658 13464 -4598
rect 13525 -4658 13555 -4490
rect 13901 -4456 13931 -4420
rect 13890 -4486 13931 -4456
rect 13682 -4524 13712 -4492
rect 13890 -4524 13920 -4486
rect 14197 -4298 14227 -4272
rect 14281 -4298 14311 -4272
rect 14548 -4292 14578 -4266
rect 14640 -4292 14670 -4266
rect 14739 -4292 14769 -4266
rect 14879 -4292 14909 -4266
rect 14976 -4292 15006 -4266
rect 15173 -4292 15203 -4266
rect 15272 -4292 15302 -4266
rect 15358 -4292 15388 -4266
rect 15442 -4292 15472 -4266
rect 15550 -4292 15580 -4266
rect 15634 -4292 15664 -4266
rect 15798 -4292 15828 -4266
rect 16017 -4292 16047 -4266
rect 16114 -4292 16144 -4266
rect 14197 -4441 14227 -4426
rect 14164 -4471 14227 -4441
rect 13998 -4524 14028 -4492
rect 14164 -4524 14194 -4471
rect 14281 -4515 14311 -4426
rect 14548 -4463 14578 -4376
rect 14640 -4414 14670 -4376
rect 13611 -4540 13920 -4524
rect 13611 -4574 13639 -4540
rect 13673 -4574 13920 -4540
rect 13611 -4590 13920 -4574
rect 13969 -4540 14028 -4524
rect 13969 -4574 13979 -4540
rect 14013 -4574 14028 -4540
rect 13969 -4590 14028 -4574
rect 14140 -4540 14194 -4524
rect 14140 -4574 14150 -4540
rect 14184 -4574 14194 -4540
rect 14236 -4525 14311 -4515
rect 14236 -4559 14252 -4525
rect 14286 -4559 14311 -4525
rect 14449 -4479 14578 -4463
rect 14624 -4424 14690 -4414
rect 14624 -4458 14640 -4424
rect 14674 -4458 14690 -4424
rect 14624 -4468 14690 -4458
rect 14449 -4513 14459 -4479
rect 14493 -4493 14578 -4479
rect 14493 -4513 14566 -4493
rect 14739 -4510 14769 -4376
rect 14879 -4434 14909 -4376
rect 14879 -4450 14934 -4434
rect 14879 -4484 14889 -4450
rect 14923 -4484 14934 -4450
rect 14879 -4500 14934 -4484
rect 14449 -4529 14566 -4513
rect 14236 -4569 14311 -4559
rect 14140 -4590 14194 -4574
rect 13713 -4612 13743 -4590
rect 13890 -4613 13920 -4590
rect 13998 -4612 14028 -4590
rect 13890 -4643 13931 -4613
rect 13901 -4658 13931 -4643
rect 14164 -4613 14194 -4590
rect 14164 -4643 14227 -4613
rect 14197 -4658 14227 -4643
rect 14281 -4658 14311 -4569
rect 14536 -4658 14566 -4529
rect 14631 -4540 14769 -4510
rect 14631 -4570 14662 -4540
rect 14608 -4586 14662 -4570
rect 14608 -4620 14618 -4586
rect 14652 -4620 14662 -4586
rect 14608 -4636 14662 -4620
rect 14704 -4592 14770 -4582
rect 14704 -4626 14720 -4592
rect 14754 -4626 14770 -4592
rect 14704 -4636 14770 -4626
rect 14631 -4670 14661 -4636
rect 14727 -4670 14757 -4636
rect 14893 -4658 14923 -4500
rect 14976 -4570 15006 -4376
rect 15173 -4475 15203 -4460
rect 15097 -4505 15203 -4475
rect 15097 -4522 15127 -4505
rect 15061 -4538 15127 -4522
rect 14965 -4586 15019 -4570
rect 14965 -4620 14975 -4586
rect 15009 -4620 15019 -4586
rect 15061 -4572 15071 -4538
rect 15105 -4572 15127 -4538
rect 15272 -4510 15302 -4376
rect 15358 -4408 15388 -4376
rect 15344 -4424 15398 -4408
rect 15344 -4458 15354 -4424
rect 15388 -4458 15398 -4424
rect 15344 -4474 15398 -4458
rect 15272 -4522 15322 -4510
rect 15272 -4534 15335 -4522
rect 15272 -4540 15359 -4534
rect 15293 -4550 15359 -4540
rect 15293 -4552 15315 -4550
rect 15061 -4588 15127 -4572
rect 15097 -4614 15127 -4588
rect 15196 -4598 15263 -4582
rect 14965 -4636 15019 -4620
rect 14965 -4658 14995 -4636
rect 15196 -4632 15219 -4598
rect 15253 -4632 15263 -4598
rect 15196 -4648 15263 -4632
rect 15305 -4584 15315 -4552
rect 15349 -4584 15359 -4550
rect 15305 -4600 15359 -4584
rect 15442 -4560 15472 -4376
rect 15550 -4532 15580 -4376
rect 15634 -4424 15664 -4376
rect 15622 -4440 15676 -4424
rect 15622 -4474 15632 -4440
rect 15666 -4474 15676 -4440
rect 15622 -4490 15676 -4474
rect 15545 -4548 15599 -4532
rect 15442 -4576 15503 -4560
rect 15442 -4596 15459 -4576
rect 15196 -4670 15226 -4648
rect 15305 -4670 15335 -4600
rect 15401 -4610 15459 -4596
rect 15493 -4610 15503 -4576
rect 15545 -4582 15555 -4548
rect 15589 -4582 15599 -4548
rect 15545 -4598 15599 -4582
rect 15401 -4626 15503 -4610
rect 15401 -4658 15431 -4626
rect 15550 -4658 15580 -4598
rect 15641 -4658 15671 -4490
rect 16017 -4456 16047 -4420
rect 16006 -4486 16047 -4456
rect 15798 -4524 15828 -4492
rect 16006 -4524 16036 -4486
rect 16313 -4298 16343 -4272
rect 16397 -4298 16427 -4272
rect 16664 -4292 16694 -4266
rect 16756 -4292 16786 -4266
rect 16855 -4292 16885 -4266
rect 16995 -4292 17025 -4266
rect 17092 -4292 17122 -4266
rect 17289 -4292 17319 -4266
rect 17388 -4292 17418 -4266
rect 17474 -4292 17504 -4266
rect 17558 -4292 17588 -4266
rect 17666 -4292 17696 -4266
rect 17750 -4292 17780 -4266
rect 17914 -4292 17944 -4266
rect 18133 -4292 18163 -4266
rect 18230 -4292 18260 -4266
rect 16313 -4441 16343 -4426
rect 16280 -4471 16343 -4441
rect 16114 -4524 16144 -4492
rect 16280 -4524 16310 -4471
rect 16397 -4515 16427 -4426
rect 16664 -4463 16694 -4376
rect 16756 -4414 16786 -4376
rect 15727 -4540 16036 -4524
rect 15727 -4574 15755 -4540
rect 15789 -4574 16036 -4540
rect 15727 -4590 16036 -4574
rect 16085 -4540 16144 -4524
rect 16085 -4574 16095 -4540
rect 16129 -4574 16144 -4540
rect 16085 -4590 16144 -4574
rect 16256 -4540 16310 -4524
rect 16256 -4574 16266 -4540
rect 16300 -4574 16310 -4540
rect 16352 -4525 16427 -4515
rect 16352 -4559 16368 -4525
rect 16402 -4559 16427 -4525
rect 16565 -4479 16694 -4463
rect 16740 -4424 16806 -4414
rect 16740 -4458 16756 -4424
rect 16790 -4458 16806 -4424
rect 16740 -4468 16806 -4458
rect 16565 -4513 16575 -4479
rect 16609 -4493 16694 -4479
rect 16609 -4513 16682 -4493
rect 16855 -4510 16885 -4376
rect 16995 -4434 17025 -4376
rect 16995 -4450 17050 -4434
rect 16995 -4484 17005 -4450
rect 17039 -4484 17050 -4450
rect 16995 -4500 17050 -4484
rect 16565 -4529 16682 -4513
rect 16352 -4569 16427 -4559
rect 16256 -4590 16310 -4574
rect 15829 -4612 15859 -4590
rect 16006 -4613 16036 -4590
rect 16114 -4612 16144 -4590
rect 16006 -4643 16047 -4613
rect 16017 -4658 16047 -4643
rect 16280 -4613 16310 -4590
rect 16280 -4643 16343 -4613
rect 16313 -4658 16343 -4643
rect 16397 -4658 16427 -4569
rect 16652 -4658 16682 -4529
rect 16747 -4540 16885 -4510
rect 16747 -4570 16778 -4540
rect 16724 -4586 16778 -4570
rect 16724 -4620 16734 -4586
rect 16768 -4620 16778 -4586
rect 16724 -4636 16778 -4620
rect 16820 -4592 16886 -4582
rect 16820 -4626 16836 -4592
rect 16870 -4626 16886 -4592
rect 16820 -4636 16886 -4626
rect 16747 -4670 16777 -4636
rect 16843 -4670 16873 -4636
rect 17009 -4658 17039 -4500
rect 17092 -4570 17122 -4376
rect 17289 -4475 17319 -4460
rect 17213 -4505 17319 -4475
rect 17213 -4522 17243 -4505
rect 17177 -4538 17243 -4522
rect 17081 -4586 17135 -4570
rect 17081 -4620 17091 -4586
rect 17125 -4620 17135 -4586
rect 17177 -4572 17187 -4538
rect 17221 -4572 17243 -4538
rect 17388 -4510 17418 -4376
rect 17474 -4408 17504 -4376
rect 17460 -4424 17514 -4408
rect 17460 -4458 17470 -4424
rect 17504 -4458 17514 -4424
rect 17460 -4474 17514 -4458
rect 17388 -4522 17438 -4510
rect 17388 -4534 17451 -4522
rect 17388 -4540 17475 -4534
rect 17409 -4550 17475 -4540
rect 17409 -4552 17431 -4550
rect 17177 -4588 17243 -4572
rect 17213 -4614 17243 -4588
rect 17312 -4598 17379 -4582
rect 17081 -4636 17135 -4620
rect 17081 -4658 17111 -4636
rect 17312 -4632 17335 -4598
rect 17369 -4632 17379 -4598
rect 17312 -4648 17379 -4632
rect 17421 -4584 17431 -4552
rect 17465 -4584 17475 -4550
rect 17421 -4600 17475 -4584
rect 17558 -4560 17588 -4376
rect 17666 -4532 17696 -4376
rect 17750 -4424 17780 -4376
rect 17738 -4440 17792 -4424
rect 17738 -4474 17748 -4440
rect 17782 -4474 17792 -4440
rect 17738 -4490 17792 -4474
rect 17661 -4548 17715 -4532
rect 17558 -4576 17619 -4560
rect 17558 -4596 17575 -4576
rect 17312 -4670 17342 -4648
rect 17421 -4670 17451 -4600
rect 17517 -4610 17575 -4596
rect 17609 -4610 17619 -4576
rect 17661 -4582 17671 -4548
rect 17705 -4582 17715 -4548
rect 17661 -4598 17715 -4582
rect 17517 -4626 17619 -4610
rect 17517 -4658 17547 -4626
rect 17666 -4658 17696 -4598
rect 17757 -4658 17787 -4490
rect 18133 -4456 18163 -4420
rect 18122 -4486 18163 -4456
rect 17914 -4524 17944 -4492
rect 18122 -4524 18152 -4486
rect 18429 -4298 18459 -4272
rect 18513 -4298 18543 -4272
rect 18780 -4292 18810 -4266
rect 18872 -4292 18902 -4266
rect 18971 -4292 19001 -4266
rect 19111 -4292 19141 -4266
rect 19208 -4292 19238 -4266
rect 19405 -4292 19435 -4266
rect 19504 -4292 19534 -4266
rect 19590 -4292 19620 -4266
rect 19674 -4292 19704 -4266
rect 19782 -4292 19812 -4266
rect 19866 -4292 19896 -4266
rect 20030 -4292 20060 -4266
rect 20249 -4292 20279 -4266
rect 20346 -4292 20376 -4266
rect 18429 -4441 18459 -4426
rect 18396 -4471 18459 -4441
rect 18230 -4524 18260 -4492
rect 18396 -4524 18426 -4471
rect 18513 -4515 18543 -4426
rect 18780 -4463 18810 -4376
rect 18872 -4414 18902 -4376
rect 17843 -4540 18152 -4524
rect 17843 -4574 17871 -4540
rect 17905 -4574 18152 -4540
rect 17843 -4590 18152 -4574
rect 18201 -4540 18260 -4524
rect 18201 -4574 18211 -4540
rect 18245 -4574 18260 -4540
rect 18201 -4590 18260 -4574
rect 18372 -4540 18426 -4524
rect 18372 -4574 18382 -4540
rect 18416 -4574 18426 -4540
rect 18468 -4525 18543 -4515
rect 18468 -4559 18484 -4525
rect 18518 -4559 18543 -4525
rect 18681 -4479 18810 -4463
rect 18856 -4424 18922 -4414
rect 18856 -4458 18872 -4424
rect 18906 -4458 18922 -4424
rect 18856 -4468 18922 -4458
rect 18681 -4513 18691 -4479
rect 18725 -4493 18810 -4479
rect 18725 -4513 18798 -4493
rect 18971 -4510 19001 -4376
rect 19111 -4434 19141 -4376
rect 19111 -4450 19166 -4434
rect 19111 -4484 19121 -4450
rect 19155 -4484 19166 -4450
rect 19111 -4500 19166 -4484
rect 18681 -4529 18798 -4513
rect 18468 -4569 18543 -4559
rect 18372 -4590 18426 -4574
rect 17945 -4612 17975 -4590
rect 18122 -4613 18152 -4590
rect 18230 -4612 18260 -4590
rect 18122 -4643 18163 -4613
rect 18133 -4658 18163 -4643
rect 18396 -4613 18426 -4590
rect 18396 -4643 18459 -4613
rect 18429 -4658 18459 -4643
rect 18513 -4658 18543 -4569
rect 18768 -4658 18798 -4529
rect 18863 -4540 19001 -4510
rect 18863 -4570 18894 -4540
rect 18840 -4586 18894 -4570
rect 18840 -4620 18850 -4586
rect 18884 -4620 18894 -4586
rect 18840 -4636 18894 -4620
rect 18936 -4592 19002 -4582
rect 18936 -4626 18952 -4592
rect 18986 -4626 19002 -4592
rect 18936 -4636 19002 -4626
rect 18863 -4670 18893 -4636
rect 18959 -4670 18989 -4636
rect 19125 -4658 19155 -4500
rect 19208 -4570 19238 -4376
rect 19405 -4475 19435 -4460
rect 19329 -4505 19435 -4475
rect 19329 -4522 19359 -4505
rect 19293 -4538 19359 -4522
rect 19197 -4586 19251 -4570
rect 19197 -4620 19207 -4586
rect 19241 -4620 19251 -4586
rect 19293 -4572 19303 -4538
rect 19337 -4572 19359 -4538
rect 19504 -4510 19534 -4376
rect 19590 -4408 19620 -4376
rect 19576 -4424 19630 -4408
rect 19576 -4458 19586 -4424
rect 19620 -4458 19630 -4424
rect 19576 -4474 19630 -4458
rect 19504 -4522 19554 -4510
rect 19504 -4534 19567 -4522
rect 19504 -4540 19591 -4534
rect 19525 -4550 19591 -4540
rect 19525 -4552 19547 -4550
rect 19293 -4588 19359 -4572
rect 19329 -4614 19359 -4588
rect 19428 -4598 19495 -4582
rect 19197 -4636 19251 -4620
rect 19197 -4658 19227 -4636
rect 19428 -4632 19451 -4598
rect 19485 -4632 19495 -4598
rect 19428 -4648 19495 -4632
rect 19537 -4584 19547 -4552
rect 19581 -4584 19591 -4550
rect 19537 -4600 19591 -4584
rect 19674 -4560 19704 -4376
rect 19782 -4532 19812 -4376
rect 19866 -4424 19896 -4376
rect 19854 -4440 19908 -4424
rect 19854 -4474 19864 -4440
rect 19898 -4474 19908 -4440
rect 19854 -4490 19908 -4474
rect 19777 -4548 19831 -4532
rect 19674 -4576 19735 -4560
rect 19674 -4596 19691 -4576
rect 19428 -4670 19458 -4648
rect 19537 -4670 19567 -4600
rect 19633 -4610 19691 -4596
rect 19725 -4610 19735 -4576
rect 19777 -4582 19787 -4548
rect 19821 -4582 19831 -4548
rect 19777 -4598 19831 -4582
rect 19633 -4626 19735 -4610
rect 19633 -4658 19663 -4626
rect 19782 -4658 19812 -4598
rect 19873 -4658 19903 -4490
rect 20249 -4456 20279 -4420
rect 20238 -4486 20279 -4456
rect 20030 -4524 20060 -4492
rect 20238 -4524 20268 -4486
rect 20545 -4298 20575 -4272
rect 20629 -4298 20659 -4272
rect 20896 -4292 20926 -4266
rect 20988 -4292 21018 -4266
rect 21087 -4292 21117 -4266
rect 21227 -4292 21257 -4266
rect 21324 -4292 21354 -4266
rect 21521 -4292 21551 -4266
rect 21620 -4292 21650 -4266
rect 21706 -4292 21736 -4266
rect 21790 -4292 21820 -4266
rect 21898 -4292 21928 -4266
rect 21982 -4292 22012 -4266
rect 22146 -4292 22176 -4266
rect 22365 -4292 22395 -4266
rect 22462 -4292 22492 -4266
rect 20545 -4441 20575 -4426
rect 20512 -4471 20575 -4441
rect 20346 -4524 20376 -4492
rect 20512 -4524 20542 -4471
rect 20629 -4515 20659 -4426
rect 20896 -4463 20926 -4376
rect 20988 -4414 21018 -4376
rect 19959 -4540 20268 -4524
rect 19959 -4574 19987 -4540
rect 20021 -4574 20268 -4540
rect 19959 -4590 20268 -4574
rect 20317 -4540 20376 -4524
rect 20317 -4574 20327 -4540
rect 20361 -4574 20376 -4540
rect 20317 -4590 20376 -4574
rect 20488 -4540 20542 -4524
rect 20488 -4574 20498 -4540
rect 20532 -4574 20542 -4540
rect 20584 -4525 20659 -4515
rect 20584 -4559 20600 -4525
rect 20634 -4559 20659 -4525
rect 20797 -4479 20926 -4463
rect 20972 -4424 21038 -4414
rect 20972 -4458 20988 -4424
rect 21022 -4458 21038 -4424
rect 20972 -4468 21038 -4458
rect 20797 -4513 20807 -4479
rect 20841 -4493 20926 -4479
rect 20841 -4513 20914 -4493
rect 21087 -4510 21117 -4376
rect 21227 -4434 21257 -4376
rect 21227 -4450 21282 -4434
rect 21227 -4484 21237 -4450
rect 21271 -4484 21282 -4450
rect 21227 -4500 21282 -4484
rect 20797 -4529 20914 -4513
rect 20584 -4569 20659 -4559
rect 20488 -4590 20542 -4574
rect 20061 -4612 20091 -4590
rect 20238 -4613 20268 -4590
rect 20346 -4612 20376 -4590
rect 20238 -4643 20279 -4613
rect 20249 -4658 20279 -4643
rect 20512 -4613 20542 -4590
rect 20512 -4643 20575 -4613
rect 20545 -4658 20575 -4643
rect 20629 -4658 20659 -4569
rect 20884 -4658 20914 -4529
rect 20979 -4540 21117 -4510
rect 20979 -4570 21010 -4540
rect 20956 -4586 21010 -4570
rect 20956 -4620 20966 -4586
rect 21000 -4620 21010 -4586
rect 20956 -4636 21010 -4620
rect 21052 -4592 21118 -4582
rect 21052 -4626 21068 -4592
rect 21102 -4626 21118 -4592
rect 21052 -4636 21118 -4626
rect 20979 -4670 21009 -4636
rect 21075 -4670 21105 -4636
rect 21241 -4658 21271 -4500
rect 21324 -4570 21354 -4376
rect 21521 -4475 21551 -4460
rect 21445 -4505 21551 -4475
rect 21445 -4522 21475 -4505
rect 21409 -4538 21475 -4522
rect 21313 -4586 21367 -4570
rect 21313 -4620 21323 -4586
rect 21357 -4620 21367 -4586
rect 21409 -4572 21419 -4538
rect 21453 -4572 21475 -4538
rect 21620 -4510 21650 -4376
rect 21706 -4408 21736 -4376
rect 21692 -4424 21746 -4408
rect 21692 -4458 21702 -4424
rect 21736 -4458 21746 -4424
rect 21692 -4474 21746 -4458
rect 21620 -4522 21670 -4510
rect 21620 -4534 21683 -4522
rect 21620 -4540 21707 -4534
rect 21641 -4550 21707 -4540
rect 21641 -4552 21663 -4550
rect 21409 -4588 21475 -4572
rect 21445 -4614 21475 -4588
rect 21544 -4598 21611 -4582
rect 21313 -4636 21367 -4620
rect 21313 -4658 21343 -4636
rect 21544 -4632 21567 -4598
rect 21601 -4632 21611 -4598
rect 21544 -4648 21611 -4632
rect 21653 -4584 21663 -4552
rect 21697 -4584 21707 -4550
rect 21653 -4600 21707 -4584
rect 21790 -4560 21820 -4376
rect 21898 -4532 21928 -4376
rect 21982 -4424 22012 -4376
rect 21970 -4440 22024 -4424
rect 21970 -4474 21980 -4440
rect 22014 -4474 22024 -4440
rect 21970 -4490 22024 -4474
rect 21893 -4548 21947 -4532
rect 21790 -4576 21851 -4560
rect 21790 -4596 21807 -4576
rect 21544 -4670 21574 -4648
rect 21653 -4670 21683 -4600
rect 21749 -4610 21807 -4596
rect 21841 -4610 21851 -4576
rect 21893 -4582 21903 -4548
rect 21937 -4582 21947 -4548
rect 21893 -4598 21947 -4582
rect 21749 -4626 21851 -4610
rect 21749 -4658 21779 -4626
rect 21898 -4658 21928 -4598
rect 21989 -4658 22019 -4490
rect 22365 -4456 22395 -4420
rect 22354 -4486 22395 -4456
rect 22146 -4524 22176 -4492
rect 22354 -4524 22384 -4486
rect 22661 -4298 22691 -4272
rect 22745 -4298 22775 -4272
rect 23012 -4292 23042 -4266
rect 23104 -4292 23134 -4266
rect 23203 -4292 23233 -4266
rect 23343 -4292 23373 -4266
rect 23440 -4292 23470 -4266
rect 23637 -4292 23667 -4266
rect 23736 -4292 23766 -4266
rect 23822 -4292 23852 -4266
rect 23906 -4292 23936 -4266
rect 24014 -4292 24044 -4266
rect 24098 -4292 24128 -4266
rect 24262 -4292 24292 -4266
rect 24481 -4292 24511 -4266
rect 24578 -4292 24608 -4266
rect 22661 -4441 22691 -4426
rect 22628 -4471 22691 -4441
rect 22462 -4524 22492 -4492
rect 22628 -4524 22658 -4471
rect 22745 -4515 22775 -4426
rect 23012 -4463 23042 -4376
rect 23104 -4414 23134 -4376
rect 22075 -4540 22384 -4524
rect 22075 -4574 22103 -4540
rect 22137 -4574 22384 -4540
rect 22075 -4590 22384 -4574
rect 22433 -4540 22492 -4524
rect 22433 -4574 22443 -4540
rect 22477 -4574 22492 -4540
rect 22433 -4590 22492 -4574
rect 22604 -4540 22658 -4524
rect 22604 -4574 22614 -4540
rect 22648 -4574 22658 -4540
rect 22700 -4525 22775 -4515
rect 22700 -4559 22716 -4525
rect 22750 -4559 22775 -4525
rect 22913 -4479 23042 -4463
rect 23088 -4424 23154 -4414
rect 23088 -4458 23104 -4424
rect 23138 -4458 23154 -4424
rect 23088 -4468 23154 -4458
rect 22913 -4513 22923 -4479
rect 22957 -4493 23042 -4479
rect 22957 -4513 23030 -4493
rect 23203 -4510 23233 -4376
rect 23343 -4434 23373 -4376
rect 23343 -4450 23398 -4434
rect 23343 -4484 23353 -4450
rect 23387 -4484 23398 -4450
rect 23343 -4500 23398 -4484
rect 22913 -4529 23030 -4513
rect 22700 -4569 22775 -4559
rect 22604 -4590 22658 -4574
rect 22177 -4612 22207 -4590
rect 22354 -4613 22384 -4590
rect 22462 -4612 22492 -4590
rect 22354 -4643 22395 -4613
rect 22365 -4658 22395 -4643
rect 22628 -4613 22658 -4590
rect 22628 -4643 22691 -4613
rect 22661 -4658 22691 -4643
rect 22745 -4658 22775 -4569
rect 23000 -4658 23030 -4529
rect 23095 -4540 23233 -4510
rect 23095 -4570 23126 -4540
rect 23072 -4586 23126 -4570
rect 23072 -4620 23082 -4586
rect 23116 -4620 23126 -4586
rect 23072 -4636 23126 -4620
rect 23168 -4592 23234 -4582
rect 23168 -4626 23184 -4592
rect 23218 -4626 23234 -4592
rect 23168 -4636 23234 -4626
rect 23095 -4670 23125 -4636
rect 23191 -4670 23221 -4636
rect 23357 -4658 23387 -4500
rect 23440 -4570 23470 -4376
rect 23637 -4475 23667 -4460
rect 23561 -4505 23667 -4475
rect 23561 -4522 23591 -4505
rect 23525 -4538 23591 -4522
rect 23429 -4586 23483 -4570
rect 23429 -4620 23439 -4586
rect 23473 -4620 23483 -4586
rect 23525 -4572 23535 -4538
rect 23569 -4572 23591 -4538
rect 23736 -4510 23766 -4376
rect 23822 -4408 23852 -4376
rect 23808 -4424 23862 -4408
rect 23808 -4458 23818 -4424
rect 23852 -4458 23862 -4424
rect 23808 -4474 23862 -4458
rect 23736 -4522 23786 -4510
rect 23736 -4534 23799 -4522
rect 23736 -4540 23823 -4534
rect 23757 -4550 23823 -4540
rect 23757 -4552 23779 -4550
rect 23525 -4588 23591 -4572
rect 23561 -4614 23591 -4588
rect 23660 -4598 23727 -4582
rect 23429 -4636 23483 -4620
rect 23429 -4658 23459 -4636
rect 23660 -4632 23683 -4598
rect 23717 -4632 23727 -4598
rect 23660 -4648 23727 -4632
rect 23769 -4584 23779 -4552
rect 23813 -4584 23823 -4550
rect 23769 -4600 23823 -4584
rect 23906 -4560 23936 -4376
rect 24014 -4532 24044 -4376
rect 24098 -4424 24128 -4376
rect 24086 -4440 24140 -4424
rect 24086 -4474 24096 -4440
rect 24130 -4474 24140 -4440
rect 24086 -4490 24140 -4474
rect 24009 -4548 24063 -4532
rect 23906 -4576 23967 -4560
rect 23906 -4596 23923 -4576
rect 23660 -4670 23690 -4648
rect 23769 -4670 23799 -4600
rect 23865 -4610 23923 -4596
rect 23957 -4610 23967 -4576
rect 24009 -4582 24019 -4548
rect 24053 -4582 24063 -4548
rect 24009 -4598 24063 -4582
rect 23865 -4626 23967 -4610
rect 23865 -4658 23895 -4626
rect 24014 -4658 24044 -4598
rect 24105 -4658 24135 -4490
rect 24481 -4456 24511 -4420
rect 24470 -4486 24511 -4456
rect 24262 -4524 24292 -4492
rect 24470 -4524 24500 -4486
rect 24777 -4298 24807 -4272
rect 24861 -4298 24891 -4272
rect 25128 -4292 25158 -4266
rect 25220 -4292 25250 -4266
rect 25319 -4292 25349 -4266
rect 25459 -4292 25489 -4266
rect 25556 -4292 25586 -4266
rect 25753 -4292 25783 -4266
rect 25852 -4292 25882 -4266
rect 25938 -4292 25968 -4266
rect 26022 -4292 26052 -4266
rect 26130 -4292 26160 -4266
rect 26214 -4292 26244 -4266
rect 26378 -4292 26408 -4266
rect 26597 -4292 26627 -4266
rect 26694 -4292 26724 -4266
rect 24777 -4441 24807 -4426
rect 24744 -4471 24807 -4441
rect 24578 -4524 24608 -4492
rect 24744 -4524 24774 -4471
rect 24861 -4515 24891 -4426
rect 25128 -4463 25158 -4376
rect 25220 -4414 25250 -4376
rect 24191 -4540 24500 -4524
rect 24191 -4574 24219 -4540
rect 24253 -4574 24500 -4540
rect 24191 -4590 24500 -4574
rect 24549 -4540 24608 -4524
rect 24549 -4574 24559 -4540
rect 24593 -4574 24608 -4540
rect 24549 -4590 24608 -4574
rect 24720 -4540 24774 -4524
rect 24720 -4574 24730 -4540
rect 24764 -4574 24774 -4540
rect 24816 -4525 24891 -4515
rect 24816 -4559 24832 -4525
rect 24866 -4559 24891 -4525
rect 25029 -4479 25158 -4463
rect 25204 -4424 25270 -4414
rect 25204 -4458 25220 -4424
rect 25254 -4458 25270 -4424
rect 25204 -4468 25270 -4458
rect 25029 -4513 25039 -4479
rect 25073 -4493 25158 -4479
rect 25073 -4513 25146 -4493
rect 25319 -4510 25349 -4376
rect 25459 -4434 25489 -4376
rect 25459 -4450 25514 -4434
rect 25459 -4484 25469 -4450
rect 25503 -4484 25514 -4450
rect 25459 -4500 25514 -4484
rect 25029 -4529 25146 -4513
rect 24816 -4569 24891 -4559
rect 24720 -4590 24774 -4574
rect 24293 -4612 24323 -4590
rect 24470 -4613 24500 -4590
rect 24578 -4612 24608 -4590
rect 24470 -4643 24511 -4613
rect 24481 -4658 24511 -4643
rect 24744 -4613 24774 -4590
rect 24744 -4643 24807 -4613
rect 24777 -4658 24807 -4643
rect 24861 -4658 24891 -4569
rect 25116 -4658 25146 -4529
rect 25211 -4540 25349 -4510
rect 25211 -4570 25242 -4540
rect 25188 -4586 25242 -4570
rect 25188 -4620 25198 -4586
rect 25232 -4620 25242 -4586
rect 25188 -4636 25242 -4620
rect 25284 -4592 25350 -4582
rect 25284 -4626 25300 -4592
rect 25334 -4626 25350 -4592
rect 25284 -4636 25350 -4626
rect 25211 -4670 25241 -4636
rect 25307 -4670 25337 -4636
rect 25473 -4658 25503 -4500
rect 25556 -4570 25586 -4376
rect 25753 -4475 25783 -4460
rect 25677 -4505 25783 -4475
rect 25677 -4522 25707 -4505
rect 25641 -4538 25707 -4522
rect 25545 -4586 25599 -4570
rect 25545 -4620 25555 -4586
rect 25589 -4620 25599 -4586
rect 25641 -4572 25651 -4538
rect 25685 -4572 25707 -4538
rect 25852 -4510 25882 -4376
rect 25938 -4408 25968 -4376
rect 25924 -4424 25978 -4408
rect 25924 -4458 25934 -4424
rect 25968 -4458 25978 -4424
rect 25924 -4474 25978 -4458
rect 25852 -4522 25902 -4510
rect 25852 -4534 25915 -4522
rect 25852 -4540 25939 -4534
rect 25873 -4550 25939 -4540
rect 25873 -4552 25895 -4550
rect 25641 -4588 25707 -4572
rect 25677 -4614 25707 -4588
rect 25776 -4598 25843 -4582
rect 25545 -4636 25599 -4620
rect 25545 -4658 25575 -4636
rect 25776 -4632 25799 -4598
rect 25833 -4632 25843 -4598
rect 25776 -4648 25843 -4632
rect 25885 -4584 25895 -4552
rect 25929 -4584 25939 -4550
rect 25885 -4600 25939 -4584
rect 26022 -4560 26052 -4376
rect 26130 -4532 26160 -4376
rect 26214 -4424 26244 -4376
rect 26202 -4440 26256 -4424
rect 26202 -4474 26212 -4440
rect 26246 -4474 26256 -4440
rect 26202 -4490 26256 -4474
rect 26125 -4548 26179 -4532
rect 26022 -4576 26083 -4560
rect 26022 -4596 26039 -4576
rect 25776 -4670 25806 -4648
rect 25885 -4670 25915 -4600
rect 25981 -4610 26039 -4596
rect 26073 -4610 26083 -4576
rect 26125 -4582 26135 -4548
rect 26169 -4582 26179 -4548
rect 26125 -4598 26179 -4582
rect 25981 -4626 26083 -4610
rect 25981 -4658 26011 -4626
rect 26130 -4658 26160 -4598
rect 26221 -4658 26251 -4490
rect 26597 -4456 26627 -4420
rect 26586 -4486 26627 -4456
rect 26378 -4524 26408 -4492
rect 26586 -4524 26616 -4486
rect 26893 -4298 26923 -4272
rect 26977 -4298 27007 -4272
rect 27244 -4292 27274 -4266
rect 27336 -4292 27366 -4266
rect 27435 -4292 27465 -4266
rect 27575 -4292 27605 -4266
rect 27672 -4292 27702 -4266
rect 27869 -4292 27899 -4266
rect 27968 -4292 27998 -4266
rect 28054 -4292 28084 -4266
rect 28138 -4292 28168 -4266
rect 28246 -4292 28276 -4266
rect 28330 -4292 28360 -4266
rect 28494 -4292 28524 -4266
rect 28713 -4292 28743 -4266
rect 28810 -4292 28840 -4266
rect 26893 -4441 26923 -4426
rect 26860 -4471 26923 -4441
rect 26694 -4524 26724 -4492
rect 26860 -4524 26890 -4471
rect 26977 -4515 27007 -4426
rect 27244 -4463 27274 -4376
rect 27336 -4414 27366 -4376
rect 26307 -4540 26616 -4524
rect 26307 -4574 26335 -4540
rect 26369 -4574 26616 -4540
rect 26307 -4590 26616 -4574
rect 26665 -4540 26724 -4524
rect 26665 -4574 26675 -4540
rect 26709 -4574 26724 -4540
rect 26665 -4590 26724 -4574
rect 26836 -4540 26890 -4524
rect 26836 -4574 26846 -4540
rect 26880 -4574 26890 -4540
rect 26932 -4525 27007 -4515
rect 26932 -4559 26948 -4525
rect 26982 -4559 27007 -4525
rect 27145 -4479 27274 -4463
rect 27320 -4424 27386 -4414
rect 27320 -4458 27336 -4424
rect 27370 -4458 27386 -4424
rect 27320 -4468 27386 -4458
rect 27145 -4513 27155 -4479
rect 27189 -4493 27274 -4479
rect 27189 -4513 27262 -4493
rect 27435 -4510 27465 -4376
rect 27575 -4434 27605 -4376
rect 27575 -4450 27630 -4434
rect 27575 -4484 27585 -4450
rect 27619 -4484 27630 -4450
rect 27575 -4500 27630 -4484
rect 27145 -4529 27262 -4513
rect 26932 -4569 27007 -4559
rect 26836 -4590 26890 -4574
rect 26409 -4612 26439 -4590
rect 26586 -4613 26616 -4590
rect 26694 -4612 26724 -4590
rect 26586 -4643 26627 -4613
rect 26597 -4658 26627 -4643
rect 26860 -4613 26890 -4590
rect 26860 -4643 26923 -4613
rect 26893 -4658 26923 -4643
rect 26977 -4658 27007 -4569
rect 27232 -4658 27262 -4529
rect 27327 -4540 27465 -4510
rect 27327 -4570 27358 -4540
rect 27304 -4586 27358 -4570
rect 27304 -4620 27314 -4586
rect 27348 -4620 27358 -4586
rect 27304 -4636 27358 -4620
rect 27400 -4592 27466 -4582
rect 27400 -4626 27416 -4592
rect 27450 -4626 27466 -4592
rect 27400 -4636 27466 -4626
rect 27327 -4670 27357 -4636
rect 27423 -4670 27453 -4636
rect 27589 -4658 27619 -4500
rect 27672 -4570 27702 -4376
rect 27869 -4475 27899 -4460
rect 27793 -4505 27899 -4475
rect 27793 -4522 27823 -4505
rect 27757 -4538 27823 -4522
rect 27661 -4586 27715 -4570
rect 27661 -4620 27671 -4586
rect 27705 -4620 27715 -4586
rect 27757 -4572 27767 -4538
rect 27801 -4572 27823 -4538
rect 27968 -4510 27998 -4376
rect 28054 -4408 28084 -4376
rect 28040 -4424 28094 -4408
rect 28040 -4458 28050 -4424
rect 28084 -4458 28094 -4424
rect 28040 -4474 28094 -4458
rect 27968 -4522 28018 -4510
rect 27968 -4534 28031 -4522
rect 27968 -4540 28055 -4534
rect 27989 -4550 28055 -4540
rect 27989 -4552 28011 -4550
rect 27757 -4588 27823 -4572
rect 27793 -4614 27823 -4588
rect 27892 -4598 27959 -4582
rect 27661 -4636 27715 -4620
rect 27661 -4658 27691 -4636
rect 27892 -4632 27915 -4598
rect 27949 -4632 27959 -4598
rect 27892 -4648 27959 -4632
rect 28001 -4584 28011 -4552
rect 28045 -4584 28055 -4550
rect 28001 -4600 28055 -4584
rect 28138 -4560 28168 -4376
rect 28246 -4532 28276 -4376
rect 28330 -4424 28360 -4376
rect 28318 -4440 28372 -4424
rect 28318 -4474 28328 -4440
rect 28362 -4474 28372 -4440
rect 28318 -4490 28372 -4474
rect 28241 -4548 28295 -4532
rect 28138 -4576 28199 -4560
rect 28138 -4596 28155 -4576
rect 27892 -4670 27922 -4648
rect 28001 -4670 28031 -4600
rect 28097 -4610 28155 -4596
rect 28189 -4610 28199 -4576
rect 28241 -4582 28251 -4548
rect 28285 -4582 28295 -4548
rect 28241 -4598 28295 -4582
rect 28097 -4626 28199 -4610
rect 28097 -4658 28127 -4626
rect 28246 -4658 28276 -4598
rect 28337 -4658 28367 -4490
rect 28713 -4456 28743 -4420
rect 28702 -4486 28743 -4456
rect 28494 -4524 28524 -4492
rect 28702 -4524 28732 -4486
rect 29009 -4298 29039 -4272
rect 29093 -4298 29123 -4272
rect 29360 -4292 29390 -4266
rect 29452 -4292 29482 -4266
rect 29551 -4292 29581 -4266
rect 29691 -4292 29721 -4266
rect 29788 -4292 29818 -4266
rect 29985 -4292 30015 -4266
rect 30084 -4292 30114 -4266
rect 30170 -4292 30200 -4266
rect 30254 -4292 30284 -4266
rect 30362 -4292 30392 -4266
rect 30446 -4292 30476 -4266
rect 30610 -4292 30640 -4266
rect 30829 -4292 30859 -4266
rect 30926 -4292 30956 -4266
rect 29009 -4441 29039 -4426
rect 28976 -4471 29039 -4441
rect 28810 -4524 28840 -4492
rect 28976 -4524 29006 -4471
rect 29093 -4515 29123 -4426
rect 29360 -4463 29390 -4376
rect 29452 -4414 29482 -4376
rect 28423 -4540 28732 -4524
rect 28423 -4574 28451 -4540
rect 28485 -4574 28732 -4540
rect 28423 -4590 28732 -4574
rect 28781 -4540 28840 -4524
rect 28781 -4574 28791 -4540
rect 28825 -4574 28840 -4540
rect 28781 -4590 28840 -4574
rect 28952 -4540 29006 -4524
rect 28952 -4574 28962 -4540
rect 28996 -4574 29006 -4540
rect 29048 -4525 29123 -4515
rect 29048 -4559 29064 -4525
rect 29098 -4559 29123 -4525
rect 29261 -4479 29390 -4463
rect 29436 -4424 29502 -4414
rect 29436 -4458 29452 -4424
rect 29486 -4458 29502 -4424
rect 29436 -4468 29502 -4458
rect 29261 -4513 29271 -4479
rect 29305 -4493 29390 -4479
rect 29305 -4513 29378 -4493
rect 29551 -4510 29581 -4376
rect 29691 -4434 29721 -4376
rect 29691 -4450 29746 -4434
rect 29691 -4484 29701 -4450
rect 29735 -4484 29746 -4450
rect 29691 -4500 29746 -4484
rect 29261 -4529 29378 -4513
rect 29048 -4569 29123 -4559
rect 28952 -4590 29006 -4574
rect 28525 -4612 28555 -4590
rect 28702 -4613 28732 -4590
rect 28810 -4612 28840 -4590
rect 28702 -4643 28743 -4613
rect 28713 -4658 28743 -4643
rect 28976 -4613 29006 -4590
rect 28976 -4643 29039 -4613
rect 29009 -4658 29039 -4643
rect 29093 -4658 29123 -4569
rect 29348 -4658 29378 -4529
rect 29443 -4540 29581 -4510
rect 29443 -4570 29474 -4540
rect 29420 -4586 29474 -4570
rect 29420 -4620 29430 -4586
rect 29464 -4620 29474 -4586
rect 29420 -4636 29474 -4620
rect 29516 -4592 29582 -4582
rect 29516 -4626 29532 -4592
rect 29566 -4626 29582 -4592
rect 29516 -4636 29582 -4626
rect 29443 -4670 29473 -4636
rect 29539 -4670 29569 -4636
rect 29705 -4658 29735 -4500
rect 29788 -4570 29818 -4376
rect 29985 -4475 30015 -4460
rect 29909 -4505 30015 -4475
rect 29909 -4522 29939 -4505
rect 29873 -4538 29939 -4522
rect 29777 -4586 29831 -4570
rect 29777 -4620 29787 -4586
rect 29821 -4620 29831 -4586
rect 29873 -4572 29883 -4538
rect 29917 -4572 29939 -4538
rect 30084 -4510 30114 -4376
rect 30170 -4408 30200 -4376
rect 30156 -4424 30210 -4408
rect 30156 -4458 30166 -4424
rect 30200 -4458 30210 -4424
rect 30156 -4474 30210 -4458
rect 30084 -4522 30134 -4510
rect 30084 -4534 30147 -4522
rect 30084 -4540 30171 -4534
rect 30105 -4550 30171 -4540
rect 30105 -4552 30127 -4550
rect 29873 -4588 29939 -4572
rect 29909 -4614 29939 -4588
rect 30008 -4598 30075 -4582
rect 29777 -4636 29831 -4620
rect 29777 -4658 29807 -4636
rect 30008 -4632 30031 -4598
rect 30065 -4632 30075 -4598
rect 30008 -4648 30075 -4632
rect 30117 -4584 30127 -4552
rect 30161 -4584 30171 -4550
rect 30117 -4600 30171 -4584
rect 30254 -4560 30284 -4376
rect 30362 -4532 30392 -4376
rect 30446 -4424 30476 -4376
rect 30434 -4440 30488 -4424
rect 30434 -4474 30444 -4440
rect 30478 -4474 30488 -4440
rect 30434 -4490 30488 -4474
rect 30357 -4548 30411 -4532
rect 30254 -4576 30315 -4560
rect 30254 -4596 30271 -4576
rect 30008 -4670 30038 -4648
rect 30117 -4670 30147 -4600
rect 30213 -4610 30271 -4596
rect 30305 -4610 30315 -4576
rect 30357 -4582 30367 -4548
rect 30401 -4582 30411 -4548
rect 30357 -4598 30411 -4582
rect 30213 -4626 30315 -4610
rect 30213 -4658 30243 -4626
rect 30362 -4658 30392 -4598
rect 30453 -4658 30483 -4490
rect 30829 -4456 30859 -4420
rect 30818 -4486 30859 -4456
rect 30610 -4524 30640 -4492
rect 30818 -4524 30848 -4486
rect 31125 -4298 31155 -4272
rect 31209 -4298 31239 -4272
rect 31476 -4292 31506 -4266
rect 31568 -4292 31598 -4266
rect 31667 -4292 31697 -4266
rect 31807 -4292 31837 -4266
rect 31904 -4292 31934 -4266
rect 32101 -4292 32131 -4266
rect 32200 -4292 32230 -4266
rect 32286 -4292 32316 -4266
rect 32370 -4292 32400 -4266
rect 32478 -4292 32508 -4266
rect 32562 -4292 32592 -4266
rect 32726 -4292 32756 -4266
rect 32945 -4292 32975 -4266
rect 33042 -4292 33072 -4266
rect 31125 -4441 31155 -4426
rect 31092 -4471 31155 -4441
rect 30926 -4524 30956 -4492
rect 31092 -4524 31122 -4471
rect 31209 -4515 31239 -4426
rect 31476 -4463 31506 -4376
rect 31568 -4414 31598 -4376
rect 30539 -4540 30848 -4524
rect 30539 -4574 30567 -4540
rect 30601 -4574 30848 -4540
rect 30539 -4590 30848 -4574
rect 30897 -4540 30956 -4524
rect 30897 -4574 30907 -4540
rect 30941 -4574 30956 -4540
rect 30897 -4590 30956 -4574
rect 31068 -4540 31122 -4524
rect 31068 -4574 31078 -4540
rect 31112 -4574 31122 -4540
rect 31164 -4525 31239 -4515
rect 31164 -4559 31180 -4525
rect 31214 -4559 31239 -4525
rect 31377 -4479 31506 -4463
rect 31552 -4424 31618 -4414
rect 31552 -4458 31568 -4424
rect 31602 -4458 31618 -4424
rect 31552 -4468 31618 -4458
rect 31377 -4513 31387 -4479
rect 31421 -4493 31506 -4479
rect 31421 -4513 31494 -4493
rect 31667 -4510 31697 -4376
rect 31807 -4434 31837 -4376
rect 31807 -4450 31862 -4434
rect 31807 -4484 31817 -4450
rect 31851 -4484 31862 -4450
rect 31807 -4500 31862 -4484
rect 31377 -4529 31494 -4513
rect 31164 -4569 31239 -4559
rect 31068 -4590 31122 -4574
rect 30641 -4612 30671 -4590
rect 30818 -4613 30848 -4590
rect 30926 -4612 30956 -4590
rect 30818 -4643 30859 -4613
rect 30829 -4658 30859 -4643
rect 31092 -4613 31122 -4590
rect 31092 -4643 31155 -4613
rect 31125 -4658 31155 -4643
rect 31209 -4658 31239 -4569
rect 31464 -4658 31494 -4529
rect 31559 -4540 31697 -4510
rect 31559 -4570 31590 -4540
rect 31536 -4586 31590 -4570
rect 31536 -4620 31546 -4586
rect 31580 -4620 31590 -4586
rect 31536 -4636 31590 -4620
rect 31632 -4592 31698 -4582
rect 31632 -4626 31648 -4592
rect 31682 -4626 31698 -4592
rect 31632 -4636 31698 -4626
rect 31559 -4670 31589 -4636
rect 31655 -4670 31685 -4636
rect 31821 -4658 31851 -4500
rect 31904 -4570 31934 -4376
rect 32101 -4475 32131 -4460
rect 32025 -4505 32131 -4475
rect 32025 -4522 32055 -4505
rect 31989 -4538 32055 -4522
rect 31893 -4586 31947 -4570
rect 31893 -4620 31903 -4586
rect 31937 -4620 31947 -4586
rect 31989 -4572 31999 -4538
rect 32033 -4572 32055 -4538
rect 32200 -4510 32230 -4376
rect 32286 -4408 32316 -4376
rect 32272 -4424 32326 -4408
rect 32272 -4458 32282 -4424
rect 32316 -4458 32326 -4424
rect 32272 -4474 32326 -4458
rect 32200 -4522 32250 -4510
rect 32200 -4534 32263 -4522
rect 32200 -4540 32287 -4534
rect 32221 -4550 32287 -4540
rect 32221 -4552 32243 -4550
rect 31989 -4588 32055 -4572
rect 32025 -4614 32055 -4588
rect 32124 -4598 32191 -4582
rect 31893 -4636 31947 -4620
rect 31893 -4658 31923 -4636
rect 32124 -4632 32147 -4598
rect 32181 -4632 32191 -4598
rect 32124 -4648 32191 -4632
rect 32233 -4584 32243 -4552
rect 32277 -4584 32287 -4550
rect 32233 -4600 32287 -4584
rect 32370 -4560 32400 -4376
rect 32478 -4532 32508 -4376
rect 32562 -4424 32592 -4376
rect 32550 -4440 32604 -4424
rect 32550 -4474 32560 -4440
rect 32594 -4474 32604 -4440
rect 32550 -4490 32604 -4474
rect 32473 -4548 32527 -4532
rect 32370 -4576 32431 -4560
rect 32370 -4596 32387 -4576
rect 32124 -4670 32154 -4648
rect 32233 -4670 32263 -4600
rect 32329 -4610 32387 -4596
rect 32421 -4610 32431 -4576
rect 32473 -4582 32483 -4548
rect 32517 -4582 32527 -4548
rect 32473 -4598 32527 -4582
rect 32329 -4626 32431 -4610
rect 32329 -4658 32359 -4626
rect 32478 -4658 32508 -4598
rect 32569 -4658 32599 -4490
rect 32945 -4456 32975 -4420
rect 32934 -4486 32975 -4456
rect 32726 -4524 32756 -4492
rect 32934 -4524 32964 -4486
rect 33042 -4524 33072 -4492
rect 32655 -4540 32964 -4524
rect 32655 -4574 32683 -4540
rect 32717 -4574 32964 -4540
rect 32655 -4590 32964 -4574
rect 33013 -4540 33072 -4524
rect 33013 -4574 33023 -4540
rect 33057 -4574 33072 -4540
rect 33013 -4590 33072 -4574
rect 32757 -4612 32787 -4590
rect 32934 -4613 32964 -4590
rect 33042 -4612 33072 -4590
rect 32934 -4643 32975 -4613
rect 32945 -4658 32975 -4643
rect -9079 -4768 -9049 -4742
rect -8995 -4768 -8965 -4742
rect -8740 -4768 -8710 -4742
rect -8645 -4768 -8615 -4742
rect -8549 -4768 -8519 -4742
rect -8383 -4768 -8353 -4742
rect -8311 -4768 -8281 -4742
rect -8179 -4768 -8149 -4742
rect -8080 -4768 -8050 -4742
rect -7971 -4768 -7941 -4742
rect -7875 -4768 -7845 -4742
rect -7726 -4768 -7696 -4742
rect -7635 -4768 -7605 -4742
rect -7447 -4768 -7417 -4742
rect -7259 -4768 -7229 -4742
rect -7162 -4768 -7132 -4742
rect -6963 -4768 -6933 -4742
rect -6879 -4768 -6849 -4742
rect -6624 -4768 -6594 -4742
rect -6529 -4768 -6499 -4742
rect -6433 -4768 -6403 -4742
rect -6267 -4768 -6237 -4742
rect -6195 -4768 -6165 -4742
rect -6063 -4768 -6033 -4742
rect -5964 -4768 -5934 -4742
rect -5855 -4768 -5825 -4742
rect -5759 -4768 -5729 -4742
rect -5610 -4768 -5580 -4742
rect -5519 -4768 -5489 -4742
rect -5331 -4768 -5301 -4742
rect -5143 -4768 -5113 -4742
rect -5046 -4768 -5016 -4742
rect -4847 -4768 -4817 -4742
rect -4763 -4768 -4733 -4742
rect -4508 -4768 -4478 -4742
rect -4413 -4768 -4383 -4742
rect -4317 -4768 -4287 -4742
rect -4151 -4768 -4121 -4742
rect -4079 -4768 -4049 -4742
rect -3947 -4768 -3917 -4742
rect -3848 -4768 -3818 -4742
rect -3739 -4768 -3709 -4742
rect -3643 -4768 -3613 -4742
rect -3494 -4768 -3464 -4742
rect -3403 -4768 -3373 -4742
rect -3215 -4768 -3185 -4742
rect -3027 -4768 -2997 -4742
rect -2930 -4768 -2900 -4742
rect -2731 -4768 -2701 -4742
rect -2647 -4768 -2617 -4742
rect -2392 -4768 -2362 -4742
rect -2297 -4768 -2267 -4742
rect -2201 -4768 -2171 -4742
rect -2035 -4768 -2005 -4742
rect -1963 -4768 -1933 -4742
rect -1831 -4768 -1801 -4742
rect -1732 -4768 -1702 -4742
rect -1623 -4768 -1593 -4742
rect -1527 -4768 -1497 -4742
rect -1378 -4768 -1348 -4742
rect -1287 -4768 -1257 -4742
rect -1099 -4768 -1069 -4742
rect -911 -4768 -881 -4742
rect -814 -4768 -784 -4742
rect -615 -4768 -585 -4742
rect -531 -4768 -501 -4742
rect -276 -4768 -246 -4742
rect -181 -4768 -151 -4742
rect -85 -4768 -55 -4742
rect 81 -4768 111 -4742
rect 153 -4768 183 -4742
rect 285 -4768 315 -4742
rect 384 -4768 414 -4742
rect 493 -4768 523 -4742
rect 589 -4768 619 -4742
rect 738 -4768 768 -4742
rect 829 -4768 859 -4742
rect 1017 -4768 1047 -4742
rect 1205 -4768 1235 -4742
rect 1302 -4768 1332 -4742
rect 1501 -4768 1531 -4742
rect 1585 -4768 1615 -4742
rect 1840 -4768 1870 -4742
rect 1935 -4768 1965 -4742
rect 2031 -4768 2061 -4742
rect 2197 -4768 2227 -4742
rect 2269 -4768 2299 -4742
rect 2401 -4768 2431 -4742
rect 2500 -4768 2530 -4742
rect 2609 -4768 2639 -4742
rect 2705 -4768 2735 -4742
rect 2854 -4768 2884 -4742
rect 2945 -4768 2975 -4742
rect 3133 -4768 3163 -4742
rect 3321 -4768 3351 -4742
rect 3418 -4768 3448 -4742
rect 3617 -4768 3647 -4742
rect 3701 -4768 3731 -4742
rect 3956 -4768 3986 -4742
rect 4051 -4768 4081 -4742
rect 4147 -4768 4177 -4742
rect 4313 -4768 4343 -4742
rect 4385 -4768 4415 -4742
rect 4517 -4768 4547 -4742
rect 4616 -4768 4646 -4742
rect 4725 -4768 4755 -4742
rect 4821 -4768 4851 -4742
rect 4970 -4768 5000 -4742
rect 5061 -4768 5091 -4742
rect 5249 -4768 5279 -4742
rect 5437 -4768 5467 -4742
rect 5534 -4768 5564 -4742
rect 5733 -4768 5763 -4742
rect 5817 -4768 5847 -4742
rect 6072 -4768 6102 -4742
rect 6167 -4768 6197 -4742
rect 6263 -4768 6293 -4742
rect 6429 -4768 6459 -4742
rect 6501 -4768 6531 -4742
rect 6633 -4768 6663 -4742
rect 6732 -4768 6762 -4742
rect 6841 -4768 6871 -4742
rect 6937 -4768 6967 -4742
rect 7086 -4768 7116 -4742
rect 7177 -4768 7207 -4742
rect 7365 -4768 7395 -4742
rect 7553 -4768 7583 -4742
rect 7650 -4768 7680 -4742
rect 7849 -4768 7879 -4742
rect 7933 -4768 7963 -4742
rect 8188 -4768 8218 -4742
rect 8283 -4768 8313 -4742
rect 8379 -4768 8409 -4742
rect 8545 -4768 8575 -4742
rect 8617 -4768 8647 -4742
rect 8749 -4768 8779 -4742
rect 8848 -4768 8878 -4742
rect 8957 -4768 8987 -4742
rect 9053 -4768 9083 -4742
rect 9202 -4768 9232 -4742
rect 9293 -4768 9323 -4742
rect 9481 -4768 9511 -4742
rect 9669 -4768 9699 -4742
rect 9766 -4768 9796 -4742
rect 9965 -4768 9995 -4742
rect 10049 -4768 10079 -4742
rect 10304 -4768 10334 -4742
rect 10399 -4768 10429 -4742
rect 10495 -4768 10525 -4742
rect 10661 -4768 10691 -4742
rect 10733 -4768 10763 -4742
rect 10865 -4768 10895 -4742
rect 10964 -4768 10994 -4742
rect 11073 -4768 11103 -4742
rect 11169 -4768 11199 -4742
rect 11318 -4768 11348 -4742
rect 11409 -4768 11439 -4742
rect 11597 -4768 11627 -4742
rect 11785 -4768 11815 -4742
rect 11882 -4768 11912 -4742
rect 12081 -4768 12111 -4742
rect 12165 -4768 12195 -4742
rect 12420 -4768 12450 -4742
rect 12515 -4768 12545 -4742
rect 12611 -4768 12641 -4742
rect 12777 -4768 12807 -4742
rect 12849 -4768 12879 -4742
rect 12981 -4768 13011 -4742
rect 13080 -4768 13110 -4742
rect 13189 -4768 13219 -4742
rect 13285 -4768 13315 -4742
rect 13434 -4768 13464 -4742
rect 13525 -4768 13555 -4742
rect 13713 -4768 13743 -4742
rect 13901 -4768 13931 -4742
rect 13998 -4768 14028 -4742
rect 14197 -4768 14227 -4742
rect 14281 -4768 14311 -4742
rect 14536 -4768 14566 -4742
rect 14631 -4768 14661 -4742
rect 14727 -4768 14757 -4742
rect 14893 -4768 14923 -4742
rect 14965 -4768 14995 -4742
rect 15097 -4768 15127 -4742
rect 15196 -4768 15226 -4742
rect 15305 -4768 15335 -4742
rect 15401 -4768 15431 -4742
rect 15550 -4768 15580 -4742
rect 15641 -4768 15671 -4742
rect 15829 -4768 15859 -4742
rect 16017 -4768 16047 -4742
rect 16114 -4768 16144 -4742
rect 16313 -4768 16343 -4742
rect 16397 -4768 16427 -4742
rect 16652 -4768 16682 -4742
rect 16747 -4768 16777 -4742
rect 16843 -4768 16873 -4742
rect 17009 -4768 17039 -4742
rect 17081 -4768 17111 -4742
rect 17213 -4768 17243 -4742
rect 17312 -4768 17342 -4742
rect 17421 -4768 17451 -4742
rect 17517 -4768 17547 -4742
rect 17666 -4768 17696 -4742
rect 17757 -4768 17787 -4742
rect 17945 -4768 17975 -4742
rect 18133 -4768 18163 -4742
rect 18230 -4768 18260 -4742
rect 18429 -4768 18459 -4742
rect 18513 -4768 18543 -4742
rect 18768 -4768 18798 -4742
rect 18863 -4768 18893 -4742
rect 18959 -4768 18989 -4742
rect 19125 -4768 19155 -4742
rect 19197 -4768 19227 -4742
rect 19329 -4768 19359 -4742
rect 19428 -4768 19458 -4742
rect 19537 -4768 19567 -4742
rect 19633 -4768 19663 -4742
rect 19782 -4768 19812 -4742
rect 19873 -4768 19903 -4742
rect 20061 -4768 20091 -4742
rect 20249 -4768 20279 -4742
rect 20346 -4768 20376 -4742
rect 20545 -4768 20575 -4742
rect 20629 -4768 20659 -4742
rect 20884 -4768 20914 -4742
rect 20979 -4768 21009 -4742
rect 21075 -4768 21105 -4742
rect 21241 -4768 21271 -4742
rect 21313 -4768 21343 -4742
rect 21445 -4768 21475 -4742
rect 21544 -4768 21574 -4742
rect 21653 -4768 21683 -4742
rect 21749 -4768 21779 -4742
rect 21898 -4768 21928 -4742
rect 21989 -4768 22019 -4742
rect 22177 -4768 22207 -4742
rect 22365 -4768 22395 -4742
rect 22462 -4768 22492 -4742
rect 22661 -4768 22691 -4742
rect 22745 -4768 22775 -4742
rect 23000 -4768 23030 -4742
rect 23095 -4768 23125 -4742
rect 23191 -4768 23221 -4742
rect 23357 -4768 23387 -4742
rect 23429 -4768 23459 -4742
rect 23561 -4768 23591 -4742
rect 23660 -4768 23690 -4742
rect 23769 -4768 23799 -4742
rect 23865 -4768 23895 -4742
rect 24014 -4768 24044 -4742
rect 24105 -4768 24135 -4742
rect 24293 -4768 24323 -4742
rect 24481 -4768 24511 -4742
rect 24578 -4768 24608 -4742
rect 24777 -4768 24807 -4742
rect 24861 -4768 24891 -4742
rect 25116 -4768 25146 -4742
rect 25211 -4768 25241 -4742
rect 25307 -4768 25337 -4742
rect 25473 -4768 25503 -4742
rect 25545 -4768 25575 -4742
rect 25677 -4768 25707 -4742
rect 25776 -4768 25806 -4742
rect 25885 -4768 25915 -4742
rect 25981 -4768 26011 -4742
rect 26130 -4768 26160 -4742
rect 26221 -4768 26251 -4742
rect 26409 -4768 26439 -4742
rect 26597 -4768 26627 -4742
rect 26694 -4768 26724 -4742
rect 26893 -4768 26923 -4742
rect 26977 -4768 27007 -4742
rect 27232 -4768 27262 -4742
rect 27327 -4768 27357 -4742
rect 27423 -4768 27453 -4742
rect 27589 -4768 27619 -4742
rect 27661 -4768 27691 -4742
rect 27793 -4768 27823 -4742
rect 27892 -4768 27922 -4742
rect 28001 -4768 28031 -4742
rect 28097 -4768 28127 -4742
rect 28246 -4768 28276 -4742
rect 28337 -4768 28367 -4742
rect 28525 -4768 28555 -4742
rect 28713 -4768 28743 -4742
rect 28810 -4768 28840 -4742
rect 29009 -4768 29039 -4742
rect 29093 -4768 29123 -4742
rect 29348 -4768 29378 -4742
rect 29443 -4768 29473 -4742
rect 29539 -4768 29569 -4742
rect 29705 -4768 29735 -4742
rect 29777 -4768 29807 -4742
rect 29909 -4768 29939 -4742
rect 30008 -4768 30038 -4742
rect 30117 -4768 30147 -4742
rect 30213 -4768 30243 -4742
rect 30362 -4768 30392 -4742
rect 30453 -4768 30483 -4742
rect 30641 -4768 30671 -4742
rect 30829 -4768 30859 -4742
rect 30926 -4768 30956 -4742
rect 31125 -4768 31155 -4742
rect 31209 -4768 31239 -4742
rect 31464 -4768 31494 -4742
rect 31559 -4768 31589 -4742
rect 31655 -4768 31685 -4742
rect 31821 -4768 31851 -4742
rect 31893 -4768 31923 -4742
rect 32025 -4768 32055 -4742
rect 32124 -4768 32154 -4742
rect 32233 -4768 32263 -4742
rect 32329 -4768 32359 -4742
rect 32478 -4768 32508 -4742
rect 32569 -4768 32599 -4742
rect 32757 -4768 32787 -4742
rect 32945 -4768 32975 -4742
rect 33042 -4768 33072 -4742
rect 4415 -7551 6015 -7535
rect 4415 -7585 4431 -7551
rect 5796 -7585 6015 -7551
rect 4415 -7623 6015 -7585
rect 6073 -7551 7673 -7535
rect 6073 -7585 6290 -7551
rect 7657 -7585 7673 -7551
rect 6073 -7623 7673 -7585
rect 4415 -9061 6015 -9023
rect 4415 -9095 4431 -9061
rect 5796 -9095 6015 -9061
rect 4415 -9133 6015 -9095
rect 6073 -9061 7673 -9023
rect 6073 -9095 6290 -9061
rect 7657 -9095 7673 -9061
rect 6073 -9133 7673 -9095
rect 4415 -10571 6015 -10533
rect 4415 -10605 4431 -10571
rect 5796 -10605 6015 -10571
rect 4415 -10643 6015 -10605
rect 6073 -10571 7673 -10533
rect 6073 -10605 6290 -10571
rect 7657 -10605 7673 -10571
rect 6073 -10643 7673 -10605
rect 4415 -12081 6015 -12043
rect 4415 -12115 4431 -12081
rect 5796 -12115 6015 -12081
rect 4415 -12153 6015 -12115
rect 6073 -12081 7673 -12043
rect 6073 -12115 6290 -12081
rect 7657 -12115 7673 -12081
rect 6073 -12153 7673 -12115
rect 4415 -13591 6015 -13553
rect 4415 -13625 4431 -13591
rect 5796 -13625 6015 -13591
rect 4415 -13663 6015 -13625
rect 6073 -13591 7673 -13553
rect 6073 -13625 6290 -13591
rect 7657 -13625 7673 -13591
rect 6073 -13663 7673 -13625
rect 4415 -15101 6015 -15063
rect 4415 -15135 4431 -15101
rect 5796 -15135 6015 -15101
rect 4415 -15173 6015 -15135
rect 6073 -15101 7673 -15063
rect 6073 -15135 6290 -15101
rect 7657 -15135 7673 -15101
rect 6073 -15173 7673 -15135
rect 4415 -16611 6015 -16573
rect 4415 -16645 4431 -16611
rect 5796 -16645 6015 -16611
rect 4415 -16683 6015 -16645
rect 6073 -16611 7673 -16573
rect 6073 -16645 6290 -16611
rect 7657 -16645 7673 -16611
rect 6073 -16683 7673 -16645
rect 4415 -18121 6015 -18083
rect 4415 -18155 4431 -18121
rect 5796 -18155 6015 -18121
rect 4415 -18193 6015 -18155
rect 6073 -18121 7673 -18083
rect 6073 -18155 6290 -18121
rect 7657 -18155 7673 -18121
rect 6073 -18193 7673 -18155
rect 4415 -19631 6015 -19593
rect 4415 -19665 4431 -19631
rect 5796 -19665 6015 -19631
rect 4415 -19703 6015 -19665
rect 6073 -19631 7673 -19593
rect 6073 -19665 6290 -19631
rect 7657 -19665 7673 -19631
rect 6073 -19703 7673 -19665
rect 4415 -21141 6015 -21103
rect 4415 -21175 4431 -21141
rect 5796 -21175 6015 -21141
rect 4415 -21213 6015 -21175
rect 6073 -21141 7673 -21103
rect 6073 -21175 6290 -21141
rect 7657 -21175 7673 -21141
rect 6073 -21213 7673 -21175
rect 4415 -22651 6015 -22613
rect 4415 -22685 4431 -22651
rect 5796 -22685 6015 -22651
rect 4415 -22723 6015 -22685
rect 6073 -22651 7673 -22613
rect 6073 -22685 6290 -22651
rect 7657 -22685 7673 -22651
rect 6073 -22723 7673 -22685
rect 4415 -24161 6015 -24123
rect 4415 -24195 4431 -24161
rect 5796 -24195 6015 -24161
rect 4415 -24233 6015 -24195
rect 6073 -24161 7673 -24123
rect 6073 -24195 6290 -24161
rect 7657 -24195 7673 -24161
rect 6073 -24233 7673 -24195
rect 4415 -25671 6015 -25633
rect 4415 -25705 4431 -25671
rect 5796 -25705 6015 -25671
rect 4415 -25721 6015 -25705
rect 6073 -25671 7673 -25633
rect 6073 -25705 6290 -25671
rect 7657 -25705 7673 -25671
rect 6073 -25721 7673 -25705
rect 9500 -7594 9566 -7578
rect 9500 -7611 9516 -7594
rect 9433 -7628 9516 -7611
rect 9550 -7611 9566 -7594
rect 10160 -7594 10226 -7578
rect 10160 -7611 10176 -7594
rect 9550 -7628 9633 -7611
rect 9433 -7675 9633 -7628
rect 10093 -7628 10176 -7611
rect 10210 -7611 10226 -7594
rect 10630 -7594 10696 -7578
rect 10630 -7611 10646 -7594
rect 10210 -7628 10293 -7611
rect 10093 -7675 10293 -7628
rect 10563 -7628 10646 -7611
rect 10680 -7611 10696 -7594
rect 11233 -7595 11299 -7579
rect 10680 -7628 10763 -7611
rect 11233 -7612 11249 -7595
rect 10563 -7675 10763 -7628
rect 11166 -7629 11249 -7612
rect 11283 -7612 11299 -7595
rect 11491 -7595 11557 -7579
rect 11491 -7612 11507 -7595
rect 11283 -7629 11366 -7612
rect 11166 -7676 11366 -7629
rect 11424 -7629 11507 -7612
rect 11541 -7612 11557 -7595
rect 11749 -7595 11815 -7579
rect 11749 -7612 11765 -7595
rect 11541 -7629 11624 -7612
rect 11424 -7676 11624 -7629
rect 11682 -7629 11765 -7612
rect 11799 -7612 11815 -7595
rect 12007 -7595 12073 -7579
rect 12007 -7612 12023 -7595
rect 11799 -7629 11882 -7612
rect 11682 -7676 11882 -7629
rect 11940 -7629 12023 -7612
rect 12057 -7612 12073 -7595
rect 12265 -7595 12331 -7579
rect 12265 -7612 12281 -7595
rect 12057 -7629 12140 -7612
rect 11940 -7676 12140 -7629
rect 12198 -7629 12281 -7612
rect 12315 -7612 12331 -7595
rect 13048 -7595 13114 -7579
rect 13048 -7612 13064 -7595
rect 12315 -7629 12398 -7612
rect 12198 -7676 12398 -7629
rect 12981 -7629 13064 -7612
rect 13098 -7612 13114 -7595
rect 13306 -7595 13372 -7579
rect 13306 -7612 13322 -7595
rect 13098 -7629 13181 -7612
rect 12981 -7676 13181 -7629
rect 13239 -7629 13322 -7612
rect 13356 -7612 13372 -7595
rect 13564 -7595 13630 -7579
rect 13564 -7612 13580 -7595
rect 13356 -7629 13439 -7612
rect 13239 -7676 13439 -7629
rect 13497 -7629 13580 -7612
rect 13614 -7612 13630 -7595
rect 13822 -7595 13888 -7579
rect 13822 -7612 13838 -7595
rect 13614 -7629 13697 -7612
rect 13497 -7676 13697 -7629
rect 13755 -7629 13838 -7612
rect 13872 -7612 13888 -7595
rect 14080 -7595 14146 -7579
rect 14080 -7612 14096 -7595
rect 13872 -7629 13955 -7612
rect 13755 -7676 13955 -7629
rect 14013 -7629 14096 -7612
rect 14130 -7612 14146 -7595
rect 14854 -7595 14920 -7579
rect 14854 -7612 14870 -7595
rect 14130 -7629 14213 -7612
rect 14013 -7676 14213 -7629
rect 14787 -7629 14870 -7612
rect 14904 -7612 14920 -7595
rect 15112 -7595 15178 -7579
rect 15112 -7612 15128 -7595
rect 14904 -7629 14987 -7612
rect 14787 -7676 14987 -7629
rect 15045 -7629 15128 -7612
rect 15162 -7612 15178 -7595
rect 15370 -7595 15436 -7579
rect 15370 -7612 15386 -7595
rect 15162 -7629 15245 -7612
rect 15045 -7676 15245 -7629
rect 15303 -7629 15386 -7612
rect 15420 -7612 15436 -7595
rect 15628 -7595 15694 -7579
rect 15628 -7612 15644 -7595
rect 15420 -7629 15503 -7612
rect 15303 -7676 15503 -7629
rect 15561 -7629 15644 -7612
rect 15678 -7612 15694 -7595
rect 15886 -7595 15952 -7579
rect 15886 -7612 15902 -7595
rect 15678 -7629 15761 -7612
rect 15561 -7676 15761 -7629
rect 15819 -7629 15902 -7612
rect 15936 -7612 15952 -7595
rect 15936 -7629 16019 -7612
rect 15819 -7676 16019 -7629
rect 9433 -7922 9633 -7875
rect 9433 -7939 9516 -7922
rect 9500 -7956 9516 -7939
rect 9550 -7939 9633 -7922
rect 10093 -7922 10293 -7875
rect 10093 -7939 10176 -7922
rect 9550 -7956 9566 -7939
rect 9500 -7972 9566 -7956
rect 10160 -7956 10176 -7939
rect 10210 -7939 10293 -7922
rect 10563 -7922 10763 -7875
rect 10563 -7939 10646 -7922
rect 10210 -7956 10226 -7939
rect 10160 -7972 10226 -7956
rect 10630 -7956 10646 -7939
rect 10680 -7939 10763 -7922
rect 11166 -7923 11366 -7876
rect 10680 -7956 10696 -7939
rect 11166 -7940 11249 -7923
rect 10630 -7972 10696 -7956
rect 11233 -7957 11249 -7940
rect 11283 -7940 11366 -7923
rect 11424 -7923 11624 -7876
rect 11424 -7940 11507 -7923
rect 11283 -7957 11299 -7940
rect 11233 -7973 11299 -7957
rect 11491 -7957 11507 -7940
rect 11541 -7940 11624 -7923
rect 11682 -7923 11882 -7876
rect 11682 -7940 11765 -7923
rect 11541 -7957 11557 -7940
rect 11491 -7973 11557 -7957
rect 11749 -7957 11765 -7940
rect 11799 -7940 11882 -7923
rect 11940 -7923 12140 -7876
rect 11940 -7940 12023 -7923
rect 11799 -7957 11815 -7940
rect 11749 -7973 11815 -7957
rect 12007 -7957 12023 -7940
rect 12057 -7940 12140 -7923
rect 12198 -7923 12398 -7876
rect 12198 -7940 12281 -7923
rect 12057 -7957 12073 -7940
rect 12007 -7973 12073 -7957
rect 12265 -7957 12281 -7940
rect 12315 -7940 12398 -7923
rect 12981 -7923 13181 -7876
rect 12981 -7940 13064 -7923
rect 12315 -7957 12331 -7940
rect 12265 -7973 12331 -7957
rect 13048 -7957 13064 -7940
rect 13098 -7940 13181 -7923
rect 13239 -7923 13439 -7876
rect 13239 -7940 13322 -7923
rect 13098 -7957 13114 -7940
rect 13048 -7973 13114 -7957
rect 13306 -7957 13322 -7940
rect 13356 -7940 13439 -7923
rect 13497 -7923 13697 -7876
rect 13497 -7940 13580 -7923
rect 13356 -7957 13372 -7940
rect 13306 -7973 13372 -7957
rect 13564 -7957 13580 -7940
rect 13614 -7940 13697 -7923
rect 13755 -7923 13955 -7876
rect 13755 -7940 13838 -7923
rect 13614 -7957 13630 -7940
rect 13564 -7973 13630 -7957
rect 13822 -7957 13838 -7940
rect 13872 -7940 13955 -7923
rect 14013 -7923 14213 -7876
rect 14013 -7940 14096 -7923
rect 13872 -7957 13888 -7940
rect 13822 -7973 13888 -7957
rect 14080 -7957 14096 -7940
rect 14130 -7940 14213 -7923
rect 14787 -7923 14987 -7876
rect 14787 -7940 14870 -7923
rect 14130 -7957 14146 -7940
rect 14080 -7973 14146 -7957
rect 14854 -7957 14870 -7940
rect 14904 -7940 14987 -7923
rect 15045 -7923 15245 -7876
rect 15045 -7940 15128 -7923
rect 14904 -7957 14920 -7940
rect 14854 -7973 14920 -7957
rect 15112 -7957 15128 -7940
rect 15162 -7940 15245 -7923
rect 15303 -7923 15503 -7876
rect 15303 -7940 15386 -7923
rect 15162 -7957 15178 -7940
rect 15112 -7973 15178 -7957
rect 15370 -7957 15386 -7940
rect 15420 -7940 15503 -7923
rect 15561 -7923 15761 -7876
rect 15561 -7940 15644 -7923
rect 15420 -7957 15436 -7940
rect 15370 -7973 15436 -7957
rect 15628 -7957 15644 -7940
rect 15678 -7940 15761 -7923
rect 15819 -7923 16019 -7876
rect 15819 -7940 15902 -7923
rect 15678 -7957 15694 -7940
rect 15628 -7973 15694 -7957
rect 15886 -7957 15902 -7940
rect 15936 -7940 16019 -7923
rect 15936 -7957 15952 -7940
rect 15886 -7973 15952 -7957
rect 9384 -8561 9500 -8533
rect 9384 -8599 9408 -8561
rect 9474 -8599 9500 -8561
rect 10044 -8568 10230 -8552
rect 10044 -8585 10060 -8568
rect 9384 -8649 9500 -8599
rect 9737 -8602 10060 -8585
rect 10214 -8585 10230 -8568
rect 10770 -8561 10886 -8533
rect 10214 -8602 10537 -8585
rect 9737 -8649 10537 -8602
rect 10770 -8599 10794 -8561
rect 10860 -8599 10886 -8561
rect 10770 -8649 10886 -8599
rect 11140 -8561 11256 -8533
rect 11140 -8599 11164 -8561
rect 11230 -8599 11256 -8561
rect 11140 -8649 11256 -8599
rect 11562 -8561 11678 -8533
rect 11562 -8599 11586 -8561
rect 11652 -8599 11678 -8561
rect 11562 -8649 11678 -8599
rect 11984 -8561 12100 -8533
rect 11984 -8599 12008 -8561
rect 12074 -8599 12100 -8561
rect 12714 -8568 12900 -8552
rect 12714 -8585 12730 -8568
rect 11984 -8649 12100 -8599
rect 12407 -8602 12730 -8585
rect 12884 -8585 12900 -8568
rect 13484 -8561 13600 -8533
rect 12884 -8602 13207 -8585
rect 12407 -8649 13207 -8602
rect 13484 -8599 13508 -8561
rect 13574 -8599 13600 -8561
rect 13484 -8649 13600 -8599
rect 13854 -8561 13970 -8533
rect 13854 -8599 13878 -8561
rect 13944 -8599 13970 -8561
rect 13854 -8649 13970 -8599
rect 14276 -8561 14392 -8533
rect 14276 -8599 14300 -8561
rect 14366 -8599 14392 -8561
rect 14276 -8649 14392 -8599
rect 14698 -8561 14814 -8533
rect 14698 -8599 14722 -8561
rect 14788 -8599 14814 -8561
rect 15377 -8567 15563 -8551
rect 15377 -8584 15393 -8567
rect 14698 -8649 14814 -8599
rect 15070 -8601 15393 -8584
rect 15547 -8584 15563 -8567
rect 16138 -8561 16254 -8533
rect 15547 -8601 15870 -8584
rect 15070 -8648 15870 -8601
rect 16138 -8599 16162 -8561
rect 16228 -8599 16254 -8561
rect 16138 -8649 16254 -8599
rect 9384 -8823 9500 -8759
rect 9737 -8806 10537 -8759
rect 9737 -8823 10060 -8806
rect 10044 -8840 10060 -8823
rect 10214 -8823 10537 -8806
rect 10770 -8823 10886 -8759
rect 11140 -8823 11256 -8759
rect 11562 -8823 11678 -8759
rect 11984 -8823 12100 -8759
rect 12407 -8806 13207 -8759
rect 12407 -8823 12730 -8806
rect 10214 -8840 10230 -8823
rect 10044 -8856 10230 -8840
rect 12714 -8840 12730 -8823
rect 12884 -8823 13207 -8806
rect 13484 -8823 13600 -8759
rect 13854 -8823 13970 -8759
rect 14276 -8823 14392 -8759
rect 14698 -8823 14814 -8759
rect 15070 -8805 15870 -8758
rect 15070 -8822 15393 -8805
rect 12884 -8840 12900 -8823
rect 12714 -8856 12900 -8840
rect 15377 -8839 15393 -8822
rect 15547 -8822 15870 -8805
rect 15547 -8839 15563 -8822
rect 16138 -8823 16254 -8759
rect 15377 -8855 15563 -8839
rect 9226 -9564 9292 -9548
rect 9226 -9581 9242 -9564
rect 9159 -9598 9242 -9581
rect 9276 -9581 9292 -9564
rect 9484 -9564 9550 -9548
rect 9484 -9581 9500 -9564
rect 9276 -9598 9359 -9581
rect 9159 -9636 9359 -9598
rect 9417 -9598 9500 -9581
rect 9534 -9581 9550 -9564
rect 9742 -9564 9808 -9548
rect 9742 -9581 9758 -9564
rect 9534 -9598 9617 -9581
rect 9417 -9636 9617 -9598
rect 9675 -9598 9758 -9581
rect 9792 -9581 9808 -9564
rect 10000 -9564 10066 -9548
rect 10000 -9581 10016 -9564
rect 9792 -9598 9875 -9581
rect 9675 -9636 9875 -9598
rect 9933 -9598 10016 -9581
rect 10050 -9581 10066 -9564
rect 10258 -9564 10324 -9548
rect 10258 -9581 10274 -9564
rect 10050 -9598 10133 -9581
rect 9933 -9636 10133 -9598
rect 10191 -9598 10274 -9581
rect 10308 -9581 10324 -9564
rect 10516 -9564 10582 -9548
rect 10516 -9581 10532 -9564
rect 10308 -9598 10391 -9581
rect 10191 -9636 10391 -9598
rect 10449 -9598 10532 -9581
rect 10566 -9581 10582 -9564
rect 10774 -9564 10840 -9548
rect 10774 -9581 10790 -9564
rect 10566 -9598 10649 -9581
rect 10449 -9636 10649 -9598
rect 10707 -9598 10790 -9581
rect 10824 -9581 10840 -9564
rect 11032 -9564 11098 -9548
rect 11032 -9581 11048 -9564
rect 10824 -9598 10907 -9581
rect 10707 -9636 10907 -9598
rect 10965 -9598 11048 -9581
rect 11082 -9581 11098 -9564
rect 11896 -9564 11962 -9548
rect 11896 -9581 11912 -9564
rect 11082 -9598 11165 -9581
rect 10965 -9636 11165 -9598
rect 11829 -9598 11912 -9581
rect 11946 -9581 11962 -9564
rect 12154 -9564 12220 -9548
rect 12154 -9581 12170 -9564
rect 11946 -9598 12029 -9581
rect 11829 -9636 12029 -9598
rect 12087 -9598 12170 -9581
rect 12204 -9581 12220 -9564
rect 12412 -9564 12478 -9548
rect 12412 -9581 12428 -9564
rect 12204 -9598 12287 -9581
rect 12087 -9636 12287 -9598
rect 12345 -9598 12428 -9581
rect 12462 -9581 12478 -9564
rect 12670 -9564 12736 -9548
rect 12670 -9581 12686 -9564
rect 12462 -9598 12545 -9581
rect 12345 -9636 12545 -9598
rect 12603 -9598 12686 -9581
rect 12720 -9581 12736 -9564
rect 12928 -9564 12994 -9548
rect 12928 -9581 12944 -9564
rect 12720 -9598 12803 -9581
rect 12603 -9636 12803 -9598
rect 12861 -9598 12944 -9581
rect 12978 -9581 12994 -9564
rect 13186 -9564 13252 -9548
rect 13186 -9581 13202 -9564
rect 12978 -9598 13061 -9581
rect 12861 -9636 13061 -9598
rect 13119 -9598 13202 -9581
rect 13236 -9581 13252 -9564
rect 13444 -9564 13510 -9548
rect 13444 -9581 13460 -9564
rect 13236 -9598 13319 -9581
rect 13119 -9636 13319 -9598
rect 13377 -9598 13460 -9581
rect 13494 -9581 13510 -9564
rect 13702 -9564 13768 -9548
rect 13702 -9581 13718 -9564
rect 13494 -9598 13577 -9581
rect 13377 -9636 13577 -9598
rect 13635 -9598 13718 -9581
rect 13752 -9581 13768 -9564
rect 14559 -9563 14625 -9547
rect 14559 -9580 14575 -9563
rect 13752 -9598 13835 -9581
rect 13635 -9636 13835 -9598
rect 14492 -9597 14575 -9580
rect 14609 -9580 14625 -9563
rect 14817 -9563 14883 -9547
rect 14817 -9580 14833 -9563
rect 14609 -9597 14692 -9580
rect 14492 -9635 14692 -9597
rect 14750 -9597 14833 -9580
rect 14867 -9580 14883 -9563
rect 15075 -9563 15141 -9547
rect 15075 -9580 15091 -9563
rect 14867 -9597 14950 -9580
rect 14750 -9635 14950 -9597
rect 15008 -9597 15091 -9580
rect 15125 -9580 15141 -9563
rect 15333 -9563 15399 -9547
rect 15333 -9580 15349 -9563
rect 15125 -9597 15208 -9580
rect 15008 -9635 15208 -9597
rect 15266 -9597 15349 -9580
rect 15383 -9580 15399 -9563
rect 15591 -9563 15657 -9547
rect 15591 -9580 15607 -9563
rect 15383 -9597 15466 -9580
rect 15266 -9635 15466 -9597
rect 15524 -9597 15607 -9580
rect 15641 -9580 15657 -9563
rect 15849 -9563 15915 -9547
rect 15849 -9580 15865 -9563
rect 15641 -9597 15724 -9580
rect 15524 -9635 15724 -9597
rect 15782 -9597 15865 -9580
rect 15899 -9580 15915 -9563
rect 16107 -9563 16173 -9547
rect 16107 -9580 16123 -9563
rect 15899 -9597 15982 -9580
rect 15782 -9635 15982 -9597
rect 16040 -9597 16123 -9580
rect 16157 -9580 16173 -9563
rect 16365 -9563 16431 -9547
rect 16365 -9580 16381 -9563
rect 16157 -9597 16240 -9580
rect 16040 -9635 16240 -9597
rect 16298 -9597 16381 -9580
rect 16415 -9580 16431 -9563
rect 16415 -9597 16498 -9580
rect 16298 -9635 16498 -9597
rect 9159 -9874 9359 -9836
rect 9159 -9891 9242 -9874
rect 9226 -9908 9242 -9891
rect 9276 -9891 9359 -9874
rect 9417 -9874 9617 -9836
rect 9417 -9891 9500 -9874
rect 9276 -9908 9292 -9891
rect 9226 -9924 9292 -9908
rect 9484 -9908 9500 -9891
rect 9534 -9891 9617 -9874
rect 9675 -9874 9875 -9836
rect 9675 -9891 9758 -9874
rect 9534 -9908 9550 -9891
rect 9484 -9924 9550 -9908
rect 9742 -9908 9758 -9891
rect 9792 -9891 9875 -9874
rect 9933 -9874 10133 -9836
rect 9933 -9891 10016 -9874
rect 9792 -9908 9808 -9891
rect 9742 -9924 9808 -9908
rect 10000 -9908 10016 -9891
rect 10050 -9891 10133 -9874
rect 10191 -9874 10391 -9836
rect 10191 -9891 10274 -9874
rect 10050 -9908 10066 -9891
rect 10000 -9924 10066 -9908
rect 10258 -9908 10274 -9891
rect 10308 -9891 10391 -9874
rect 10449 -9874 10649 -9836
rect 10449 -9891 10532 -9874
rect 10308 -9908 10324 -9891
rect 10258 -9924 10324 -9908
rect 10516 -9908 10532 -9891
rect 10566 -9891 10649 -9874
rect 10707 -9874 10907 -9836
rect 10707 -9891 10790 -9874
rect 10566 -9908 10582 -9891
rect 10516 -9924 10582 -9908
rect 10774 -9908 10790 -9891
rect 10824 -9891 10907 -9874
rect 10965 -9874 11165 -9836
rect 10965 -9891 11048 -9874
rect 10824 -9908 10840 -9891
rect 10774 -9924 10840 -9908
rect 11032 -9908 11048 -9891
rect 11082 -9891 11165 -9874
rect 11829 -9874 12029 -9836
rect 11829 -9891 11912 -9874
rect 11082 -9908 11098 -9891
rect 11032 -9924 11098 -9908
rect 11896 -9908 11912 -9891
rect 11946 -9891 12029 -9874
rect 12087 -9874 12287 -9836
rect 12087 -9891 12170 -9874
rect 11946 -9908 11962 -9891
rect 11896 -9924 11962 -9908
rect 12154 -9908 12170 -9891
rect 12204 -9891 12287 -9874
rect 12345 -9874 12545 -9836
rect 12345 -9891 12428 -9874
rect 12204 -9908 12220 -9891
rect 12154 -9924 12220 -9908
rect 12412 -9908 12428 -9891
rect 12462 -9891 12545 -9874
rect 12603 -9874 12803 -9836
rect 12603 -9891 12686 -9874
rect 12462 -9908 12478 -9891
rect 12412 -9924 12478 -9908
rect 12670 -9908 12686 -9891
rect 12720 -9891 12803 -9874
rect 12861 -9874 13061 -9836
rect 12861 -9891 12944 -9874
rect 12720 -9908 12736 -9891
rect 12670 -9924 12736 -9908
rect 12928 -9908 12944 -9891
rect 12978 -9891 13061 -9874
rect 13119 -9874 13319 -9836
rect 13119 -9891 13202 -9874
rect 12978 -9908 12994 -9891
rect 12928 -9924 12994 -9908
rect 13186 -9908 13202 -9891
rect 13236 -9891 13319 -9874
rect 13377 -9874 13577 -9836
rect 13377 -9891 13460 -9874
rect 13236 -9908 13252 -9891
rect 13186 -9924 13252 -9908
rect 13444 -9908 13460 -9891
rect 13494 -9891 13577 -9874
rect 13635 -9874 13835 -9836
rect 13635 -9891 13718 -9874
rect 13494 -9908 13510 -9891
rect 13444 -9924 13510 -9908
rect 13702 -9908 13718 -9891
rect 13752 -9891 13835 -9874
rect 14492 -9873 14692 -9835
rect 14492 -9890 14575 -9873
rect 13752 -9908 13768 -9891
rect 13702 -9924 13768 -9908
rect 14559 -9907 14575 -9890
rect 14609 -9890 14692 -9873
rect 14750 -9873 14950 -9835
rect 14750 -9890 14833 -9873
rect 14609 -9907 14625 -9890
rect 14559 -9923 14625 -9907
rect 14817 -9907 14833 -9890
rect 14867 -9890 14950 -9873
rect 15008 -9873 15208 -9835
rect 15008 -9890 15091 -9873
rect 14867 -9907 14883 -9890
rect 14817 -9923 14883 -9907
rect 15075 -9907 15091 -9890
rect 15125 -9890 15208 -9873
rect 15266 -9873 15466 -9835
rect 15266 -9890 15349 -9873
rect 15125 -9907 15141 -9890
rect 15075 -9923 15141 -9907
rect 15333 -9907 15349 -9890
rect 15383 -9890 15466 -9873
rect 15524 -9873 15724 -9835
rect 15524 -9890 15607 -9873
rect 15383 -9907 15399 -9890
rect 15333 -9923 15399 -9907
rect 15591 -9907 15607 -9890
rect 15641 -9890 15724 -9873
rect 15782 -9873 15982 -9835
rect 15782 -9890 15865 -9873
rect 15641 -9907 15657 -9890
rect 15591 -9923 15657 -9907
rect 15849 -9907 15865 -9890
rect 15899 -9890 15982 -9873
rect 16040 -9873 16240 -9835
rect 16040 -9890 16123 -9873
rect 15899 -9907 15915 -9890
rect 15849 -9923 15915 -9907
rect 16107 -9907 16123 -9890
rect 16157 -9890 16240 -9873
rect 16298 -9873 16498 -9835
rect 16298 -9890 16381 -9873
rect 16157 -9907 16173 -9890
rect 16107 -9923 16173 -9907
rect 16365 -9907 16381 -9890
rect 16415 -9890 16498 -9873
rect 16415 -9907 16431 -9890
rect 16365 -9923 16431 -9907
rect 9226 -9982 9292 -9966
rect 9226 -9999 9242 -9982
rect 9159 -10016 9242 -9999
rect 9276 -9999 9292 -9982
rect 9484 -9982 9550 -9966
rect 9484 -9999 9500 -9982
rect 9276 -10016 9359 -9999
rect 9159 -10054 9359 -10016
rect 9417 -10016 9500 -9999
rect 9534 -9999 9550 -9982
rect 9742 -9982 9808 -9966
rect 9742 -9999 9758 -9982
rect 9534 -10016 9617 -9999
rect 9417 -10054 9617 -10016
rect 9675 -10016 9758 -9999
rect 9792 -9999 9808 -9982
rect 10000 -9982 10066 -9966
rect 10000 -9999 10016 -9982
rect 9792 -10016 9875 -9999
rect 9675 -10054 9875 -10016
rect 9933 -10016 10016 -9999
rect 10050 -9999 10066 -9982
rect 10258 -9982 10324 -9966
rect 10258 -9999 10274 -9982
rect 10050 -10016 10133 -9999
rect 9933 -10054 10133 -10016
rect 10191 -10016 10274 -9999
rect 10308 -9999 10324 -9982
rect 10516 -9982 10582 -9966
rect 10516 -9999 10532 -9982
rect 10308 -10016 10391 -9999
rect 10191 -10054 10391 -10016
rect 10449 -10016 10532 -9999
rect 10566 -9999 10582 -9982
rect 10774 -9982 10840 -9966
rect 10774 -9999 10790 -9982
rect 10566 -10016 10649 -9999
rect 10449 -10054 10649 -10016
rect 10707 -10016 10790 -9999
rect 10824 -9999 10840 -9982
rect 11032 -9982 11098 -9966
rect 11032 -9999 11048 -9982
rect 10824 -10016 10907 -9999
rect 10707 -10054 10907 -10016
rect 10965 -10016 11048 -9999
rect 11082 -9999 11098 -9982
rect 11896 -9982 11962 -9966
rect 11896 -9999 11912 -9982
rect 11082 -10016 11165 -9999
rect 10965 -10054 11165 -10016
rect 11829 -10016 11912 -9999
rect 11946 -9999 11962 -9982
rect 12154 -9982 12220 -9966
rect 12154 -9999 12170 -9982
rect 11946 -10016 12029 -9999
rect 11829 -10054 12029 -10016
rect 12087 -10016 12170 -9999
rect 12204 -9999 12220 -9982
rect 12412 -9982 12478 -9966
rect 12412 -9999 12428 -9982
rect 12204 -10016 12287 -9999
rect 12087 -10054 12287 -10016
rect 12345 -10016 12428 -9999
rect 12462 -9999 12478 -9982
rect 12670 -9982 12736 -9966
rect 12670 -9999 12686 -9982
rect 12462 -10016 12545 -9999
rect 12345 -10054 12545 -10016
rect 12603 -10016 12686 -9999
rect 12720 -9999 12736 -9982
rect 12928 -9982 12994 -9966
rect 12928 -9999 12944 -9982
rect 12720 -10016 12803 -9999
rect 12603 -10054 12803 -10016
rect 12861 -10016 12944 -9999
rect 12978 -9999 12994 -9982
rect 13186 -9982 13252 -9966
rect 13186 -9999 13202 -9982
rect 12978 -10016 13061 -9999
rect 12861 -10054 13061 -10016
rect 13119 -10016 13202 -9999
rect 13236 -9999 13252 -9982
rect 13444 -9982 13510 -9966
rect 13444 -9999 13460 -9982
rect 13236 -10016 13319 -9999
rect 13119 -10054 13319 -10016
rect 13377 -10016 13460 -9999
rect 13494 -9999 13510 -9982
rect 13702 -9982 13768 -9966
rect 13702 -9999 13718 -9982
rect 13494 -10016 13577 -9999
rect 13377 -10054 13577 -10016
rect 13635 -10016 13718 -9999
rect 13752 -9999 13768 -9982
rect 14559 -9981 14625 -9965
rect 14559 -9998 14575 -9981
rect 13752 -10016 13835 -9999
rect 13635 -10054 13835 -10016
rect 14492 -10015 14575 -9998
rect 14609 -9998 14625 -9981
rect 14817 -9981 14883 -9965
rect 14817 -9998 14833 -9981
rect 14609 -10015 14692 -9998
rect 14492 -10053 14692 -10015
rect 14750 -10015 14833 -9998
rect 14867 -9998 14883 -9981
rect 15075 -9981 15141 -9965
rect 15075 -9998 15091 -9981
rect 14867 -10015 14950 -9998
rect 14750 -10053 14950 -10015
rect 15008 -10015 15091 -9998
rect 15125 -9998 15141 -9981
rect 15333 -9981 15399 -9965
rect 15333 -9998 15349 -9981
rect 15125 -10015 15208 -9998
rect 15008 -10053 15208 -10015
rect 15266 -10015 15349 -9998
rect 15383 -9998 15399 -9981
rect 15591 -9981 15657 -9965
rect 15591 -9998 15607 -9981
rect 15383 -10015 15466 -9998
rect 15266 -10053 15466 -10015
rect 15524 -10015 15607 -9998
rect 15641 -9998 15657 -9981
rect 15849 -9981 15915 -9965
rect 15849 -9998 15865 -9981
rect 15641 -10015 15724 -9998
rect 15524 -10053 15724 -10015
rect 15782 -10015 15865 -9998
rect 15899 -9998 15915 -9981
rect 16107 -9981 16173 -9965
rect 16107 -9998 16123 -9981
rect 15899 -10015 15982 -9998
rect 15782 -10053 15982 -10015
rect 16040 -10015 16123 -9998
rect 16157 -9998 16173 -9981
rect 16365 -9981 16431 -9965
rect 16365 -9998 16381 -9981
rect 16157 -10015 16240 -9998
rect 16040 -10053 16240 -10015
rect 16298 -10015 16381 -9998
rect 16415 -9998 16431 -9981
rect 16415 -10015 16498 -9998
rect 16298 -10053 16498 -10015
rect 9159 -10292 9359 -10254
rect 9159 -10309 9242 -10292
rect 9226 -10326 9242 -10309
rect 9276 -10309 9359 -10292
rect 9417 -10292 9617 -10254
rect 9417 -10309 9500 -10292
rect 9276 -10326 9292 -10309
rect 9226 -10342 9292 -10326
rect 9484 -10326 9500 -10309
rect 9534 -10309 9617 -10292
rect 9675 -10292 9875 -10254
rect 9675 -10309 9758 -10292
rect 9534 -10326 9550 -10309
rect 9484 -10342 9550 -10326
rect 9742 -10326 9758 -10309
rect 9792 -10309 9875 -10292
rect 9933 -10292 10133 -10254
rect 9933 -10309 10016 -10292
rect 9792 -10326 9808 -10309
rect 9742 -10342 9808 -10326
rect 10000 -10326 10016 -10309
rect 10050 -10309 10133 -10292
rect 10191 -10292 10391 -10254
rect 10191 -10309 10274 -10292
rect 10050 -10326 10066 -10309
rect 10000 -10342 10066 -10326
rect 10258 -10326 10274 -10309
rect 10308 -10309 10391 -10292
rect 10449 -10292 10649 -10254
rect 10449 -10309 10532 -10292
rect 10308 -10326 10324 -10309
rect 10258 -10342 10324 -10326
rect 10516 -10326 10532 -10309
rect 10566 -10309 10649 -10292
rect 10707 -10292 10907 -10254
rect 10707 -10309 10790 -10292
rect 10566 -10326 10582 -10309
rect 10516 -10342 10582 -10326
rect 10774 -10326 10790 -10309
rect 10824 -10309 10907 -10292
rect 10965 -10292 11165 -10254
rect 10965 -10309 11048 -10292
rect 10824 -10326 10840 -10309
rect 10774 -10342 10840 -10326
rect 11032 -10326 11048 -10309
rect 11082 -10309 11165 -10292
rect 11829 -10292 12029 -10254
rect 11829 -10309 11912 -10292
rect 11082 -10326 11098 -10309
rect 11032 -10342 11098 -10326
rect 11896 -10326 11912 -10309
rect 11946 -10309 12029 -10292
rect 12087 -10292 12287 -10254
rect 12087 -10309 12170 -10292
rect 11946 -10326 11962 -10309
rect 11896 -10342 11962 -10326
rect 12154 -10326 12170 -10309
rect 12204 -10309 12287 -10292
rect 12345 -10292 12545 -10254
rect 12345 -10309 12428 -10292
rect 12204 -10326 12220 -10309
rect 12154 -10342 12220 -10326
rect 12412 -10326 12428 -10309
rect 12462 -10309 12545 -10292
rect 12603 -10292 12803 -10254
rect 12603 -10309 12686 -10292
rect 12462 -10326 12478 -10309
rect 12412 -10342 12478 -10326
rect 12670 -10326 12686 -10309
rect 12720 -10309 12803 -10292
rect 12861 -10292 13061 -10254
rect 12861 -10309 12944 -10292
rect 12720 -10326 12736 -10309
rect 12670 -10342 12736 -10326
rect 12928 -10326 12944 -10309
rect 12978 -10309 13061 -10292
rect 13119 -10292 13319 -10254
rect 13119 -10309 13202 -10292
rect 12978 -10326 12994 -10309
rect 12928 -10342 12994 -10326
rect 13186 -10326 13202 -10309
rect 13236 -10309 13319 -10292
rect 13377 -10292 13577 -10254
rect 13377 -10309 13460 -10292
rect 13236 -10326 13252 -10309
rect 13186 -10342 13252 -10326
rect 13444 -10326 13460 -10309
rect 13494 -10309 13577 -10292
rect 13635 -10292 13835 -10254
rect 13635 -10309 13718 -10292
rect 13494 -10326 13510 -10309
rect 13444 -10342 13510 -10326
rect 13702 -10326 13718 -10309
rect 13752 -10309 13835 -10292
rect 14492 -10291 14692 -10253
rect 14492 -10308 14575 -10291
rect 13752 -10326 13768 -10309
rect 13702 -10342 13768 -10326
rect 14559 -10325 14575 -10308
rect 14609 -10308 14692 -10291
rect 14750 -10291 14950 -10253
rect 14750 -10308 14833 -10291
rect 14609 -10325 14625 -10308
rect 14559 -10341 14625 -10325
rect 14817 -10325 14833 -10308
rect 14867 -10308 14950 -10291
rect 15008 -10291 15208 -10253
rect 15008 -10308 15091 -10291
rect 14867 -10325 14883 -10308
rect 14817 -10341 14883 -10325
rect 15075 -10325 15091 -10308
rect 15125 -10308 15208 -10291
rect 15266 -10291 15466 -10253
rect 15266 -10308 15349 -10291
rect 15125 -10325 15141 -10308
rect 15075 -10341 15141 -10325
rect 15333 -10325 15349 -10308
rect 15383 -10308 15466 -10291
rect 15524 -10291 15724 -10253
rect 15524 -10308 15607 -10291
rect 15383 -10325 15399 -10308
rect 15333 -10341 15399 -10325
rect 15591 -10325 15607 -10308
rect 15641 -10308 15724 -10291
rect 15782 -10291 15982 -10253
rect 15782 -10308 15865 -10291
rect 15641 -10325 15657 -10308
rect 15591 -10341 15657 -10325
rect 15849 -10325 15865 -10308
rect 15899 -10308 15982 -10291
rect 16040 -10291 16240 -10253
rect 16040 -10308 16123 -10291
rect 15899 -10325 15915 -10308
rect 15849 -10341 15915 -10325
rect 16107 -10325 16123 -10308
rect 16157 -10308 16240 -10291
rect 16298 -10291 16498 -10253
rect 16298 -10308 16381 -10291
rect 16157 -10325 16173 -10308
rect 16107 -10341 16173 -10325
rect 16365 -10325 16381 -10308
rect 16415 -10308 16498 -10291
rect 16415 -10325 16431 -10308
rect 16365 -10341 16431 -10325
rect 9226 -10400 9292 -10384
rect 9226 -10417 9242 -10400
rect 9159 -10434 9242 -10417
rect 9276 -10417 9292 -10400
rect 9484 -10400 9550 -10384
rect 9484 -10417 9500 -10400
rect 9276 -10434 9359 -10417
rect 9159 -10472 9359 -10434
rect 9417 -10434 9500 -10417
rect 9534 -10417 9550 -10400
rect 9742 -10400 9808 -10384
rect 9742 -10417 9758 -10400
rect 9534 -10434 9617 -10417
rect 9417 -10472 9617 -10434
rect 9675 -10434 9758 -10417
rect 9792 -10417 9808 -10400
rect 10000 -10400 10066 -10384
rect 10000 -10417 10016 -10400
rect 9792 -10434 9875 -10417
rect 9675 -10472 9875 -10434
rect 9933 -10434 10016 -10417
rect 10050 -10417 10066 -10400
rect 10258 -10400 10324 -10384
rect 10258 -10417 10274 -10400
rect 10050 -10434 10133 -10417
rect 9933 -10472 10133 -10434
rect 10191 -10434 10274 -10417
rect 10308 -10417 10324 -10400
rect 10516 -10400 10582 -10384
rect 10516 -10417 10532 -10400
rect 10308 -10434 10391 -10417
rect 10191 -10472 10391 -10434
rect 10449 -10434 10532 -10417
rect 10566 -10417 10582 -10400
rect 10774 -10400 10840 -10384
rect 10774 -10417 10790 -10400
rect 10566 -10434 10649 -10417
rect 10449 -10472 10649 -10434
rect 10707 -10434 10790 -10417
rect 10824 -10417 10840 -10400
rect 11032 -10400 11098 -10384
rect 11032 -10417 11048 -10400
rect 10824 -10434 10907 -10417
rect 10707 -10472 10907 -10434
rect 10965 -10434 11048 -10417
rect 11082 -10417 11098 -10400
rect 11896 -10400 11962 -10384
rect 11896 -10417 11912 -10400
rect 11082 -10434 11165 -10417
rect 10965 -10472 11165 -10434
rect 11829 -10434 11912 -10417
rect 11946 -10417 11962 -10400
rect 12154 -10400 12220 -10384
rect 12154 -10417 12170 -10400
rect 11946 -10434 12029 -10417
rect 11829 -10472 12029 -10434
rect 12087 -10434 12170 -10417
rect 12204 -10417 12220 -10400
rect 12412 -10400 12478 -10384
rect 12412 -10417 12428 -10400
rect 12204 -10434 12287 -10417
rect 12087 -10472 12287 -10434
rect 12345 -10434 12428 -10417
rect 12462 -10417 12478 -10400
rect 12670 -10400 12736 -10384
rect 12670 -10417 12686 -10400
rect 12462 -10434 12545 -10417
rect 12345 -10472 12545 -10434
rect 12603 -10434 12686 -10417
rect 12720 -10417 12736 -10400
rect 12928 -10400 12994 -10384
rect 12928 -10417 12944 -10400
rect 12720 -10434 12803 -10417
rect 12603 -10472 12803 -10434
rect 12861 -10434 12944 -10417
rect 12978 -10417 12994 -10400
rect 13186 -10400 13252 -10384
rect 13186 -10417 13202 -10400
rect 12978 -10434 13061 -10417
rect 12861 -10472 13061 -10434
rect 13119 -10434 13202 -10417
rect 13236 -10417 13252 -10400
rect 13444 -10400 13510 -10384
rect 13444 -10417 13460 -10400
rect 13236 -10434 13319 -10417
rect 13119 -10472 13319 -10434
rect 13377 -10434 13460 -10417
rect 13494 -10417 13510 -10400
rect 13702 -10400 13768 -10384
rect 13702 -10417 13718 -10400
rect 13494 -10434 13577 -10417
rect 13377 -10472 13577 -10434
rect 13635 -10434 13718 -10417
rect 13752 -10417 13768 -10400
rect 14559 -10399 14625 -10383
rect 14559 -10416 14575 -10399
rect 13752 -10434 13835 -10417
rect 13635 -10472 13835 -10434
rect 14492 -10433 14575 -10416
rect 14609 -10416 14625 -10399
rect 14817 -10399 14883 -10383
rect 14817 -10416 14833 -10399
rect 14609 -10433 14692 -10416
rect 14492 -10471 14692 -10433
rect 14750 -10433 14833 -10416
rect 14867 -10416 14883 -10399
rect 15075 -10399 15141 -10383
rect 15075 -10416 15091 -10399
rect 14867 -10433 14950 -10416
rect 14750 -10471 14950 -10433
rect 15008 -10433 15091 -10416
rect 15125 -10416 15141 -10399
rect 15333 -10399 15399 -10383
rect 15333 -10416 15349 -10399
rect 15125 -10433 15208 -10416
rect 15008 -10471 15208 -10433
rect 15266 -10433 15349 -10416
rect 15383 -10416 15399 -10399
rect 15591 -10399 15657 -10383
rect 15591 -10416 15607 -10399
rect 15383 -10433 15466 -10416
rect 15266 -10471 15466 -10433
rect 15524 -10433 15607 -10416
rect 15641 -10416 15657 -10399
rect 15849 -10399 15915 -10383
rect 15849 -10416 15865 -10399
rect 15641 -10433 15724 -10416
rect 15524 -10471 15724 -10433
rect 15782 -10433 15865 -10416
rect 15899 -10416 15915 -10399
rect 16107 -10399 16173 -10383
rect 16107 -10416 16123 -10399
rect 15899 -10433 15982 -10416
rect 15782 -10471 15982 -10433
rect 16040 -10433 16123 -10416
rect 16157 -10416 16173 -10399
rect 16365 -10399 16431 -10383
rect 16365 -10416 16381 -10399
rect 16157 -10433 16240 -10416
rect 16040 -10471 16240 -10433
rect 16298 -10433 16381 -10416
rect 16415 -10416 16431 -10399
rect 16415 -10433 16498 -10416
rect 16298 -10471 16498 -10433
rect 9159 -10710 9359 -10672
rect 9159 -10727 9242 -10710
rect 9226 -10744 9242 -10727
rect 9276 -10727 9359 -10710
rect 9417 -10710 9617 -10672
rect 9417 -10727 9500 -10710
rect 9276 -10744 9292 -10727
rect 9226 -10760 9292 -10744
rect 9484 -10744 9500 -10727
rect 9534 -10727 9617 -10710
rect 9675 -10710 9875 -10672
rect 9675 -10727 9758 -10710
rect 9534 -10744 9550 -10727
rect 9484 -10760 9550 -10744
rect 9742 -10744 9758 -10727
rect 9792 -10727 9875 -10710
rect 9933 -10710 10133 -10672
rect 9933 -10727 10016 -10710
rect 9792 -10744 9808 -10727
rect 9742 -10760 9808 -10744
rect 10000 -10744 10016 -10727
rect 10050 -10727 10133 -10710
rect 10191 -10710 10391 -10672
rect 10191 -10727 10274 -10710
rect 10050 -10744 10066 -10727
rect 10000 -10760 10066 -10744
rect 10258 -10744 10274 -10727
rect 10308 -10727 10391 -10710
rect 10449 -10710 10649 -10672
rect 10449 -10727 10532 -10710
rect 10308 -10744 10324 -10727
rect 10258 -10760 10324 -10744
rect 10516 -10744 10532 -10727
rect 10566 -10727 10649 -10710
rect 10707 -10710 10907 -10672
rect 10707 -10727 10790 -10710
rect 10566 -10744 10582 -10727
rect 10516 -10760 10582 -10744
rect 10774 -10744 10790 -10727
rect 10824 -10727 10907 -10710
rect 10965 -10710 11165 -10672
rect 10965 -10727 11048 -10710
rect 10824 -10744 10840 -10727
rect 10774 -10760 10840 -10744
rect 11032 -10744 11048 -10727
rect 11082 -10727 11165 -10710
rect 11829 -10710 12029 -10672
rect 11829 -10727 11912 -10710
rect 11082 -10744 11098 -10727
rect 11032 -10760 11098 -10744
rect 11896 -10744 11912 -10727
rect 11946 -10727 12029 -10710
rect 12087 -10710 12287 -10672
rect 12087 -10727 12170 -10710
rect 11946 -10744 11962 -10727
rect 11896 -10760 11962 -10744
rect 12154 -10744 12170 -10727
rect 12204 -10727 12287 -10710
rect 12345 -10710 12545 -10672
rect 12345 -10727 12428 -10710
rect 12204 -10744 12220 -10727
rect 12154 -10760 12220 -10744
rect 12412 -10744 12428 -10727
rect 12462 -10727 12545 -10710
rect 12603 -10710 12803 -10672
rect 12603 -10727 12686 -10710
rect 12462 -10744 12478 -10727
rect 12412 -10760 12478 -10744
rect 12670 -10744 12686 -10727
rect 12720 -10727 12803 -10710
rect 12861 -10710 13061 -10672
rect 12861 -10727 12944 -10710
rect 12720 -10744 12736 -10727
rect 12670 -10760 12736 -10744
rect 12928 -10744 12944 -10727
rect 12978 -10727 13061 -10710
rect 13119 -10710 13319 -10672
rect 13119 -10727 13202 -10710
rect 12978 -10744 12994 -10727
rect 12928 -10760 12994 -10744
rect 13186 -10744 13202 -10727
rect 13236 -10727 13319 -10710
rect 13377 -10710 13577 -10672
rect 13377 -10727 13460 -10710
rect 13236 -10744 13252 -10727
rect 13186 -10760 13252 -10744
rect 13444 -10744 13460 -10727
rect 13494 -10727 13577 -10710
rect 13635 -10710 13835 -10672
rect 13635 -10727 13718 -10710
rect 13494 -10744 13510 -10727
rect 13444 -10760 13510 -10744
rect 13702 -10744 13718 -10727
rect 13752 -10727 13835 -10710
rect 14492 -10709 14692 -10671
rect 14492 -10726 14575 -10709
rect 13752 -10744 13768 -10727
rect 13702 -10760 13768 -10744
rect 14559 -10743 14575 -10726
rect 14609 -10726 14692 -10709
rect 14750 -10709 14950 -10671
rect 14750 -10726 14833 -10709
rect 14609 -10743 14625 -10726
rect 14559 -10759 14625 -10743
rect 14817 -10743 14833 -10726
rect 14867 -10726 14950 -10709
rect 15008 -10709 15208 -10671
rect 15008 -10726 15091 -10709
rect 14867 -10743 14883 -10726
rect 14817 -10759 14883 -10743
rect 15075 -10743 15091 -10726
rect 15125 -10726 15208 -10709
rect 15266 -10709 15466 -10671
rect 15266 -10726 15349 -10709
rect 15125 -10743 15141 -10726
rect 15075 -10759 15141 -10743
rect 15333 -10743 15349 -10726
rect 15383 -10726 15466 -10709
rect 15524 -10709 15724 -10671
rect 15524 -10726 15607 -10709
rect 15383 -10743 15399 -10726
rect 15333 -10759 15399 -10743
rect 15591 -10743 15607 -10726
rect 15641 -10726 15724 -10709
rect 15782 -10709 15982 -10671
rect 15782 -10726 15865 -10709
rect 15641 -10743 15657 -10726
rect 15591 -10759 15657 -10743
rect 15849 -10743 15865 -10726
rect 15899 -10726 15982 -10709
rect 16040 -10709 16240 -10671
rect 16040 -10726 16123 -10709
rect 15899 -10743 15915 -10726
rect 15849 -10759 15915 -10743
rect 16107 -10743 16123 -10726
rect 16157 -10726 16240 -10709
rect 16298 -10709 16498 -10671
rect 16298 -10726 16381 -10709
rect 16157 -10743 16173 -10726
rect 16107 -10759 16173 -10743
rect 16365 -10743 16381 -10726
rect 16415 -10726 16498 -10709
rect 16415 -10743 16431 -10726
rect 16365 -10759 16431 -10743
rect 9226 -10818 9292 -10802
rect 9226 -10835 9242 -10818
rect 9159 -10852 9242 -10835
rect 9276 -10835 9292 -10818
rect 9484 -10818 9550 -10802
rect 9484 -10835 9500 -10818
rect 9276 -10852 9359 -10835
rect 9159 -10890 9359 -10852
rect 9417 -10852 9500 -10835
rect 9534 -10835 9550 -10818
rect 9742 -10818 9808 -10802
rect 9742 -10835 9758 -10818
rect 9534 -10852 9617 -10835
rect 9417 -10890 9617 -10852
rect 9675 -10852 9758 -10835
rect 9792 -10835 9808 -10818
rect 10000 -10818 10066 -10802
rect 10000 -10835 10016 -10818
rect 9792 -10852 9875 -10835
rect 9675 -10890 9875 -10852
rect 9933 -10852 10016 -10835
rect 10050 -10835 10066 -10818
rect 10258 -10818 10324 -10802
rect 10258 -10835 10274 -10818
rect 10050 -10852 10133 -10835
rect 9933 -10890 10133 -10852
rect 10191 -10852 10274 -10835
rect 10308 -10835 10324 -10818
rect 10516 -10818 10582 -10802
rect 10516 -10835 10532 -10818
rect 10308 -10852 10391 -10835
rect 10191 -10890 10391 -10852
rect 10449 -10852 10532 -10835
rect 10566 -10835 10582 -10818
rect 10774 -10818 10840 -10802
rect 10774 -10835 10790 -10818
rect 10566 -10852 10649 -10835
rect 10449 -10890 10649 -10852
rect 10707 -10852 10790 -10835
rect 10824 -10835 10840 -10818
rect 11032 -10818 11098 -10802
rect 11032 -10835 11048 -10818
rect 10824 -10852 10907 -10835
rect 10707 -10890 10907 -10852
rect 10965 -10852 11048 -10835
rect 11082 -10835 11098 -10818
rect 11896 -10818 11962 -10802
rect 11896 -10835 11912 -10818
rect 11082 -10852 11165 -10835
rect 10965 -10890 11165 -10852
rect 11829 -10852 11912 -10835
rect 11946 -10835 11962 -10818
rect 12154 -10818 12220 -10802
rect 12154 -10835 12170 -10818
rect 11946 -10852 12029 -10835
rect 11829 -10890 12029 -10852
rect 12087 -10852 12170 -10835
rect 12204 -10835 12220 -10818
rect 12412 -10818 12478 -10802
rect 12412 -10835 12428 -10818
rect 12204 -10852 12287 -10835
rect 12087 -10890 12287 -10852
rect 12345 -10852 12428 -10835
rect 12462 -10835 12478 -10818
rect 12670 -10818 12736 -10802
rect 12670 -10835 12686 -10818
rect 12462 -10852 12545 -10835
rect 12345 -10890 12545 -10852
rect 12603 -10852 12686 -10835
rect 12720 -10835 12736 -10818
rect 12928 -10818 12994 -10802
rect 12928 -10835 12944 -10818
rect 12720 -10852 12803 -10835
rect 12603 -10890 12803 -10852
rect 12861 -10852 12944 -10835
rect 12978 -10835 12994 -10818
rect 13186 -10818 13252 -10802
rect 13186 -10835 13202 -10818
rect 12978 -10852 13061 -10835
rect 12861 -10890 13061 -10852
rect 13119 -10852 13202 -10835
rect 13236 -10835 13252 -10818
rect 13444 -10818 13510 -10802
rect 13444 -10835 13460 -10818
rect 13236 -10852 13319 -10835
rect 13119 -10890 13319 -10852
rect 13377 -10852 13460 -10835
rect 13494 -10835 13510 -10818
rect 13702 -10818 13768 -10802
rect 13702 -10835 13718 -10818
rect 13494 -10852 13577 -10835
rect 13377 -10890 13577 -10852
rect 13635 -10852 13718 -10835
rect 13752 -10835 13768 -10818
rect 14559 -10817 14625 -10801
rect 14559 -10834 14575 -10817
rect 13752 -10852 13835 -10835
rect 13635 -10890 13835 -10852
rect 14492 -10851 14575 -10834
rect 14609 -10834 14625 -10817
rect 14817 -10817 14883 -10801
rect 14817 -10834 14833 -10817
rect 14609 -10851 14692 -10834
rect 14492 -10889 14692 -10851
rect 14750 -10851 14833 -10834
rect 14867 -10834 14883 -10817
rect 15075 -10817 15141 -10801
rect 15075 -10834 15091 -10817
rect 14867 -10851 14950 -10834
rect 14750 -10889 14950 -10851
rect 15008 -10851 15091 -10834
rect 15125 -10834 15141 -10817
rect 15333 -10817 15399 -10801
rect 15333 -10834 15349 -10817
rect 15125 -10851 15208 -10834
rect 15008 -10889 15208 -10851
rect 15266 -10851 15349 -10834
rect 15383 -10834 15399 -10817
rect 15591 -10817 15657 -10801
rect 15591 -10834 15607 -10817
rect 15383 -10851 15466 -10834
rect 15266 -10889 15466 -10851
rect 15524 -10851 15607 -10834
rect 15641 -10834 15657 -10817
rect 15849 -10817 15915 -10801
rect 15849 -10834 15865 -10817
rect 15641 -10851 15724 -10834
rect 15524 -10889 15724 -10851
rect 15782 -10851 15865 -10834
rect 15899 -10834 15915 -10817
rect 16107 -10817 16173 -10801
rect 16107 -10834 16123 -10817
rect 15899 -10851 15982 -10834
rect 15782 -10889 15982 -10851
rect 16040 -10851 16123 -10834
rect 16157 -10834 16173 -10817
rect 16365 -10817 16431 -10801
rect 16365 -10834 16381 -10817
rect 16157 -10851 16240 -10834
rect 16040 -10889 16240 -10851
rect 16298 -10851 16381 -10834
rect 16415 -10834 16431 -10817
rect 16415 -10851 16498 -10834
rect 16298 -10889 16498 -10851
rect 9159 -11128 9359 -11090
rect 9159 -11145 9242 -11128
rect 9226 -11162 9242 -11145
rect 9276 -11145 9359 -11128
rect 9417 -11128 9617 -11090
rect 9417 -11145 9500 -11128
rect 9276 -11162 9292 -11145
rect 9226 -11178 9292 -11162
rect 9484 -11162 9500 -11145
rect 9534 -11145 9617 -11128
rect 9675 -11128 9875 -11090
rect 9675 -11145 9758 -11128
rect 9534 -11162 9550 -11145
rect 9484 -11178 9550 -11162
rect 9742 -11162 9758 -11145
rect 9792 -11145 9875 -11128
rect 9933 -11128 10133 -11090
rect 9933 -11145 10016 -11128
rect 9792 -11162 9808 -11145
rect 9742 -11178 9808 -11162
rect 10000 -11162 10016 -11145
rect 10050 -11145 10133 -11128
rect 10191 -11128 10391 -11090
rect 10191 -11145 10274 -11128
rect 10050 -11162 10066 -11145
rect 10000 -11178 10066 -11162
rect 10258 -11162 10274 -11145
rect 10308 -11145 10391 -11128
rect 10449 -11128 10649 -11090
rect 10449 -11145 10532 -11128
rect 10308 -11162 10324 -11145
rect 10258 -11178 10324 -11162
rect 10516 -11162 10532 -11145
rect 10566 -11145 10649 -11128
rect 10707 -11128 10907 -11090
rect 10707 -11145 10790 -11128
rect 10566 -11162 10582 -11145
rect 10516 -11178 10582 -11162
rect 10774 -11162 10790 -11145
rect 10824 -11145 10907 -11128
rect 10965 -11128 11165 -11090
rect 10965 -11145 11048 -11128
rect 10824 -11162 10840 -11145
rect 10774 -11178 10840 -11162
rect 11032 -11162 11048 -11145
rect 11082 -11145 11165 -11128
rect 11829 -11128 12029 -11090
rect 11829 -11145 11912 -11128
rect 11082 -11162 11098 -11145
rect 11032 -11178 11098 -11162
rect 11896 -11162 11912 -11145
rect 11946 -11145 12029 -11128
rect 12087 -11128 12287 -11090
rect 12087 -11145 12170 -11128
rect 11946 -11162 11962 -11145
rect 11896 -11178 11962 -11162
rect 12154 -11162 12170 -11145
rect 12204 -11145 12287 -11128
rect 12345 -11128 12545 -11090
rect 12345 -11145 12428 -11128
rect 12204 -11162 12220 -11145
rect 12154 -11178 12220 -11162
rect 12412 -11162 12428 -11145
rect 12462 -11145 12545 -11128
rect 12603 -11128 12803 -11090
rect 12603 -11145 12686 -11128
rect 12462 -11162 12478 -11145
rect 12412 -11178 12478 -11162
rect 12670 -11162 12686 -11145
rect 12720 -11145 12803 -11128
rect 12861 -11128 13061 -11090
rect 12861 -11145 12944 -11128
rect 12720 -11162 12736 -11145
rect 12670 -11178 12736 -11162
rect 12928 -11162 12944 -11145
rect 12978 -11145 13061 -11128
rect 13119 -11128 13319 -11090
rect 13119 -11145 13202 -11128
rect 12978 -11162 12994 -11145
rect 12928 -11178 12994 -11162
rect 13186 -11162 13202 -11145
rect 13236 -11145 13319 -11128
rect 13377 -11128 13577 -11090
rect 13377 -11145 13460 -11128
rect 13236 -11162 13252 -11145
rect 13186 -11178 13252 -11162
rect 13444 -11162 13460 -11145
rect 13494 -11145 13577 -11128
rect 13635 -11128 13835 -11090
rect 13635 -11145 13718 -11128
rect 13494 -11162 13510 -11145
rect 13444 -11178 13510 -11162
rect 13702 -11162 13718 -11145
rect 13752 -11145 13835 -11128
rect 14492 -11127 14692 -11089
rect 14492 -11144 14575 -11127
rect 13752 -11162 13768 -11145
rect 13702 -11178 13768 -11162
rect 14559 -11161 14575 -11144
rect 14609 -11144 14692 -11127
rect 14750 -11127 14950 -11089
rect 14750 -11144 14833 -11127
rect 14609 -11161 14625 -11144
rect 14559 -11177 14625 -11161
rect 14817 -11161 14833 -11144
rect 14867 -11144 14950 -11127
rect 15008 -11127 15208 -11089
rect 15008 -11144 15091 -11127
rect 14867 -11161 14883 -11144
rect 14817 -11177 14883 -11161
rect 15075 -11161 15091 -11144
rect 15125 -11144 15208 -11127
rect 15266 -11127 15466 -11089
rect 15266 -11144 15349 -11127
rect 15125 -11161 15141 -11144
rect 15075 -11177 15141 -11161
rect 15333 -11161 15349 -11144
rect 15383 -11144 15466 -11127
rect 15524 -11127 15724 -11089
rect 15524 -11144 15607 -11127
rect 15383 -11161 15399 -11144
rect 15333 -11177 15399 -11161
rect 15591 -11161 15607 -11144
rect 15641 -11144 15724 -11127
rect 15782 -11127 15982 -11089
rect 15782 -11144 15865 -11127
rect 15641 -11161 15657 -11144
rect 15591 -11177 15657 -11161
rect 15849 -11161 15865 -11144
rect 15899 -11144 15982 -11127
rect 16040 -11127 16240 -11089
rect 16040 -11144 16123 -11127
rect 15899 -11161 15915 -11144
rect 15849 -11177 15915 -11161
rect 16107 -11161 16123 -11144
rect 16157 -11144 16240 -11127
rect 16298 -11127 16498 -11089
rect 16298 -11144 16381 -11127
rect 16157 -11161 16173 -11144
rect 16107 -11177 16173 -11161
rect 16365 -11161 16381 -11144
rect 16415 -11144 16498 -11127
rect 16415 -11161 16431 -11144
rect 16365 -11177 16431 -11161
rect 9226 -11236 9292 -11220
rect 9226 -11253 9242 -11236
rect 9159 -11270 9242 -11253
rect 9276 -11253 9292 -11236
rect 9484 -11236 9550 -11220
rect 9484 -11253 9500 -11236
rect 9276 -11270 9359 -11253
rect 9159 -11308 9359 -11270
rect 9417 -11270 9500 -11253
rect 9534 -11253 9550 -11236
rect 9742 -11236 9808 -11220
rect 9742 -11253 9758 -11236
rect 9534 -11270 9617 -11253
rect 9417 -11308 9617 -11270
rect 9675 -11270 9758 -11253
rect 9792 -11253 9808 -11236
rect 10000 -11236 10066 -11220
rect 10000 -11253 10016 -11236
rect 9792 -11270 9875 -11253
rect 9675 -11308 9875 -11270
rect 9933 -11270 10016 -11253
rect 10050 -11253 10066 -11236
rect 10258 -11236 10324 -11220
rect 10258 -11253 10274 -11236
rect 10050 -11270 10133 -11253
rect 9933 -11308 10133 -11270
rect 10191 -11270 10274 -11253
rect 10308 -11253 10324 -11236
rect 10516 -11236 10582 -11220
rect 10516 -11253 10532 -11236
rect 10308 -11270 10391 -11253
rect 10191 -11308 10391 -11270
rect 10449 -11270 10532 -11253
rect 10566 -11253 10582 -11236
rect 10774 -11236 10840 -11220
rect 10774 -11253 10790 -11236
rect 10566 -11270 10649 -11253
rect 10449 -11308 10649 -11270
rect 10707 -11270 10790 -11253
rect 10824 -11253 10840 -11236
rect 11032 -11236 11098 -11220
rect 11032 -11253 11048 -11236
rect 10824 -11270 10907 -11253
rect 10707 -11308 10907 -11270
rect 10965 -11270 11048 -11253
rect 11082 -11253 11098 -11236
rect 11896 -11236 11962 -11220
rect 11896 -11253 11912 -11236
rect 11082 -11270 11165 -11253
rect 10965 -11308 11165 -11270
rect 11829 -11270 11912 -11253
rect 11946 -11253 11962 -11236
rect 12154 -11236 12220 -11220
rect 12154 -11253 12170 -11236
rect 11946 -11270 12029 -11253
rect 11829 -11308 12029 -11270
rect 12087 -11270 12170 -11253
rect 12204 -11253 12220 -11236
rect 12412 -11236 12478 -11220
rect 12412 -11253 12428 -11236
rect 12204 -11270 12287 -11253
rect 12087 -11308 12287 -11270
rect 12345 -11270 12428 -11253
rect 12462 -11253 12478 -11236
rect 12670 -11236 12736 -11220
rect 12670 -11253 12686 -11236
rect 12462 -11270 12545 -11253
rect 12345 -11308 12545 -11270
rect 12603 -11270 12686 -11253
rect 12720 -11253 12736 -11236
rect 12928 -11236 12994 -11220
rect 12928 -11253 12944 -11236
rect 12720 -11270 12803 -11253
rect 12603 -11308 12803 -11270
rect 12861 -11270 12944 -11253
rect 12978 -11253 12994 -11236
rect 13186 -11236 13252 -11220
rect 13186 -11253 13202 -11236
rect 12978 -11270 13061 -11253
rect 12861 -11308 13061 -11270
rect 13119 -11270 13202 -11253
rect 13236 -11253 13252 -11236
rect 13444 -11236 13510 -11220
rect 13444 -11253 13460 -11236
rect 13236 -11270 13319 -11253
rect 13119 -11308 13319 -11270
rect 13377 -11270 13460 -11253
rect 13494 -11253 13510 -11236
rect 13702 -11236 13768 -11220
rect 13702 -11253 13718 -11236
rect 13494 -11270 13577 -11253
rect 13377 -11308 13577 -11270
rect 13635 -11270 13718 -11253
rect 13752 -11253 13768 -11236
rect 14559 -11235 14625 -11219
rect 14559 -11252 14575 -11235
rect 13752 -11270 13835 -11253
rect 13635 -11308 13835 -11270
rect 14492 -11269 14575 -11252
rect 14609 -11252 14625 -11235
rect 14817 -11235 14883 -11219
rect 14817 -11252 14833 -11235
rect 14609 -11269 14692 -11252
rect 14492 -11307 14692 -11269
rect 14750 -11269 14833 -11252
rect 14867 -11252 14883 -11235
rect 15075 -11235 15141 -11219
rect 15075 -11252 15091 -11235
rect 14867 -11269 14950 -11252
rect 14750 -11307 14950 -11269
rect 15008 -11269 15091 -11252
rect 15125 -11252 15141 -11235
rect 15333 -11235 15399 -11219
rect 15333 -11252 15349 -11235
rect 15125 -11269 15208 -11252
rect 15008 -11307 15208 -11269
rect 15266 -11269 15349 -11252
rect 15383 -11252 15399 -11235
rect 15591 -11235 15657 -11219
rect 15591 -11252 15607 -11235
rect 15383 -11269 15466 -11252
rect 15266 -11307 15466 -11269
rect 15524 -11269 15607 -11252
rect 15641 -11252 15657 -11235
rect 15849 -11235 15915 -11219
rect 15849 -11252 15865 -11235
rect 15641 -11269 15724 -11252
rect 15524 -11307 15724 -11269
rect 15782 -11269 15865 -11252
rect 15899 -11252 15915 -11235
rect 16107 -11235 16173 -11219
rect 16107 -11252 16123 -11235
rect 15899 -11269 15982 -11252
rect 15782 -11307 15982 -11269
rect 16040 -11269 16123 -11252
rect 16157 -11252 16173 -11235
rect 16365 -11235 16431 -11219
rect 16365 -11252 16381 -11235
rect 16157 -11269 16240 -11252
rect 16040 -11307 16240 -11269
rect 16298 -11269 16381 -11252
rect 16415 -11252 16431 -11235
rect 16415 -11269 16498 -11252
rect 16298 -11307 16498 -11269
rect 9159 -11546 9359 -11508
rect 9159 -11563 9242 -11546
rect 9226 -11580 9242 -11563
rect 9276 -11563 9359 -11546
rect 9417 -11546 9617 -11508
rect 9417 -11563 9500 -11546
rect 9276 -11580 9292 -11563
rect 9226 -11596 9292 -11580
rect 9484 -11580 9500 -11563
rect 9534 -11563 9617 -11546
rect 9675 -11546 9875 -11508
rect 9675 -11563 9758 -11546
rect 9534 -11580 9550 -11563
rect 9484 -11596 9550 -11580
rect 9742 -11580 9758 -11563
rect 9792 -11563 9875 -11546
rect 9933 -11546 10133 -11508
rect 9933 -11563 10016 -11546
rect 9792 -11580 9808 -11563
rect 9742 -11596 9808 -11580
rect 10000 -11580 10016 -11563
rect 10050 -11563 10133 -11546
rect 10191 -11546 10391 -11508
rect 10191 -11563 10274 -11546
rect 10050 -11580 10066 -11563
rect 10000 -11596 10066 -11580
rect 10258 -11580 10274 -11563
rect 10308 -11563 10391 -11546
rect 10449 -11546 10649 -11508
rect 10449 -11563 10532 -11546
rect 10308 -11580 10324 -11563
rect 10258 -11596 10324 -11580
rect 10516 -11580 10532 -11563
rect 10566 -11563 10649 -11546
rect 10707 -11546 10907 -11508
rect 10707 -11563 10790 -11546
rect 10566 -11580 10582 -11563
rect 10516 -11596 10582 -11580
rect 10774 -11580 10790 -11563
rect 10824 -11563 10907 -11546
rect 10965 -11546 11165 -11508
rect 10965 -11563 11048 -11546
rect 10824 -11580 10840 -11563
rect 10774 -11596 10840 -11580
rect 11032 -11580 11048 -11563
rect 11082 -11563 11165 -11546
rect 11829 -11546 12029 -11508
rect 11829 -11563 11912 -11546
rect 11082 -11580 11098 -11563
rect 11032 -11596 11098 -11580
rect 11896 -11580 11912 -11563
rect 11946 -11563 12029 -11546
rect 12087 -11546 12287 -11508
rect 12087 -11563 12170 -11546
rect 11946 -11580 11962 -11563
rect 11896 -11596 11962 -11580
rect 12154 -11580 12170 -11563
rect 12204 -11563 12287 -11546
rect 12345 -11546 12545 -11508
rect 12345 -11563 12428 -11546
rect 12204 -11580 12220 -11563
rect 12154 -11596 12220 -11580
rect 12412 -11580 12428 -11563
rect 12462 -11563 12545 -11546
rect 12603 -11546 12803 -11508
rect 12603 -11563 12686 -11546
rect 12462 -11580 12478 -11563
rect 12412 -11596 12478 -11580
rect 12670 -11580 12686 -11563
rect 12720 -11563 12803 -11546
rect 12861 -11546 13061 -11508
rect 12861 -11563 12944 -11546
rect 12720 -11580 12736 -11563
rect 12670 -11596 12736 -11580
rect 12928 -11580 12944 -11563
rect 12978 -11563 13061 -11546
rect 13119 -11546 13319 -11508
rect 13119 -11563 13202 -11546
rect 12978 -11580 12994 -11563
rect 12928 -11596 12994 -11580
rect 13186 -11580 13202 -11563
rect 13236 -11563 13319 -11546
rect 13377 -11546 13577 -11508
rect 13377 -11563 13460 -11546
rect 13236 -11580 13252 -11563
rect 13186 -11596 13252 -11580
rect 13444 -11580 13460 -11563
rect 13494 -11563 13577 -11546
rect 13635 -11546 13835 -11508
rect 13635 -11563 13718 -11546
rect 13494 -11580 13510 -11563
rect 13444 -11596 13510 -11580
rect 13702 -11580 13718 -11563
rect 13752 -11563 13835 -11546
rect 14492 -11545 14692 -11507
rect 14492 -11562 14575 -11545
rect 13752 -11580 13768 -11563
rect 13702 -11596 13768 -11580
rect 14559 -11579 14575 -11562
rect 14609 -11562 14692 -11545
rect 14750 -11545 14950 -11507
rect 14750 -11562 14833 -11545
rect 14609 -11579 14625 -11562
rect 14559 -11595 14625 -11579
rect 14817 -11579 14833 -11562
rect 14867 -11562 14950 -11545
rect 15008 -11545 15208 -11507
rect 15008 -11562 15091 -11545
rect 14867 -11579 14883 -11562
rect 14817 -11595 14883 -11579
rect 15075 -11579 15091 -11562
rect 15125 -11562 15208 -11545
rect 15266 -11545 15466 -11507
rect 15266 -11562 15349 -11545
rect 15125 -11579 15141 -11562
rect 15075 -11595 15141 -11579
rect 15333 -11579 15349 -11562
rect 15383 -11562 15466 -11545
rect 15524 -11545 15724 -11507
rect 15524 -11562 15607 -11545
rect 15383 -11579 15399 -11562
rect 15333 -11595 15399 -11579
rect 15591 -11579 15607 -11562
rect 15641 -11562 15724 -11545
rect 15782 -11545 15982 -11507
rect 15782 -11562 15865 -11545
rect 15641 -11579 15657 -11562
rect 15591 -11595 15657 -11579
rect 15849 -11579 15865 -11562
rect 15899 -11562 15982 -11545
rect 16040 -11545 16240 -11507
rect 16040 -11562 16123 -11545
rect 15899 -11579 15915 -11562
rect 15849 -11595 15915 -11579
rect 16107 -11579 16123 -11562
rect 16157 -11562 16240 -11545
rect 16298 -11545 16498 -11507
rect 16298 -11562 16381 -11545
rect 16157 -11579 16173 -11562
rect 16107 -11595 16173 -11579
rect 16365 -11579 16381 -11562
rect 16415 -11562 16498 -11545
rect 16415 -11579 16431 -11562
rect 16365 -11595 16431 -11579
rect 9226 -11654 9292 -11638
rect 9226 -11671 9242 -11654
rect 9159 -11688 9242 -11671
rect 9276 -11671 9292 -11654
rect 9484 -11654 9550 -11638
rect 9484 -11671 9500 -11654
rect 9276 -11688 9359 -11671
rect 9159 -11726 9359 -11688
rect 9417 -11688 9500 -11671
rect 9534 -11671 9550 -11654
rect 9742 -11654 9808 -11638
rect 9742 -11671 9758 -11654
rect 9534 -11688 9617 -11671
rect 9417 -11726 9617 -11688
rect 9675 -11688 9758 -11671
rect 9792 -11671 9808 -11654
rect 10000 -11654 10066 -11638
rect 10000 -11671 10016 -11654
rect 9792 -11688 9875 -11671
rect 9675 -11726 9875 -11688
rect 9933 -11688 10016 -11671
rect 10050 -11671 10066 -11654
rect 10258 -11654 10324 -11638
rect 10258 -11671 10274 -11654
rect 10050 -11688 10133 -11671
rect 9933 -11726 10133 -11688
rect 10191 -11688 10274 -11671
rect 10308 -11671 10324 -11654
rect 10516 -11654 10582 -11638
rect 10516 -11671 10532 -11654
rect 10308 -11688 10391 -11671
rect 10191 -11726 10391 -11688
rect 10449 -11688 10532 -11671
rect 10566 -11671 10582 -11654
rect 10774 -11654 10840 -11638
rect 10774 -11671 10790 -11654
rect 10566 -11688 10649 -11671
rect 10449 -11726 10649 -11688
rect 10707 -11688 10790 -11671
rect 10824 -11671 10840 -11654
rect 11032 -11654 11098 -11638
rect 11032 -11671 11048 -11654
rect 10824 -11688 10907 -11671
rect 10707 -11726 10907 -11688
rect 10965 -11688 11048 -11671
rect 11082 -11671 11098 -11654
rect 11896 -11654 11962 -11638
rect 11896 -11671 11912 -11654
rect 11082 -11688 11165 -11671
rect 10965 -11726 11165 -11688
rect 11829 -11688 11912 -11671
rect 11946 -11671 11962 -11654
rect 12154 -11654 12220 -11638
rect 12154 -11671 12170 -11654
rect 11946 -11688 12029 -11671
rect 11829 -11726 12029 -11688
rect 12087 -11688 12170 -11671
rect 12204 -11671 12220 -11654
rect 12412 -11654 12478 -11638
rect 12412 -11671 12428 -11654
rect 12204 -11688 12287 -11671
rect 12087 -11726 12287 -11688
rect 12345 -11688 12428 -11671
rect 12462 -11671 12478 -11654
rect 12670 -11654 12736 -11638
rect 12670 -11671 12686 -11654
rect 12462 -11688 12545 -11671
rect 12345 -11726 12545 -11688
rect 12603 -11688 12686 -11671
rect 12720 -11671 12736 -11654
rect 12928 -11654 12994 -11638
rect 12928 -11671 12944 -11654
rect 12720 -11688 12803 -11671
rect 12603 -11726 12803 -11688
rect 12861 -11688 12944 -11671
rect 12978 -11671 12994 -11654
rect 13186 -11654 13252 -11638
rect 13186 -11671 13202 -11654
rect 12978 -11688 13061 -11671
rect 12861 -11726 13061 -11688
rect 13119 -11688 13202 -11671
rect 13236 -11671 13252 -11654
rect 13444 -11654 13510 -11638
rect 13444 -11671 13460 -11654
rect 13236 -11688 13319 -11671
rect 13119 -11726 13319 -11688
rect 13377 -11688 13460 -11671
rect 13494 -11671 13510 -11654
rect 13702 -11654 13768 -11638
rect 13702 -11671 13718 -11654
rect 13494 -11688 13577 -11671
rect 13377 -11726 13577 -11688
rect 13635 -11688 13718 -11671
rect 13752 -11671 13768 -11654
rect 14559 -11653 14625 -11637
rect 14559 -11670 14575 -11653
rect 13752 -11688 13835 -11671
rect 13635 -11726 13835 -11688
rect 14492 -11687 14575 -11670
rect 14609 -11670 14625 -11653
rect 14817 -11653 14883 -11637
rect 14817 -11670 14833 -11653
rect 14609 -11687 14692 -11670
rect 14492 -11725 14692 -11687
rect 14750 -11687 14833 -11670
rect 14867 -11670 14883 -11653
rect 15075 -11653 15141 -11637
rect 15075 -11670 15091 -11653
rect 14867 -11687 14950 -11670
rect 14750 -11725 14950 -11687
rect 15008 -11687 15091 -11670
rect 15125 -11670 15141 -11653
rect 15333 -11653 15399 -11637
rect 15333 -11670 15349 -11653
rect 15125 -11687 15208 -11670
rect 15008 -11725 15208 -11687
rect 15266 -11687 15349 -11670
rect 15383 -11670 15399 -11653
rect 15591 -11653 15657 -11637
rect 15591 -11670 15607 -11653
rect 15383 -11687 15466 -11670
rect 15266 -11725 15466 -11687
rect 15524 -11687 15607 -11670
rect 15641 -11670 15657 -11653
rect 15849 -11653 15915 -11637
rect 15849 -11670 15865 -11653
rect 15641 -11687 15724 -11670
rect 15524 -11725 15724 -11687
rect 15782 -11687 15865 -11670
rect 15899 -11670 15915 -11653
rect 16107 -11653 16173 -11637
rect 16107 -11670 16123 -11653
rect 15899 -11687 15982 -11670
rect 15782 -11725 15982 -11687
rect 16040 -11687 16123 -11670
rect 16157 -11670 16173 -11653
rect 16365 -11653 16431 -11637
rect 16365 -11670 16381 -11653
rect 16157 -11687 16240 -11670
rect 16040 -11725 16240 -11687
rect 16298 -11687 16381 -11670
rect 16415 -11670 16431 -11653
rect 16415 -11687 16498 -11670
rect 16298 -11725 16498 -11687
rect 9159 -11964 9359 -11926
rect 9159 -11981 9242 -11964
rect 9226 -11998 9242 -11981
rect 9276 -11981 9359 -11964
rect 9417 -11964 9617 -11926
rect 9417 -11981 9500 -11964
rect 9276 -11998 9292 -11981
rect 9226 -12014 9292 -11998
rect 9484 -11998 9500 -11981
rect 9534 -11981 9617 -11964
rect 9675 -11964 9875 -11926
rect 9675 -11981 9758 -11964
rect 9534 -11998 9550 -11981
rect 9484 -12014 9550 -11998
rect 9742 -11998 9758 -11981
rect 9792 -11981 9875 -11964
rect 9933 -11964 10133 -11926
rect 9933 -11981 10016 -11964
rect 9792 -11998 9808 -11981
rect 9742 -12014 9808 -11998
rect 10000 -11998 10016 -11981
rect 10050 -11981 10133 -11964
rect 10191 -11964 10391 -11926
rect 10191 -11981 10274 -11964
rect 10050 -11998 10066 -11981
rect 10000 -12014 10066 -11998
rect 10258 -11998 10274 -11981
rect 10308 -11981 10391 -11964
rect 10449 -11964 10649 -11926
rect 10449 -11981 10532 -11964
rect 10308 -11998 10324 -11981
rect 10258 -12014 10324 -11998
rect 10516 -11998 10532 -11981
rect 10566 -11981 10649 -11964
rect 10707 -11964 10907 -11926
rect 10707 -11981 10790 -11964
rect 10566 -11998 10582 -11981
rect 10516 -12014 10582 -11998
rect 10774 -11998 10790 -11981
rect 10824 -11981 10907 -11964
rect 10965 -11964 11165 -11926
rect 10965 -11981 11048 -11964
rect 10824 -11998 10840 -11981
rect 10774 -12014 10840 -11998
rect 11032 -11998 11048 -11981
rect 11082 -11981 11165 -11964
rect 11829 -11964 12029 -11926
rect 11829 -11981 11912 -11964
rect 11082 -11998 11098 -11981
rect 11032 -12014 11098 -11998
rect 11896 -11998 11912 -11981
rect 11946 -11981 12029 -11964
rect 12087 -11964 12287 -11926
rect 12087 -11981 12170 -11964
rect 11946 -11998 11962 -11981
rect 11896 -12014 11962 -11998
rect 12154 -11998 12170 -11981
rect 12204 -11981 12287 -11964
rect 12345 -11964 12545 -11926
rect 12345 -11981 12428 -11964
rect 12204 -11998 12220 -11981
rect 12154 -12014 12220 -11998
rect 12412 -11998 12428 -11981
rect 12462 -11981 12545 -11964
rect 12603 -11964 12803 -11926
rect 12603 -11981 12686 -11964
rect 12462 -11998 12478 -11981
rect 12412 -12014 12478 -11998
rect 12670 -11998 12686 -11981
rect 12720 -11981 12803 -11964
rect 12861 -11964 13061 -11926
rect 12861 -11981 12944 -11964
rect 12720 -11998 12736 -11981
rect 12670 -12014 12736 -11998
rect 12928 -11998 12944 -11981
rect 12978 -11981 13061 -11964
rect 13119 -11964 13319 -11926
rect 13119 -11981 13202 -11964
rect 12978 -11998 12994 -11981
rect 12928 -12014 12994 -11998
rect 13186 -11998 13202 -11981
rect 13236 -11981 13319 -11964
rect 13377 -11964 13577 -11926
rect 13377 -11981 13460 -11964
rect 13236 -11998 13252 -11981
rect 13186 -12014 13252 -11998
rect 13444 -11998 13460 -11981
rect 13494 -11981 13577 -11964
rect 13635 -11964 13835 -11926
rect 13635 -11981 13718 -11964
rect 13494 -11998 13510 -11981
rect 13444 -12014 13510 -11998
rect 13702 -11998 13718 -11981
rect 13752 -11981 13835 -11964
rect 14492 -11963 14692 -11925
rect 14492 -11980 14575 -11963
rect 13752 -11998 13768 -11981
rect 13702 -12014 13768 -11998
rect 14559 -11997 14575 -11980
rect 14609 -11980 14692 -11963
rect 14750 -11963 14950 -11925
rect 14750 -11980 14833 -11963
rect 14609 -11997 14625 -11980
rect 14559 -12013 14625 -11997
rect 14817 -11997 14833 -11980
rect 14867 -11980 14950 -11963
rect 15008 -11963 15208 -11925
rect 15008 -11980 15091 -11963
rect 14867 -11997 14883 -11980
rect 14817 -12013 14883 -11997
rect 15075 -11997 15091 -11980
rect 15125 -11980 15208 -11963
rect 15266 -11963 15466 -11925
rect 15266 -11980 15349 -11963
rect 15125 -11997 15141 -11980
rect 15075 -12013 15141 -11997
rect 15333 -11997 15349 -11980
rect 15383 -11980 15466 -11963
rect 15524 -11963 15724 -11925
rect 15524 -11980 15607 -11963
rect 15383 -11997 15399 -11980
rect 15333 -12013 15399 -11997
rect 15591 -11997 15607 -11980
rect 15641 -11980 15724 -11963
rect 15782 -11963 15982 -11925
rect 15782 -11980 15865 -11963
rect 15641 -11997 15657 -11980
rect 15591 -12013 15657 -11997
rect 15849 -11997 15865 -11980
rect 15899 -11980 15982 -11963
rect 16040 -11963 16240 -11925
rect 16040 -11980 16123 -11963
rect 15899 -11997 15915 -11980
rect 15849 -12013 15915 -11997
rect 16107 -11997 16123 -11980
rect 16157 -11980 16240 -11963
rect 16298 -11963 16498 -11925
rect 16298 -11980 16381 -11963
rect 16157 -11997 16173 -11980
rect 16107 -12013 16173 -11997
rect 16365 -11997 16381 -11980
rect 16415 -11980 16498 -11963
rect 16415 -11997 16431 -11980
rect 16365 -12013 16431 -11997
rect 9226 -12072 9292 -12056
rect 9226 -12089 9242 -12072
rect 9159 -12106 9242 -12089
rect 9276 -12089 9292 -12072
rect 9484 -12072 9550 -12056
rect 9484 -12089 9500 -12072
rect 9276 -12106 9359 -12089
rect 9159 -12144 9359 -12106
rect 9417 -12106 9500 -12089
rect 9534 -12089 9550 -12072
rect 9742 -12072 9808 -12056
rect 9742 -12089 9758 -12072
rect 9534 -12106 9617 -12089
rect 9417 -12144 9617 -12106
rect 9675 -12106 9758 -12089
rect 9792 -12089 9808 -12072
rect 10000 -12072 10066 -12056
rect 10000 -12089 10016 -12072
rect 9792 -12106 9875 -12089
rect 9675 -12144 9875 -12106
rect 9933 -12106 10016 -12089
rect 10050 -12089 10066 -12072
rect 10258 -12072 10324 -12056
rect 10258 -12089 10274 -12072
rect 10050 -12106 10133 -12089
rect 9933 -12144 10133 -12106
rect 10191 -12106 10274 -12089
rect 10308 -12089 10324 -12072
rect 10516 -12072 10582 -12056
rect 10516 -12089 10532 -12072
rect 10308 -12106 10391 -12089
rect 10191 -12144 10391 -12106
rect 10449 -12106 10532 -12089
rect 10566 -12089 10582 -12072
rect 10774 -12072 10840 -12056
rect 10774 -12089 10790 -12072
rect 10566 -12106 10649 -12089
rect 10449 -12144 10649 -12106
rect 10707 -12106 10790 -12089
rect 10824 -12089 10840 -12072
rect 11032 -12072 11098 -12056
rect 11032 -12089 11048 -12072
rect 10824 -12106 10907 -12089
rect 10707 -12144 10907 -12106
rect 10965 -12106 11048 -12089
rect 11082 -12089 11098 -12072
rect 11896 -12072 11962 -12056
rect 11896 -12089 11912 -12072
rect 11082 -12106 11165 -12089
rect 10965 -12144 11165 -12106
rect 11829 -12106 11912 -12089
rect 11946 -12089 11962 -12072
rect 12154 -12072 12220 -12056
rect 12154 -12089 12170 -12072
rect 11946 -12106 12029 -12089
rect 11829 -12144 12029 -12106
rect 12087 -12106 12170 -12089
rect 12204 -12089 12220 -12072
rect 12412 -12072 12478 -12056
rect 12412 -12089 12428 -12072
rect 12204 -12106 12287 -12089
rect 12087 -12144 12287 -12106
rect 12345 -12106 12428 -12089
rect 12462 -12089 12478 -12072
rect 12670 -12072 12736 -12056
rect 12670 -12089 12686 -12072
rect 12462 -12106 12545 -12089
rect 12345 -12144 12545 -12106
rect 12603 -12106 12686 -12089
rect 12720 -12089 12736 -12072
rect 12928 -12072 12994 -12056
rect 12928 -12089 12944 -12072
rect 12720 -12106 12803 -12089
rect 12603 -12144 12803 -12106
rect 12861 -12106 12944 -12089
rect 12978 -12089 12994 -12072
rect 13186 -12072 13252 -12056
rect 13186 -12089 13202 -12072
rect 12978 -12106 13061 -12089
rect 12861 -12144 13061 -12106
rect 13119 -12106 13202 -12089
rect 13236 -12089 13252 -12072
rect 13444 -12072 13510 -12056
rect 13444 -12089 13460 -12072
rect 13236 -12106 13319 -12089
rect 13119 -12144 13319 -12106
rect 13377 -12106 13460 -12089
rect 13494 -12089 13510 -12072
rect 13702 -12072 13768 -12056
rect 13702 -12089 13718 -12072
rect 13494 -12106 13577 -12089
rect 13377 -12144 13577 -12106
rect 13635 -12106 13718 -12089
rect 13752 -12089 13768 -12072
rect 14559 -12071 14625 -12055
rect 14559 -12088 14575 -12071
rect 13752 -12106 13835 -12089
rect 13635 -12144 13835 -12106
rect 14492 -12105 14575 -12088
rect 14609 -12088 14625 -12071
rect 14817 -12071 14883 -12055
rect 14817 -12088 14833 -12071
rect 14609 -12105 14692 -12088
rect 14492 -12143 14692 -12105
rect 14750 -12105 14833 -12088
rect 14867 -12088 14883 -12071
rect 15075 -12071 15141 -12055
rect 15075 -12088 15091 -12071
rect 14867 -12105 14950 -12088
rect 14750 -12143 14950 -12105
rect 15008 -12105 15091 -12088
rect 15125 -12088 15141 -12071
rect 15333 -12071 15399 -12055
rect 15333 -12088 15349 -12071
rect 15125 -12105 15208 -12088
rect 15008 -12143 15208 -12105
rect 15266 -12105 15349 -12088
rect 15383 -12088 15399 -12071
rect 15591 -12071 15657 -12055
rect 15591 -12088 15607 -12071
rect 15383 -12105 15466 -12088
rect 15266 -12143 15466 -12105
rect 15524 -12105 15607 -12088
rect 15641 -12088 15657 -12071
rect 15849 -12071 15915 -12055
rect 15849 -12088 15865 -12071
rect 15641 -12105 15724 -12088
rect 15524 -12143 15724 -12105
rect 15782 -12105 15865 -12088
rect 15899 -12088 15915 -12071
rect 16107 -12071 16173 -12055
rect 16107 -12088 16123 -12071
rect 15899 -12105 15982 -12088
rect 15782 -12143 15982 -12105
rect 16040 -12105 16123 -12088
rect 16157 -12088 16173 -12071
rect 16365 -12071 16431 -12055
rect 16365 -12088 16381 -12071
rect 16157 -12105 16240 -12088
rect 16040 -12143 16240 -12105
rect 16298 -12105 16381 -12088
rect 16415 -12088 16431 -12071
rect 16415 -12105 16498 -12088
rect 16298 -12143 16498 -12105
rect 9159 -12382 9359 -12344
rect 9159 -12399 9242 -12382
rect 9226 -12416 9242 -12399
rect 9276 -12399 9359 -12382
rect 9417 -12382 9617 -12344
rect 9417 -12399 9500 -12382
rect 9276 -12416 9292 -12399
rect 9226 -12432 9292 -12416
rect 9484 -12416 9500 -12399
rect 9534 -12399 9617 -12382
rect 9675 -12382 9875 -12344
rect 9675 -12399 9758 -12382
rect 9534 -12416 9550 -12399
rect 9484 -12432 9550 -12416
rect 9742 -12416 9758 -12399
rect 9792 -12399 9875 -12382
rect 9933 -12382 10133 -12344
rect 9933 -12399 10016 -12382
rect 9792 -12416 9808 -12399
rect 9742 -12432 9808 -12416
rect 10000 -12416 10016 -12399
rect 10050 -12399 10133 -12382
rect 10191 -12382 10391 -12344
rect 10191 -12399 10274 -12382
rect 10050 -12416 10066 -12399
rect 10000 -12432 10066 -12416
rect 10258 -12416 10274 -12399
rect 10308 -12399 10391 -12382
rect 10449 -12382 10649 -12344
rect 10449 -12399 10532 -12382
rect 10308 -12416 10324 -12399
rect 10258 -12432 10324 -12416
rect 10516 -12416 10532 -12399
rect 10566 -12399 10649 -12382
rect 10707 -12382 10907 -12344
rect 10707 -12399 10790 -12382
rect 10566 -12416 10582 -12399
rect 10516 -12432 10582 -12416
rect 10774 -12416 10790 -12399
rect 10824 -12399 10907 -12382
rect 10965 -12382 11165 -12344
rect 10965 -12399 11048 -12382
rect 10824 -12416 10840 -12399
rect 10774 -12432 10840 -12416
rect 11032 -12416 11048 -12399
rect 11082 -12399 11165 -12382
rect 11829 -12382 12029 -12344
rect 11829 -12399 11912 -12382
rect 11082 -12416 11098 -12399
rect 11032 -12432 11098 -12416
rect 11896 -12416 11912 -12399
rect 11946 -12399 12029 -12382
rect 12087 -12382 12287 -12344
rect 12087 -12399 12170 -12382
rect 11946 -12416 11962 -12399
rect 11896 -12432 11962 -12416
rect 12154 -12416 12170 -12399
rect 12204 -12399 12287 -12382
rect 12345 -12382 12545 -12344
rect 12345 -12399 12428 -12382
rect 12204 -12416 12220 -12399
rect 12154 -12432 12220 -12416
rect 12412 -12416 12428 -12399
rect 12462 -12399 12545 -12382
rect 12603 -12382 12803 -12344
rect 12603 -12399 12686 -12382
rect 12462 -12416 12478 -12399
rect 12412 -12432 12478 -12416
rect 12670 -12416 12686 -12399
rect 12720 -12399 12803 -12382
rect 12861 -12382 13061 -12344
rect 12861 -12399 12944 -12382
rect 12720 -12416 12736 -12399
rect 12670 -12432 12736 -12416
rect 12928 -12416 12944 -12399
rect 12978 -12399 13061 -12382
rect 13119 -12382 13319 -12344
rect 13119 -12399 13202 -12382
rect 12978 -12416 12994 -12399
rect 12928 -12432 12994 -12416
rect 13186 -12416 13202 -12399
rect 13236 -12399 13319 -12382
rect 13377 -12382 13577 -12344
rect 13377 -12399 13460 -12382
rect 13236 -12416 13252 -12399
rect 13186 -12432 13252 -12416
rect 13444 -12416 13460 -12399
rect 13494 -12399 13577 -12382
rect 13635 -12382 13835 -12344
rect 13635 -12399 13718 -12382
rect 13494 -12416 13510 -12399
rect 13444 -12432 13510 -12416
rect 13702 -12416 13718 -12399
rect 13752 -12399 13835 -12382
rect 14492 -12381 14692 -12343
rect 14492 -12398 14575 -12381
rect 13752 -12416 13768 -12399
rect 13702 -12432 13768 -12416
rect 14559 -12415 14575 -12398
rect 14609 -12398 14692 -12381
rect 14750 -12381 14950 -12343
rect 14750 -12398 14833 -12381
rect 14609 -12415 14625 -12398
rect 14559 -12431 14625 -12415
rect 14817 -12415 14833 -12398
rect 14867 -12398 14950 -12381
rect 15008 -12381 15208 -12343
rect 15008 -12398 15091 -12381
rect 14867 -12415 14883 -12398
rect 14817 -12431 14883 -12415
rect 15075 -12415 15091 -12398
rect 15125 -12398 15208 -12381
rect 15266 -12381 15466 -12343
rect 15266 -12398 15349 -12381
rect 15125 -12415 15141 -12398
rect 15075 -12431 15141 -12415
rect 15333 -12415 15349 -12398
rect 15383 -12398 15466 -12381
rect 15524 -12381 15724 -12343
rect 15524 -12398 15607 -12381
rect 15383 -12415 15399 -12398
rect 15333 -12431 15399 -12415
rect 15591 -12415 15607 -12398
rect 15641 -12398 15724 -12381
rect 15782 -12381 15982 -12343
rect 15782 -12398 15865 -12381
rect 15641 -12415 15657 -12398
rect 15591 -12431 15657 -12415
rect 15849 -12415 15865 -12398
rect 15899 -12398 15982 -12381
rect 16040 -12381 16240 -12343
rect 16040 -12398 16123 -12381
rect 15899 -12415 15915 -12398
rect 15849 -12431 15915 -12415
rect 16107 -12415 16123 -12398
rect 16157 -12398 16240 -12381
rect 16298 -12381 16498 -12343
rect 16298 -12398 16381 -12381
rect 16157 -12415 16173 -12398
rect 16107 -12431 16173 -12415
rect 16365 -12415 16381 -12398
rect 16415 -12398 16498 -12381
rect 16415 -12415 16431 -12398
rect 16365 -12431 16431 -12415
rect 9106 -12724 9172 -12708
rect 9106 -12741 9122 -12724
rect 9039 -12758 9122 -12741
rect 9156 -12741 9172 -12724
rect 9646 -12724 9712 -12708
rect 9646 -12741 9662 -12724
rect 9156 -12758 9239 -12741
rect 9039 -12796 9239 -12758
rect 9579 -12758 9662 -12741
rect 9696 -12741 9712 -12724
rect 10126 -12724 10192 -12708
rect 10126 -12741 10142 -12724
rect 9696 -12758 9779 -12741
rect 9579 -12796 9779 -12758
rect 10059 -12758 10142 -12741
rect 10176 -12741 10192 -12724
rect 10629 -12722 10695 -12706
rect 10629 -12739 10645 -12722
rect 10176 -12758 10259 -12741
rect 10059 -12796 10259 -12758
rect 10562 -12756 10645 -12739
rect 10679 -12739 10695 -12722
rect 11139 -12712 11205 -12696
rect 11139 -12729 11155 -12712
rect 10679 -12756 10762 -12739
rect 10562 -12794 10762 -12756
rect 11072 -12746 11155 -12729
rect 11189 -12729 11205 -12712
rect 11776 -12724 11842 -12708
rect 11189 -12746 11272 -12729
rect 11776 -12741 11792 -12724
rect 11072 -12784 11272 -12746
rect 11709 -12758 11792 -12741
rect 11826 -12741 11842 -12724
rect 12316 -12724 12382 -12708
rect 12316 -12741 12332 -12724
rect 11826 -12758 11909 -12741
rect 11709 -12796 11909 -12758
rect 12249 -12758 12332 -12741
rect 12366 -12741 12382 -12724
rect 12796 -12724 12862 -12708
rect 12796 -12741 12812 -12724
rect 12366 -12758 12449 -12741
rect 12249 -12796 12449 -12758
rect 12729 -12758 12812 -12741
rect 12846 -12741 12862 -12724
rect 13299 -12722 13365 -12706
rect 13299 -12739 13315 -12722
rect 12846 -12758 12929 -12741
rect 12729 -12796 12929 -12758
rect 13232 -12756 13315 -12739
rect 13349 -12739 13365 -12722
rect 13809 -12712 13875 -12696
rect 13809 -12729 13825 -12712
rect 13349 -12756 13432 -12739
rect 13232 -12794 13432 -12756
rect 13742 -12746 13825 -12729
rect 13859 -12729 13875 -12712
rect 14439 -12723 14505 -12707
rect 13859 -12746 13942 -12729
rect 14439 -12740 14455 -12723
rect 13742 -12784 13942 -12746
rect 14372 -12757 14455 -12740
rect 14489 -12740 14505 -12723
rect 14979 -12723 15045 -12707
rect 14979 -12740 14995 -12723
rect 14489 -12757 14572 -12740
rect 9039 -13034 9239 -12996
rect 9039 -13051 9122 -13034
rect 9106 -13068 9122 -13051
rect 9156 -13051 9239 -13034
rect 9579 -13034 9779 -12996
rect 9579 -13051 9662 -13034
rect 9156 -13068 9172 -13051
rect 9106 -13084 9172 -13068
rect 9646 -13068 9662 -13051
rect 9696 -13051 9779 -13034
rect 10059 -13034 10259 -12996
rect 10059 -13051 10142 -13034
rect 9696 -13068 9712 -13051
rect 9646 -13084 9712 -13068
rect 10126 -13068 10142 -13051
rect 10176 -13051 10259 -13034
rect 10562 -13032 10762 -12994
rect 10562 -13049 10645 -13032
rect 10176 -13068 10192 -13051
rect 10126 -13084 10192 -13068
rect 10629 -13066 10645 -13049
rect 10679 -13049 10762 -13032
rect 11072 -13022 11272 -12984
rect 14372 -12795 14572 -12757
rect 14912 -12757 14995 -12740
rect 15029 -12740 15045 -12723
rect 15459 -12723 15525 -12707
rect 15459 -12740 15475 -12723
rect 15029 -12757 15112 -12740
rect 14912 -12795 15112 -12757
rect 15392 -12757 15475 -12740
rect 15509 -12740 15525 -12723
rect 15962 -12721 16028 -12705
rect 15962 -12738 15978 -12721
rect 15509 -12757 15592 -12740
rect 15392 -12795 15592 -12757
rect 15895 -12755 15978 -12738
rect 16012 -12738 16028 -12721
rect 16472 -12711 16538 -12695
rect 16472 -12728 16488 -12711
rect 16012 -12755 16095 -12738
rect 15895 -12793 16095 -12755
rect 16405 -12745 16488 -12728
rect 16522 -12728 16538 -12711
rect 16522 -12745 16605 -12728
rect 16405 -12783 16605 -12745
rect 11072 -13039 11155 -13022
rect 10679 -13066 10695 -13049
rect 10629 -13082 10695 -13066
rect 11139 -13056 11155 -13039
rect 11189 -13039 11272 -13022
rect 11709 -13034 11909 -12996
rect 11189 -13056 11205 -13039
rect 11709 -13051 11792 -13034
rect 11139 -13072 11205 -13056
rect 11776 -13068 11792 -13051
rect 11826 -13051 11909 -13034
rect 12249 -13034 12449 -12996
rect 12249 -13051 12332 -13034
rect 11826 -13068 11842 -13051
rect 11776 -13084 11842 -13068
rect 12316 -13068 12332 -13051
rect 12366 -13051 12449 -13034
rect 12729 -13034 12929 -12996
rect 12729 -13051 12812 -13034
rect 12366 -13068 12382 -13051
rect 12316 -13084 12382 -13068
rect 12796 -13068 12812 -13051
rect 12846 -13051 12929 -13034
rect 13232 -13032 13432 -12994
rect 13232 -13049 13315 -13032
rect 12846 -13068 12862 -13051
rect 12796 -13084 12862 -13068
rect 13299 -13066 13315 -13049
rect 13349 -13049 13432 -13032
rect 13742 -13022 13942 -12984
rect 13742 -13039 13825 -13022
rect 13349 -13066 13365 -13049
rect 13299 -13082 13365 -13066
rect 13809 -13056 13825 -13039
rect 13859 -13039 13942 -13022
rect 14372 -13033 14572 -12995
rect 13859 -13056 13875 -13039
rect 14372 -13050 14455 -13033
rect 13809 -13072 13875 -13056
rect 14439 -13067 14455 -13050
rect 14489 -13050 14572 -13033
rect 14912 -13033 15112 -12995
rect 14912 -13050 14995 -13033
rect 14489 -13067 14505 -13050
rect 14439 -13083 14505 -13067
rect 14979 -13067 14995 -13050
rect 15029 -13050 15112 -13033
rect 15392 -13033 15592 -12995
rect 15392 -13050 15475 -13033
rect 15029 -13067 15045 -13050
rect 14979 -13083 15045 -13067
rect 15459 -13067 15475 -13050
rect 15509 -13050 15592 -13033
rect 15895 -13031 16095 -12993
rect 15895 -13048 15978 -13031
rect 15509 -13067 15525 -13050
rect 15459 -13083 15525 -13067
rect 15962 -13065 15978 -13048
rect 16012 -13048 16095 -13031
rect 16405 -13021 16605 -12983
rect 16405 -13038 16488 -13021
rect 16012 -13065 16028 -13048
rect 15962 -13081 16028 -13065
rect 16472 -13055 16488 -13038
rect 16522 -13038 16605 -13021
rect 16522 -13055 16538 -13038
rect 16472 -13071 16538 -13055
rect 9384 -14243 9500 -14215
rect 9384 -14281 9408 -14243
rect 9474 -14281 9500 -14243
rect 10036 -14250 10222 -14234
rect 10036 -14267 10052 -14250
rect 9384 -14331 9500 -14281
rect 9729 -14284 10052 -14267
rect 10206 -14267 10222 -14250
rect 10770 -14244 10886 -14216
rect 10206 -14284 10529 -14267
rect 9729 -14331 10529 -14284
rect 10770 -14282 10794 -14244
rect 10860 -14282 10886 -14244
rect 10770 -14332 10886 -14282
rect 11140 -14244 11256 -14216
rect 11140 -14282 11164 -14244
rect 11230 -14282 11256 -14244
rect 11140 -14332 11256 -14282
rect 11562 -14244 11678 -14216
rect 11562 -14282 11586 -14244
rect 11652 -14282 11678 -14244
rect 11562 -14332 11678 -14282
rect 11984 -14244 12100 -14216
rect 11984 -14282 12008 -14244
rect 12074 -14282 12100 -14244
rect 12713 -14250 12899 -14234
rect 12713 -14267 12729 -14250
rect 11984 -14332 12100 -14282
rect 12406 -14284 12729 -14267
rect 12883 -14267 12899 -14250
rect 13484 -14240 13600 -14212
rect 12883 -14284 13206 -14267
rect 12406 -14331 13206 -14284
rect 13484 -14278 13508 -14240
rect 13574 -14278 13600 -14240
rect 13484 -14328 13600 -14278
rect 13854 -14240 13970 -14212
rect 13854 -14278 13878 -14240
rect 13944 -14278 13970 -14240
rect 13854 -14328 13970 -14278
rect 14276 -14240 14392 -14212
rect 14276 -14278 14300 -14240
rect 14366 -14278 14392 -14240
rect 14276 -14328 14392 -14278
rect 14698 -14240 14814 -14212
rect 14698 -14278 14722 -14240
rect 14788 -14278 14814 -14240
rect 15377 -14249 15563 -14233
rect 15377 -14266 15393 -14249
rect 14698 -14328 14814 -14278
rect 15070 -14283 15393 -14266
rect 15547 -14266 15563 -14249
rect 16082 -14243 16198 -14215
rect 15547 -14283 15870 -14266
rect 9384 -14505 9500 -14441
rect 9729 -14488 10529 -14441
rect 15070 -14330 15870 -14283
rect 16082 -14281 16106 -14243
rect 16172 -14281 16198 -14243
rect 9729 -14505 10052 -14488
rect 10036 -14522 10052 -14505
rect 10206 -14505 10529 -14488
rect 10206 -14522 10222 -14505
rect 10770 -14506 10886 -14442
rect 11140 -14506 11256 -14442
rect 11562 -14506 11678 -14442
rect 11984 -14506 12100 -14442
rect 12406 -14488 13206 -14441
rect 12406 -14505 12729 -14488
rect 10036 -14538 10222 -14522
rect 12713 -14522 12729 -14505
rect 12883 -14505 13206 -14488
rect 13484 -14502 13600 -14438
rect 13854 -14502 13970 -14438
rect 14276 -14502 14392 -14438
rect 14698 -14502 14814 -14438
rect 16082 -14331 16198 -14281
rect 15070 -14487 15870 -14440
rect 15070 -14504 15393 -14487
rect 12883 -14522 12899 -14505
rect 12713 -14538 12899 -14522
rect 15377 -14521 15393 -14504
rect 15547 -14504 15870 -14487
rect 15547 -14521 15563 -14504
rect 16082 -14505 16198 -14441
rect 15377 -14537 15563 -14521
rect 9226 -15281 9292 -15265
rect 9226 -15298 9242 -15281
rect 9159 -15315 9242 -15298
rect 9276 -15298 9292 -15281
rect 9484 -15281 9550 -15265
rect 9484 -15298 9500 -15281
rect 9276 -15315 9359 -15298
rect 9159 -15353 9359 -15315
rect 9417 -15315 9500 -15298
rect 9534 -15298 9550 -15281
rect 9742 -15281 9808 -15265
rect 9742 -15298 9758 -15281
rect 9534 -15315 9617 -15298
rect 9417 -15353 9617 -15315
rect 9675 -15315 9758 -15298
rect 9792 -15298 9808 -15281
rect 10000 -15281 10066 -15265
rect 10000 -15298 10016 -15281
rect 9792 -15315 9875 -15298
rect 9675 -15353 9875 -15315
rect 9933 -15315 10016 -15298
rect 10050 -15298 10066 -15281
rect 10258 -15281 10324 -15265
rect 10258 -15298 10274 -15281
rect 10050 -15315 10133 -15298
rect 9933 -15353 10133 -15315
rect 10191 -15315 10274 -15298
rect 10308 -15298 10324 -15281
rect 10516 -15281 10582 -15265
rect 10516 -15298 10532 -15281
rect 10308 -15315 10391 -15298
rect 10191 -15353 10391 -15315
rect 10449 -15315 10532 -15298
rect 10566 -15298 10582 -15281
rect 10774 -15281 10840 -15265
rect 10774 -15298 10790 -15281
rect 10566 -15315 10649 -15298
rect 10449 -15353 10649 -15315
rect 10707 -15315 10790 -15298
rect 10824 -15298 10840 -15281
rect 11032 -15281 11098 -15265
rect 11032 -15298 11048 -15281
rect 10824 -15315 10907 -15298
rect 10707 -15353 10907 -15315
rect 10965 -15315 11048 -15298
rect 11082 -15298 11098 -15281
rect 11896 -15281 11962 -15265
rect 11896 -15298 11912 -15281
rect 11082 -15315 11165 -15298
rect 10965 -15353 11165 -15315
rect 11829 -15315 11912 -15298
rect 11946 -15298 11962 -15281
rect 12154 -15281 12220 -15265
rect 12154 -15298 12170 -15281
rect 11946 -15315 12029 -15298
rect 11829 -15353 12029 -15315
rect 12087 -15315 12170 -15298
rect 12204 -15298 12220 -15281
rect 12412 -15281 12478 -15265
rect 12412 -15298 12428 -15281
rect 12204 -15315 12287 -15298
rect 12087 -15353 12287 -15315
rect 12345 -15315 12428 -15298
rect 12462 -15298 12478 -15281
rect 12670 -15281 12736 -15265
rect 12670 -15298 12686 -15281
rect 12462 -15315 12545 -15298
rect 12345 -15353 12545 -15315
rect 12603 -15315 12686 -15298
rect 12720 -15298 12736 -15281
rect 12928 -15281 12994 -15265
rect 12928 -15298 12944 -15281
rect 12720 -15315 12803 -15298
rect 12603 -15353 12803 -15315
rect 12861 -15315 12944 -15298
rect 12978 -15298 12994 -15281
rect 13186 -15281 13252 -15265
rect 13186 -15298 13202 -15281
rect 12978 -15315 13061 -15298
rect 12861 -15353 13061 -15315
rect 13119 -15315 13202 -15298
rect 13236 -15298 13252 -15281
rect 13444 -15281 13510 -15265
rect 13444 -15298 13460 -15281
rect 13236 -15315 13319 -15298
rect 13119 -15353 13319 -15315
rect 13377 -15315 13460 -15298
rect 13494 -15298 13510 -15281
rect 13702 -15281 13768 -15265
rect 13702 -15298 13718 -15281
rect 13494 -15315 13577 -15298
rect 13377 -15353 13577 -15315
rect 13635 -15315 13718 -15298
rect 13752 -15298 13768 -15281
rect 14559 -15280 14625 -15264
rect 14559 -15297 14575 -15280
rect 13752 -15315 13835 -15298
rect 13635 -15353 13835 -15315
rect 14492 -15314 14575 -15297
rect 14609 -15297 14625 -15280
rect 14817 -15280 14883 -15264
rect 14817 -15297 14833 -15280
rect 14609 -15314 14692 -15297
rect 14492 -15352 14692 -15314
rect 14750 -15314 14833 -15297
rect 14867 -15297 14883 -15280
rect 15075 -15280 15141 -15264
rect 15075 -15297 15091 -15280
rect 14867 -15314 14950 -15297
rect 14750 -15352 14950 -15314
rect 15008 -15314 15091 -15297
rect 15125 -15297 15141 -15280
rect 15333 -15280 15399 -15264
rect 15333 -15297 15349 -15280
rect 15125 -15314 15208 -15297
rect 15008 -15352 15208 -15314
rect 15266 -15314 15349 -15297
rect 15383 -15297 15399 -15280
rect 15591 -15280 15657 -15264
rect 15591 -15297 15607 -15280
rect 15383 -15314 15466 -15297
rect 15266 -15352 15466 -15314
rect 15524 -15314 15607 -15297
rect 15641 -15297 15657 -15280
rect 15849 -15280 15915 -15264
rect 15849 -15297 15865 -15280
rect 15641 -15314 15724 -15297
rect 15524 -15352 15724 -15314
rect 15782 -15314 15865 -15297
rect 15899 -15297 15915 -15280
rect 16107 -15280 16173 -15264
rect 16107 -15297 16123 -15280
rect 15899 -15314 15982 -15297
rect 15782 -15352 15982 -15314
rect 16040 -15314 16123 -15297
rect 16157 -15297 16173 -15280
rect 16365 -15280 16431 -15264
rect 16365 -15297 16381 -15280
rect 16157 -15314 16240 -15297
rect 16040 -15352 16240 -15314
rect 16298 -15314 16381 -15297
rect 16415 -15297 16431 -15280
rect 16415 -15314 16498 -15297
rect 16298 -15352 16498 -15314
rect 9159 -15591 9359 -15553
rect 9159 -15608 9242 -15591
rect 9226 -15625 9242 -15608
rect 9276 -15608 9359 -15591
rect 9417 -15591 9617 -15553
rect 9417 -15608 9500 -15591
rect 9276 -15625 9292 -15608
rect 9226 -15641 9292 -15625
rect 9484 -15625 9500 -15608
rect 9534 -15608 9617 -15591
rect 9675 -15591 9875 -15553
rect 9675 -15608 9758 -15591
rect 9534 -15625 9550 -15608
rect 9484 -15641 9550 -15625
rect 9742 -15625 9758 -15608
rect 9792 -15608 9875 -15591
rect 9933 -15591 10133 -15553
rect 9933 -15608 10016 -15591
rect 9792 -15625 9808 -15608
rect 9742 -15641 9808 -15625
rect 10000 -15625 10016 -15608
rect 10050 -15608 10133 -15591
rect 10191 -15591 10391 -15553
rect 10191 -15608 10274 -15591
rect 10050 -15625 10066 -15608
rect 10000 -15641 10066 -15625
rect 10258 -15625 10274 -15608
rect 10308 -15608 10391 -15591
rect 10449 -15591 10649 -15553
rect 10449 -15608 10532 -15591
rect 10308 -15625 10324 -15608
rect 10258 -15641 10324 -15625
rect 10516 -15625 10532 -15608
rect 10566 -15608 10649 -15591
rect 10707 -15591 10907 -15553
rect 10707 -15608 10790 -15591
rect 10566 -15625 10582 -15608
rect 10516 -15641 10582 -15625
rect 10774 -15625 10790 -15608
rect 10824 -15608 10907 -15591
rect 10965 -15591 11165 -15553
rect 10965 -15608 11048 -15591
rect 10824 -15625 10840 -15608
rect 10774 -15641 10840 -15625
rect 11032 -15625 11048 -15608
rect 11082 -15608 11165 -15591
rect 11829 -15591 12029 -15553
rect 11829 -15608 11912 -15591
rect 11082 -15625 11098 -15608
rect 11032 -15641 11098 -15625
rect 11896 -15625 11912 -15608
rect 11946 -15608 12029 -15591
rect 12087 -15591 12287 -15553
rect 12087 -15608 12170 -15591
rect 11946 -15625 11962 -15608
rect 11896 -15641 11962 -15625
rect 12154 -15625 12170 -15608
rect 12204 -15608 12287 -15591
rect 12345 -15591 12545 -15553
rect 12345 -15608 12428 -15591
rect 12204 -15625 12220 -15608
rect 12154 -15641 12220 -15625
rect 12412 -15625 12428 -15608
rect 12462 -15608 12545 -15591
rect 12603 -15591 12803 -15553
rect 12603 -15608 12686 -15591
rect 12462 -15625 12478 -15608
rect 12412 -15641 12478 -15625
rect 12670 -15625 12686 -15608
rect 12720 -15608 12803 -15591
rect 12861 -15591 13061 -15553
rect 12861 -15608 12944 -15591
rect 12720 -15625 12736 -15608
rect 12670 -15641 12736 -15625
rect 12928 -15625 12944 -15608
rect 12978 -15608 13061 -15591
rect 13119 -15591 13319 -15553
rect 13119 -15608 13202 -15591
rect 12978 -15625 12994 -15608
rect 12928 -15641 12994 -15625
rect 13186 -15625 13202 -15608
rect 13236 -15608 13319 -15591
rect 13377 -15591 13577 -15553
rect 13377 -15608 13460 -15591
rect 13236 -15625 13252 -15608
rect 13186 -15641 13252 -15625
rect 13444 -15625 13460 -15608
rect 13494 -15608 13577 -15591
rect 13635 -15591 13835 -15553
rect 13635 -15608 13718 -15591
rect 13494 -15625 13510 -15608
rect 13444 -15641 13510 -15625
rect 13702 -15625 13718 -15608
rect 13752 -15608 13835 -15591
rect 14492 -15590 14692 -15552
rect 14492 -15607 14575 -15590
rect 13752 -15625 13768 -15608
rect 13702 -15641 13768 -15625
rect 14559 -15624 14575 -15607
rect 14609 -15607 14692 -15590
rect 14750 -15590 14950 -15552
rect 14750 -15607 14833 -15590
rect 14609 -15624 14625 -15607
rect 14559 -15640 14625 -15624
rect 14817 -15624 14833 -15607
rect 14867 -15607 14950 -15590
rect 15008 -15590 15208 -15552
rect 15008 -15607 15091 -15590
rect 14867 -15624 14883 -15607
rect 14817 -15640 14883 -15624
rect 15075 -15624 15091 -15607
rect 15125 -15607 15208 -15590
rect 15266 -15590 15466 -15552
rect 15266 -15607 15349 -15590
rect 15125 -15624 15141 -15607
rect 15075 -15640 15141 -15624
rect 15333 -15624 15349 -15607
rect 15383 -15607 15466 -15590
rect 15524 -15590 15724 -15552
rect 15524 -15607 15607 -15590
rect 15383 -15624 15399 -15607
rect 15333 -15640 15399 -15624
rect 15591 -15624 15607 -15607
rect 15641 -15607 15724 -15590
rect 15782 -15590 15982 -15552
rect 15782 -15607 15865 -15590
rect 15641 -15624 15657 -15607
rect 15591 -15640 15657 -15624
rect 15849 -15624 15865 -15607
rect 15899 -15607 15982 -15590
rect 16040 -15590 16240 -15552
rect 16040 -15607 16123 -15590
rect 15899 -15624 15915 -15607
rect 15849 -15640 15915 -15624
rect 16107 -15624 16123 -15607
rect 16157 -15607 16240 -15590
rect 16298 -15590 16498 -15552
rect 16298 -15607 16381 -15590
rect 16157 -15624 16173 -15607
rect 16107 -15640 16173 -15624
rect 16365 -15624 16381 -15607
rect 16415 -15607 16498 -15590
rect 16415 -15624 16431 -15607
rect 16365 -15640 16431 -15624
rect 9226 -15699 9292 -15683
rect 9226 -15716 9242 -15699
rect 9159 -15733 9242 -15716
rect 9276 -15716 9292 -15699
rect 9484 -15699 9550 -15683
rect 9484 -15716 9500 -15699
rect 9276 -15733 9359 -15716
rect 9159 -15771 9359 -15733
rect 9417 -15733 9500 -15716
rect 9534 -15716 9550 -15699
rect 9742 -15699 9808 -15683
rect 9742 -15716 9758 -15699
rect 9534 -15733 9617 -15716
rect 9417 -15771 9617 -15733
rect 9675 -15733 9758 -15716
rect 9792 -15716 9808 -15699
rect 10000 -15699 10066 -15683
rect 10000 -15716 10016 -15699
rect 9792 -15733 9875 -15716
rect 9675 -15771 9875 -15733
rect 9933 -15733 10016 -15716
rect 10050 -15716 10066 -15699
rect 10258 -15699 10324 -15683
rect 10258 -15716 10274 -15699
rect 10050 -15733 10133 -15716
rect 9933 -15771 10133 -15733
rect 10191 -15733 10274 -15716
rect 10308 -15716 10324 -15699
rect 10516 -15699 10582 -15683
rect 10516 -15716 10532 -15699
rect 10308 -15733 10391 -15716
rect 10191 -15771 10391 -15733
rect 10449 -15733 10532 -15716
rect 10566 -15716 10582 -15699
rect 10774 -15699 10840 -15683
rect 10774 -15716 10790 -15699
rect 10566 -15733 10649 -15716
rect 10449 -15771 10649 -15733
rect 10707 -15733 10790 -15716
rect 10824 -15716 10840 -15699
rect 11032 -15699 11098 -15683
rect 11032 -15716 11048 -15699
rect 10824 -15733 10907 -15716
rect 10707 -15771 10907 -15733
rect 10965 -15733 11048 -15716
rect 11082 -15716 11098 -15699
rect 11896 -15699 11962 -15683
rect 11896 -15716 11912 -15699
rect 11082 -15733 11165 -15716
rect 10965 -15771 11165 -15733
rect 11829 -15733 11912 -15716
rect 11946 -15716 11962 -15699
rect 12154 -15699 12220 -15683
rect 12154 -15716 12170 -15699
rect 11946 -15733 12029 -15716
rect 11829 -15771 12029 -15733
rect 12087 -15733 12170 -15716
rect 12204 -15716 12220 -15699
rect 12412 -15699 12478 -15683
rect 12412 -15716 12428 -15699
rect 12204 -15733 12287 -15716
rect 12087 -15771 12287 -15733
rect 12345 -15733 12428 -15716
rect 12462 -15716 12478 -15699
rect 12670 -15699 12736 -15683
rect 12670 -15716 12686 -15699
rect 12462 -15733 12545 -15716
rect 12345 -15771 12545 -15733
rect 12603 -15733 12686 -15716
rect 12720 -15716 12736 -15699
rect 12928 -15699 12994 -15683
rect 12928 -15716 12944 -15699
rect 12720 -15733 12803 -15716
rect 12603 -15771 12803 -15733
rect 12861 -15733 12944 -15716
rect 12978 -15716 12994 -15699
rect 13186 -15699 13252 -15683
rect 13186 -15716 13202 -15699
rect 12978 -15733 13061 -15716
rect 12861 -15771 13061 -15733
rect 13119 -15733 13202 -15716
rect 13236 -15716 13252 -15699
rect 13444 -15699 13510 -15683
rect 13444 -15716 13460 -15699
rect 13236 -15733 13319 -15716
rect 13119 -15771 13319 -15733
rect 13377 -15733 13460 -15716
rect 13494 -15716 13510 -15699
rect 13702 -15699 13768 -15683
rect 13702 -15716 13718 -15699
rect 13494 -15733 13577 -15716
rect 13377 -15771 13577 -15733
rect 13635 -15733 13718 -15716
rect 13752 -15716 13768 -15699
rect 14559 -15698 14625 -15682
rect 14559 -15715 14575 -15698
rect 13752 -15733 13835 -15716
rect 13635 -15771 13835 -15733
rect 14492 -15732 14575 -15715
rect 14609 -15715 14625 -15698
rect 14817 -15698 14883 -15682
rect 14817 -15715 14833 -15698
rect 14609 -15732 14692 -15715
rect 14492 -15770 14692 -15732
rect 14750 -15732 14833 -15715
rect 14867 -15715 14883 -15698
rect 15075 -15698 15141 -15682
rect 15075 -15715 15091 -15698
rect 14867 -15732 14950 -15715
rect 14750 -15770 14950 -15732
rect 15008 -15732 15091 -15715
rect 15125 -15715 15141 -15698
rect 15333 -15698 15399 -15682
rect 15333 -15715 15349 -15698
rect 15125 -15732 15208 -15715
rect 15008 -15770 15208 -15732
rect 15266 -15732 15349 -15715
rect 15383 -15715 15399 -15698
rect 15591 -15698 15657 -15682
rect 15591 -15715 15607 -15698
rect 15383 -15732 15466 -15715
rect 15266 -15770 15466 -15732
rect 15524 -15732 15607 -15715
rect 15641 -15715 15657 -15698
rect 15849 -15698 15915 -15682
rect 15849 -15715 15865 -15698
rect 15641 -15732 15724 -15715
rect 15524 -15770 15724 -15732
rect 15782 -15732 15865 -15715
rect 15899 -15715 15915 -15698
rect 16107 -15698 16173 -15682
rect 16107 -15715 16123 -15698
rect 15899 -15732 15982 -15715
rect 15782 -15770 15982 -15732
rect 16040 -15732 16123 -15715
rect 16157 -15715 16173 -15698
rect 16365 -15698 16431 -15682
rect 16365 -15715 16381 -15698
rect 16157 -15732 16240 -15715
rect 16040 -15770 16240 -15732
rect 16298 -15732 16381 -15715
rect 16415 -15715 16431 -15698
rect 16415 -15732 16498 -15715
rect 16298 -15770 16498 -15732
rect 9159 -16009 9359 -15971
rect 9159 -16026 9242 -16009
rect 9226 -16043 9242 -16026
rect 9276 -16026 9359 -16009
rect 9417 -16009 9617 -15971
rect 9417 -16026 9500 -16009
rect 9276 -16043 9292 -16026
rect 9226 -16059 9292 -16043
rect 9484 -16043 9500 -16026
rect 9534 -16026 9617 -16009
rect 9675 -16009 9875 -15971
rect 9675 -16026 9758 -16009
rect 9534 -16043 9550 -16026
rect 9484 -16059 9550 -16043
rect 9742 -16043 9758 -16026
rect 9792 -16026 9875 -16009
rect 9933 -16009 10133 -15971
rect 9933 -16026 10016 -16009
rect 9792 -16043 9808 -16026
rect 9742 -16059 9808 -16043
rect 10000 -16043 10016 -16026
rect 10050 -16026 10133 -16009
rect 10191 -16009 10391 -15971
rect 10191 -16026 10274 -16009
rect 10050 -16043 10066 -16026
rect 10000 -16059 10066 -16043
rect 10258 -16043 10274 -16026
rect 10308 -16026 10391 -16009
rect 10449 -16009 10649 -15971
rect 10449 -16026 10532 -16009
rect 10308 -16043 10324 -16026
rect 10258 -16059 10324 -16043
rect 10516 -16043 10532 -16026
rect 10566 -16026 10649 -16009
rect 10707 -16009 10907 -15971
rect 10707 -16026 10790 -16009
rect 10566 -16043 10582 -16026
rect 10516 -16059 10582 -16043
rect 10774 -16043 10790 -16026
rect 10824 -16026 10907 -16009
rect 10965 -16009 11165 -15971
rect 10965 -16026 11048 -16009
rect 10824 -16043 10840 -16026
rect 10774 -16059 10840 -16043
rect 11032 -16043 11048 -16026
rect 11082 -16026 11165 -16009
rect 11829 -16009 12029 -15971
rect 11829 -16026 11912 -16009
rect 11082 -16043 11098 -16026
rect 11032 -16059 11098 -16043
rect 11896 -16043 11912 -16026
rect 11946 -16026 12029 -16009
rect 12087 -16009 12287 -15971
rect 12087 -16026 12170 -16009
rect 11946 -16043 11962 -16026
rect 11896 -16059 11962 -16043
rect 12154 -16043 12170 -16026
rect 12204 -16026 12287 -16009
rect 12345 -16009 12545 -15971
rect 12345 -16026 12428 -16009
rect 12204 -16043 12220 -16026
rect 12154 -16059 12220 -16043
rect 12412 -16043 12428 -16026
rect 12462 -16026 12545 -16009
rect 12603 -16009 12803 -15971
rect 12603 -16026 12686 -16009
rect 12462 -16043 12478 -16026
rect 12412 -16059 12478 -16043
rect 12670 -16043 12686 -16026
rect 12720 -16026 12803 -16009
rect 12861 -16009 13061 -15971
rect 12861 -16026 12944 -16009
rect 12720 -16043 12736 -16026
rect 12670 -16059 12736 -16043
rect 12928 -16043 12944 -16026
rect 12978 -16026 13061 -16009
rect 13119 -16009 13319 -15971
rect 13119 -16026 13202 -16009
rect 12978 -16043 12994 -16026
rect 12928 -16059 12994 -16043
rect 13186 -16043 13202 -16026
rect 13236 -16026 13319 -16009
rect 13377 -16009 13577 -15971
rect 13377 -16026 13460 -16009
rect 13236 -16043 13252 -16026
rect 13186 -16059 13252 -16043
rect 13444 -16043 13460 -16026
rect 13494 -16026 13577 -16009
rect 13635 -16009 13835 -15971
rect 13635 -16026 13718 -16009
rect 13494 -16043 13510 -16026
rect 13444 -16059 13510 -16043
rect 13702 -16043 13718 -16026
rect 13752 -16026 13835 -16009
rect 14492 -16008 14692 -15970
rect 14492 -16025 14575 -16008
rect 13752 -16043 13768 -16026
rect 13702 -16059 13768 -16043
rect 14559 -16042 14575 -16025
rect 14609 -16025 14692 -16008
rect 14750 -16008 14950 -15970
rect 14750 -16025 14833 -16008
rect 14609 -16042 14625 -16025
rect 14559 -16058 14625 -16042
rect 14817 -16042 14833 -16025
rect 14867 -16025 14950 -16008
rect 15008 -16008 15208 -15970
rect 15008 -16025 15091 -16008
rect 14867 -16042 14883 -16025
rect 14817 -16058 14883 -16042
rect 15075 -16042 15091 -16025
rect 15125 -16025 15208 -16008
rect 15266 -16008 15466 -15970
rect 15266 -16025 15349 -16008
rect 15125 -16042 15141 -16025
rect 15075 -16058 15141 -16042
rect 15333 -16042 15349 -16025
rect 15383 -16025 15466 -16008
rect 15524 -16008 15724 -15970
rect 15524 -16025 15607 -16008
rect 15383 -16042 15399 -16025
rect 15333 -16058 15399 -16042
rect 15591 -16042 15607 -16025
rect 15641 -16025 15724 -16008
rect 15782 -16008 15982 -15970
rect 15782 -16025 15865 -16008
rect 15641 -16042 15657 -16025
rect 15591 -16058 15657 -16042
rect 15849 -16042 15865 -16025
rect 15899 -16025 15982 -16008
rect 16040 -16008 16240 -15970
rect 16040 -16025 16123 -16008
rect 15899 -16042 15915 -16025
rect 15849 -16058 15915 -16042
rect 16107 -16042 16123 -16025
rect 16157 -16025 16240 -16008
rect 16298 -16008 16498 -15970
rect 16298 -16025 16381 -16008
rect 16157 -16042 16173 -16025
rect 16107 -16058 16173 -16042
rect 16365 -16042 16381 -16025
rect 16415 -16025 16498 -16008
rect 16415 -16042 16431 -16025
rect 16365 -16058 16431 -16042
rect 9226 -16117 9292 -16101
rect 9226 -16134 9242 -16117
rect 9159 -16151 9242 -16134
rect 9276 -16134 9292 -16117
rect 9484 -16117 9550 -16101
rect 9484 -16134 9500 -16117
rect 9276 -16151 9359 -16134
rect 9159 -16189 9359 -16151
rect 9417 -16151 9500 -16134
rect 9534 -16134 9550 -16117
rect 9742 -16117 9808 -16101
rect 9742 -16134 9758 -16117
rect 9534 -16151 9617 -16134
rect 9417 -16189 9617 -16151
rect 9675 -16151 9758 -16134
rect 9792 -16134 9808 -16117
rect 10000 -16117 10066 -16101
rect 10000 -16134 10016 -16117
rect 9792 -16151 9875 -16134
rect 9675 -16189 9875 -16151
rect 9933 -16151 10016 -16134
rect 10050 -16134 10066 -16117
rect 10258 -16117 10324 -16101
rect 10258 -16134 10274 -16117
rect 10050 -16151 10133 -16134
rect 9933 -16189 10133 -16151
rect 10191 -16151 10274 -16134
rect 10308 -16134 10324 -16117
rect 10516 -16117 10582 -16101
rect 10516 -16134 10532 -16117
rect 10308 -16151 10391 -16134
rect 10191 -16189 10391 -16151
rect 10449 -16151 10532 -16134
rect 10566 -16134 10582 -16117
rect 10774 -16117 10840 -16101
rect 10774 -16134 10790 -16117
rect 10566 -16151 10649 -16134
rect 10449 -16189 10649 -16151
rect 10707 -16151 10790 -16134
rect 10824 -16134 10840 -16117
rect 11032 -16117 11098 -16101
rect 11032 -16134 11048 -16117
rect 10824 -16151 10907 -16134
rect 10707 -16189 10907 -16151
rect 10965 -16151 11048 -16134
rect 11082 -16134 11098 -16117
rect 11896 -16117 11962 -16101
rect 11896 -16134 11912 -16117
rect 11082 -16151 11165 -16134
rect 10965 -16189 11165 -16151
rect 11829 -16151 11912 -16134
rect 11946 -16134 11962 -16117
rect 12154 -16117 12220 -16101
rect 12154 -16134 12170 -16117
rect 11946 -16151 12029 -16134
rect 11829 -16189 12029 -16151
rect 12087 -16151 12170 -16134
rect 12204 -16134 12220 -16117
rect 12412 -16117 12478 -16101
rect 12412 -16134 12428 -16117
rect 12204 -16151 12287 -16134
rect 12087 -16189 12287 -16151
rect 12345 -16151 12428 -16134
rect 12462 -16134 12478 -16117
rect 12670 -16117 12736 -16101
rect 12670 -16134 12686 -16117
rect 12462 -16151 12545 -16134
rect 12345 -16189 12545 -16151
rect 12603 -16151 12686 -16134
rect 12720 -16134 12736 -16117
rect 12928 -16117 12994 -16101
rect 12928 -16134 12944 -16117
rect 12720 -16151 12803 -16134
rect 12603 -16189 12803 -16151
rect 12861 -16151 12944 -16134
rect 12978 -16134 12994 -16117
rect 13186 -16117 13252 -16101
rect 13186 -16134 13202 -16117
rect 12978 -16151 13061 -16134
rect 12861 -16189 13061 -16151
rect 13119 -16151 13202 -16134
rect 13236 -16134 13252 -16117
rect 13444 -16117 13510 -16101
rect 13444 -16134 13460 -16117
rect 13236 -16151 13319 -16134
rect 13119 -16189 13319 -16151
rect 13377 -16151 13460 -16134
rect 13494 -16134 13510 -16117
rect 13702 -16117 13768 -16101
rect 13702 -16134 13718 -16117
rect 13494 -16151 13577 -16134
rect 13377 -16189 13577 -16151
rect 13635 -16151 13718 -16134
rect 13752 -16134 13768 -16117
rect 14559 -16116 14625 -16100
rect 14559 -16133 14575 -16116
rect 13752 -16151 13835 -16134
rect 13635 -16189 13835 -16151
rect 14492 -16150 14575 -16133
rect 14609 -16133 14625 -16116
rect 14817 -16116 14883 -16100
rect 14817 -16133 14833 -16116
rect 14609 -16150 14692 -16133
rect 14492 -16188 14692 -16150
rect 14750 -16150 14833 -16133
rect 14867 -16133 14883 -16116
rect 15075 -16116 15141 -16100
rect 15075 -16133 15091 -16116
rect 14867 -16150 14950 -16133
rect 14750 -16188 14950 -16150
rect 15008 -16150 15091 -16133
rect 15125 -16133 15141 -16116
rect 15333 -16116 15399 -16100
rect 15333 -16133 15349 -16116
rect 15125 -16150 15208 -16133
rect 15008 -16188 15208 -16150
rect 15266 -16150 15349 -16133
rect 15383 -16133 15399 -16116
rect 15591 -16116 15657 -16100
rect 15591 -16133 15607 -16116
rect 15383 -16150 15466 -16133
rect 15266 -16188 15466 -16150
rect 15524 -16150 15607 -16133
rect 15641 -16133 15657 -16116
rect 15849 -16116 15915 -16100
rect 15849 -16133 15865 -16116
rect 15641 -16150 15724 -16133
rect 15524 -16188 15724 -16150
rect 15782 -16150 15865 -16133
rect 15899 -16133 15915 -16116
rect 16107 -16116 16173 -16100
rect 16107 -16133 16123 -16116
rect 15899 -16150 15982 -16133
rect 15782 -16188 15982 -16150
rect 16040 -16150 16123 -16133
rect 16157 -16133 16173 -16116
rect 16365 -16116 16431 -16100
rect 16365 -16133 16381 -16116
rect 16157 -16150 16240 -16133
rect 16040 -16188 16240 -16150
rect 16298 -16150 16381 -16133
rect 16415 -16133 16431 -16116
rect 16415 -16150 16498 -16133
rect 16298 -16188 16498 -16150
rect 9159 -16427 9359 -16389
rect 9159 -16444 9242 -16427
rect 9226 -16461 9242 -16444
rect 9276 -16444 9359 -16427
rect 9417 -16427 9617 -16389
rect 9417 -16444 9500 -16427
rect 9276 -16461 9292 -16444
rect 9226 -16477 9292 -16461
rect 9484 -16461 9500 -16444
rect 9534 -16444 9617 -16427
rect 9675 -16427 9875 -16389
rect 9675 -16444 9758 -16427
rect 9534 -16461 9550 -16444
rect 9484 -16477 9550 -16461
rect 9742 -16461 9758 -16444
rect 9792 -16444 9875 -16427
rect 9933 -16427 10133 -16389
rect 9933 -16444 10016 -16427
rect 9792 -16461 9808 -16444
rect 9742 -16477 9808 -16461
rect 10000 -16461 10016 -16444
rect 10050 -16444 10133 -16427
rect 10191 -16427 10391 -16389
rect 10191 -16444 10274 -16427
rect 10050 -16461 10066 -16444
rect 10000 -16477 10066 -16461
rect 10258 -16461 10274 -16444
rect 10308 -16444 10391 -16427
rect 10449 -16427 10649 -16389
rect 10449 -16444 10532 -16427
rect 10308 -16461 10324 -16444
rect 10258 -16477 10324 -16461
rect 10516 -16461 10532 -16444
rect 10566 -16444 10649 -16427
rect 10707 -16427 10907 -16389
rect 10707 -16444 10790 -16427
rect 10566 -16461 10582 -16444
rect 10516 -16477 10582 -16461
rect 10774 -16461 10790 -16444
rect 10824 -16444 10907 -16427
rect 10965 -16427 11165 -16389
rect 10965 -16444 11048 -16427
rect 10824 -16461 10840 -16444
rect 10774 -16477 10840 -16461
rect 11032 -16461 11048 -16444
rect 11082 -16444 11165 -16427
rect 11829 -16427 12029 -16389
rect 11829 -16444 11912 -16427
rect 11082 -16461 11098 -16444
rect 11032 -16477 11098 -16461
rect 11896 -16461 11912 -16444
rect 11946 -16444 12029 -16427
rect 12087 -16427 12287 -16389
rect 12087 -16444 12170 -16427
rect 11946 -16461 11962 -16444
rect 11896 -16477 11962 -16461
rect 12154 -16461 12170 -16444
rect 12204 -16444 12287 -16427
rect 12345 -16427 12545 -16389
rect 12345 -16444 12428 -16427
rect 12204 -16461 12220 -16444
rect 12154 -16477 12220 -16461
rect 12412 -16461 12428 -16444
rect 12462 -16444 12545 -16427
rect 12603 -16427 12803 -16389
rect 12603 -16444 12686 -16427
rect 12462 -16461 12478 -16444
rect 12412 -16477 12478 -16461
rect 12670 -16461 12686 -16444
rect 12720 -16444 12803 -16427
rect 12861 -16427 13061 -16389
rect 12861 -16444 12944 -16427
rect 12720 -16461 12736 -16444
rect 12670 -16477 12736 -16461
rect 12928 -16461 12944 -16444
rect 12978 -16444 13061 -16427
rect 13119 -16427 13319 -16389
rect 13119 -16444 13202 -16427
rect 12978 -16461 12994 -16444
rect 12928 -16477 12994 -16461
rect 13186 -16461 13202 -16444
rect 13236 -16444 13319 -16427
rect 13377 -16427 13577 -16389
rect 13377 -16444 13460 -16427
rect 13236 -16461 13252 -16444
rect 13186 -16477 13252 -16461
rect 13444 -16461 13460 -16444
rect 13494 -16444 13577 -16427
rect 13635 -16427 13835 -16389
rect 13635 -16444 13718 -16427
rect 13494 -16461 13510 -16444
rect 13444 -16477 13510 -16461
rect 13702 -16461 13718 -16444
rect 13752 -16444 13835 -16427
rect 14492 -16426 14692 -16388
rect 14492 -16443 14575 -16426
rect 13752 -16461 13768 -16444
rect 13702 -16477 13768 -16461
rect 14559 -16460 14575 -16443
rect 14609 -16443 14692 -16426
rect 14750 -16426 14950 -16388
rect 14750 -16443 14833 -16426
rect 14609 -16460 14625 -16443
rect 14559 -16476 14625 -16460
rect 14817 -16460 14833 -16443
rect 14867 -16443 14950 -16426
rect 15008 -16426 15208 -16388
rect 15008 -16443 15091 -16426
rect 14867 -16460 14883 -16443
rect 14817 -16476 14883 -16460
rect 15075 -16460 15091 -16443
rect 15125 -16443 15208 -16426
rect 15266 -16426 15466 -16388
rect 15266 -16443 15349 -16426
rect 15125 -16460 15141 -16443
rect 15075 -16476 15141 -16460
rect 15333 -16460 15349 -16443
rect 15383 -16443 15466 -16426
rect 15524 -16426 15724 -16388
rect 15524 -16443 15607 -16426
rect 15383 -16460 15399 -16443
rect 15333 -16476 15399 -16460
rect 15591 -16460 15607 -16443
rect 15641 -16443 15724 -16426
rect 15782 -16426 15982 -16388
rect 15782 -16443 15865 -16426
rect 15641 -16460 15657 -16443
rect 15591 -16476 15657 -16460
rect 15849 -16460 15865 -16443
rect 15899 -16443 15982 -16426
rect 16040 -16426 16240 -16388
rect 16040 -16443 16123 -16426
rect 15899 -16460 15915 -16443
rect 15849 -16476 15915 -16460
rect 16107 -16460 16123 -16443
rect 16157 -16443 16240 -16426
rect 16298 -16426 16498 -16388
rect 16298 -16443 16381 -16426
rect 16157 -16460 16173 -16443
rect 16107 -16476 16173 -16460
rect 16365 -16460 16381 -16443
rect 16415 -16443 16498 -16426
rect 16415 -16460 16431 -16443
rect 16365 -16476 16431 -16460
rect 9226 -16535 9292 -16519
rect 9226 -16552 9242 -16535
rect 9159 -16569 9242 -16552
rect 9276 -16552 9292 -16535
rect 9484 -16535 9550 -16519
rect 9484 -16552 9500 -16535
rect 9276 -16569 9359 -16552
rect 9159 -16607 9359 -16569
rect 9417 -16569 9500 -16552
rect 9534 -16552 9550 -16535
rect 9742 -16535 9808 -16519
rect 9742 -16552 9758 -16535
rect 9534 -16569 9617 -16552
rect 9417 -16607 9617 -16569
rect 9675 -16569 9758 -16552
rect 9792 -16552 9808 -16535
rect 10000 -16535 10066 -16519
rect 10000 -16552 10016 -16535
rect 9792 -16569 9875 -16552
rect 9675 -16607 9875 -16569
rect 9933 -16569 10016 -16552
rect 10050 -16552 10066 -16535
rect 10258 -16535 10324 -16519
rect 10258 -16552 10274 -16535
rect 10050 -16569 10133 -16552
rect 9933 -16607 10133 -16569
rect 10191 -16569 10274 -16552
rect 10308 -16552 10324 -16535
rect 10516 -16535 10582 -16519
rect 10516 -16552 10532 -16535
rect 10308 -16569 10391 -16552
rect 10191 -16607 10391 -16569
rect 10449 -16569 10532 -16552
rect 10566 -16552 10582 -16535
rect 10774 -16535 10840 -16519
rect 10774 -16552 10790 -16535
rect 10566 -16569 10649 -16552
rect 10449 -16607 10649 -16569
rect 10707 -16569 10790 -16552
rect 10824 -16552 10840 -16535
rect 11032 -16535 11098 -16519
rect 11032 -16552 11048 -16535
rect 10824 -16569 10907 -16552
rect 10707 -16607 10907 -16569
rect 10965 -16569 11048 -16552
rect 11082 -16552 11098 -16535
rect 11896 -16535 11962 -16519
rect 11896 -16552 11912 -16535
rect 11082 -16569 11165 -16552
rect 10965 -16607 11165 -16569
rect 11829 -16569 11912 -16552
rect 11946 -16552 11962 -16535
rect 12154 -16535 12220 -16519
rect 12154 -16552 12170 -16535
rect 11946 -16569 12029 -16552
rect 11829 -16607 12029 -16569
rect 12087 -16569 12170 -16552
rect 12204 -16552 12220 -16535
rect 12412 -16535 12478 -16519
rect 12412 -16552 12428 -16535
rect 12204 -16569 12287 -16552
rect 12087 -16607 12287 -16569
rect 12345 -16569 12428 -16552
rect 12462 -16552 12478 -16535
rect 12670 -16535 12736 -16519
rect 12670 -16552 12686 -16535
rect 12462 -16569 12545 -16552
rect 12345 -16607 12545 -16569
rect 12603 -16569 12686 -16552
rect 12720 -16552 12736 -16535
rect 12928 -16535 12994 -16519
rect 12928 -16552 12944 -16535
rect 12720 -16569 12803 -16552
rect 12603 -16607 12803 -16569
rect 12861 -16569 12944 -16552
rect 12978 -16552 12994 -16535
rect 13186 -16535 13252 -16519
rect 13186 -16552 13202 -16535
rect 12978 -16569 13061 -16552
rect 12861 -16607 13061 -16569
rect 13119 -16569 13202 -16552
rect 13236 -16552 13252 -16535
rect 13444 -16535 13510 -16519
rect 13444 -16552 13460 -16535
rect 13236 -16569 13319 -16552
rect 13119 -16607 13319 -16569
rect 13377 -16569 13460 -16552
rect 13494 -16552 13510 -16535
rect 13702 -16535 13768 -16519
rect 13702 -16552 13718 -16535
rect 13494 -16569 13577 -16552
rect 13377 -16607 13577 -16569
rect 13635 -16569 13718 -16552
rect 13752 -16552 13768 -16535
rect 14559 -16534 14625 -16518
rect 14559 -16551 14575 -16534
rect 13752 -16569 13835 -16552
rect 13635 -16607 13835 -16569
rect 14492 -16568 14575 -16551
rect 14609 -16551 14625 -16534
rect 14817 -16534 14883 -16518
rect 14817 -16551 14833 -16534
rect 14609 -16568 14692 -16551
rect 14492 -16606 14692 -16568
rect 14750 -16568 14833 -16551
rect 14867 -16551 14883 -16534
rect 15075 -16534 15141 -16518
rect 15075 -16551 15091 -16534
rect 14867 -16568 14950 -16551
rect 14750 -16606 14950 -16568
rect 15008 -16568 15091 -16551
rect 15125 -16551 15141 -16534
rect 15333 -16534 15399 -16518
rect 15333 -16551 15349 -16534
rect 15125 -16568 15208 -16551
rect 15008 -16606 15208 -16568
rect 15266 -16568 15349 -16551
rect 15383 -16551 15399 -16534
rect 15591 -16534 15657 -16518
rect 15591 -16551 15607 -16534
rect 15383 -16568 15466 -16551
rect 15266 -16606 15466 -16568
rect 15524 -16568 15607 -16551
rect 15641 -16551 15657 -16534
rect 15849 -16534 15915 -16518
rect 15849 -16551 15865 -16534
rect 15641 -16568 15724 -16551
rect 15524 -16606 15724 -16568
rect 15782 -16568 15865 -16551
rect 15899 -16551 15915 -16534
rect 16107 -16534 16173 -16518
rect 16107 -16551 16123 -16534
rect 15899 -16568 15982 -16551
rect 15782 -16606 15982 -16568
rect 16040 -16568 16123 -16551
rect 16157 -16551 16173 -16534
rect 16365 -16534 16431 -16518
rect 16365 -16551 16381 -16534
rect 16157 -16568 16240 -16551
rect 16040 -16606 16240 -16568
rect 16298 -16568 16381 -16551
rect 16415 -16551 16431 -16534
rect 16415 -16568 16498 -16551
rect 16298 -16606 16498 -16568
rect 9159 -16845 9359 -16807
rect 9159 -16862 9242 -16845
rect 9226 -16879 9242 -16862
rect 9276 -16862 9359 -16845
rect 9417 -16845 9617 -16807
rect 9417 -16862 9500 -16845
rect 9276 -16879 9292 -16862
rect 9226 -16895 9292 -16879
rect 9484 -16879 9500 -16862
rect 9534 -16862 9617 -16845
rect 9675 -16845 9875 -16807
rect 9675 -16862 9758 -16845
rect 9534 -16879 9550 -16862
rect 9484 -16895 9550 -16879
rect 9742 -16879 9758 -16862
rect 9792 -16862 9875 -16845
rect 9933 -16845 10133 -16807
rect 9933 -16862 10016 -16845
rect 9792 -16879 9808 -16862
rect 9742 -16895 9808 -16879
rect 10000 -16879 10016 -16862
rect 10050 -16862 10133 -16845
rect 10191 -16845 10391 -16807
rect 10191 -16862 10274 -16845
rect 10050 -16879 10066 -16862
rect 10000 -16895 10066 -16879
rect 10258 -16879 10274 -16862
rect 10308 -16862 10391 -16845
rect 10449 -16845 10649 -16807
rect 10449 -16862 10532 -16845
rect 10308 -16879 10324 -16862
rect 10258 -16895 10324 -16879
rect 10516 -16879 10532 -16862
rect 10566 -16862 10649 -16845
rect 10707 -16845 10907 -16807
rect 10707 -16862 10790 -16845
rect 10566 -16879 10582 -16862
rect 10516 -16895 10582 -16879
rect 10774 -16879 10790 -16862
rect 10824 -16862 10907 -16845
rect 10965 -16845 11165 -16807
rect 10965 -16862 11048 -16845
rect 10824 -16879 10840 -16862
rect 10774 -16895 10840 -16879
rect 11032 -16879 11048 -16862
rect 11082 -16862 11165 -16845
rect 11829 -16845 12029 -16807
rect 11829 -16862 11912 -16845
rect 11082 -16879 11098 -16862
rect 11032 -16895 11098 -16879
rect 11896 -16879 11912 -16862
rect 11946 -16862 12029 -16845
rect 12087 -16845 12287 -16807
rect 12087 -16862 12170 -16845
rect 11946 -16879 11962 -16862
rect 11896 -16895 11962 -16879
rect 12154 -16879 12170 -16862
rect 12204 -16862 12287 -16845
rect 12345 -16845 12545 -16807
rect 12345 -16862 12428 -16845
rect 12204 -16879 12220 -16862
rect 12154 -16895 12220 -16879
rect 12412 -16879 12428 -16862
rect 12462 -16862 12545 -16845
rect 12603 -16845 12803 -16807
rect 12603 -16862 12686 -16845
rect 12462 -16879 12478 -16862
rect 12412 -16895 12478 -16879
rect 12670 -16879 12686 -16862
rect 12720 -16862 12803 -16845
rect 12861 -16845 13061 -16807
rect 12861 -16862 12944 -16845
rect 12720 -16879 12736 -16862
rect 12670 -16895 12736 -16879
rect 12928 -16879 12944 -16862
rect 12978 -16862 13061 -16845
rect 13119 -16845 13319 -16807
rect 13119 -16862 13202 -16845
rect 12978 -16879 12994 -16862
rect 12928 -16895 12994 -16879
rect 13186 -16879 13202 -16862
rect 13236 -16862 13319 -16845
rect 13377 -16845 13577 -16807
rect 13377 -16862 13460 -16845
rect 13236 -16879 13252 -16862
rect 13186 -16895 13252 -16879
rect 13444 -16879 13460 -16862
rect 13494 -16862 13577 -16845
rect 13635 -16845 13835 -16807
rect 13635 -16862 13718 -16845
rect 13494 -16879 13510 -16862
rect 13444 -16895 13510 -16879
rect 13702 -16879 13718 -16862
rect 13752 -16862 13835 -16845
rect 14492 -16844 14692 -16806
rect 14492 -16861 14575 -16844
rect 13752 -16879 13768 -16862
rect 13702 -16895 13768 -16879
rect 14559 -16878 14575 -16861
rect 14609 -16861 14692 -16844
rect 14750 -16844 14950 -16806
rect 14750 -16861 14833 -16844
rect 14609 -16878 14625 -16861
rect 14559 -16894 14625 -16878
rect 14817 -16878 14833 -16861
rect 14867 -16861 14950 -16844
rect 15008 -16844 15208 -16806
rect 15008 -16861 15091 -16844
rect 14867 -16878 14883 -16861
rect 14817 -16894 14883 -16878
rect 15075 -16878 15091 -16861
rect 15125 -16861 15208 -16844
rect 15266 -16844 15466 -16806
rect 15266 -16861 15349 -16844
rect 15125 -16878 15141 -16861
rect 15075 -16894 15141 -16878
rect 15333 -16878 15349 -16861
rect 15383 -16861 15466 -16844
rect 15524 -16844 15724 -16806
rect 15524 -16861 15607 -16844
rect 15383 -16878 15399 -16861
rect 15333 -16894 15399 -16878
rect 15591 -16878 15607 -16861
rect 15641 -16861 15724 -16844
rect 15782 -16844 15982 -16806
rect 15782 -16861 15865 -16844
rect 15641 -16878 15657 -16861
rect 15591 -16894 15657 -16878
rect 15849 -16878 15865 -16861
rect 15899 -16861 15982 -16844
rect 16040 -16844 16240 -16806
rect 16040 -16861 16123 -16844
rect 15899 -16878 15915 -16861
rect 15849 -16894 15915 -16878
rect 16107 -16878 16123 -16861
rect 16157 -16861 16240 -16844
rect 16298 -16844 16498 -16806
rect 16298 -16861 16381 -16844
rect 16157 -16878 16173 -16861
rect 16107 -16894 16173 -16878
rect 16365 -16878 16381 -16861
rect 16415 -16861 16498 -16844
rect 16415 -16878 16431 -16861
rect 16365 -16894 16431 -16878
rect 9226 -16953 9292 -16937
rect 9226 -16970 9242 -16953
rect 9159 -16987 9242 -16970
rect 9276 -16970 9292 -16953
rect 9484 -16953 9550 -16937
rect 9484 -16970 9500 -16953
rect 9276 -16987 9359 -16970
rect 9159 -17025 9359 -16987
rect 9417 -16987 9500 -16970
rect 9534 -16970 9550 -16953
rect 9742 -16953 9808 -16937
rect 9742 -16970 9758 -16953
rect 9534 -16987 9617 -16970
rect 9417 -17025 9617 -16987
rect 9675 -16987 9758 -16970
rect 9792 -16970 9808 -16953
rect 10000 -16953 10066 -16937
rect 10000 -16970 10016 -16953
rect 9792 -16987 9875 -16970
rect 9675 -17025 9875 -16987
rect 9933 -16987 10016 -16970
rect 10050 -16970 10066 -16953
rect 10258 -16953 10324 -16937
rect 10258 -16970 10274 -16953
rect 10050 -16987 10133 -16970
rect 9933 -17025 10133 -16987
rect 10191 -16987 10274 -16970
rect 10308 -16970 10324 -16953
rect 10516 -16953 10582 -16937
rect 10516 -16970 10532 -16953
rect 10308 -16987 10391 -16970
rect 10191 -17025 10391 -16987
rect 10449 -16987 10532 -16970
rect 10566 -16970 10582 -16953
rect 10774 -16953 10840 -16937
rect 10774 -16970 10790 -16953
rect 10566 -16987 10649 -16970
rect 10449 -17025 10649 -16987
rect 10707 -16987 10790 -16970
rect 10824 -16970 10840 -16953
rect 11032 -16953 11098 -16937
rect 11032 -16970 11048 -16953
rect 10824 -16987 10907 -16970
rect 10707 -17025 10907 -16987
rect 10965 -16987 11048 -16970
rect 11082 -16970 11098 -16953
rect 11896 -16953 11962 -16937
rect 11896 -16970 11912 -16953
rect 11082 -16987 11165 -16970
rect 10965 -17025 11165 -16987
rect 11829 -16987 11912 -16970
rect 11946 -16970 11962 -16953
rect 12154 -16953 12220 -16937
rect 12154 -16970 12170 -16953
rect 11946 -16987 12029 -16970
rect 11829 -17025 12029 -16987
rect 12087 -16987 12170 -16970
rect 12204 -16970 12220 -16953
rect 12412 -16953 12478 -16937
rect 12412 -16970 12428 -16953
rect 12204 -16987 12287 -16970
rect 12087 -17025 12287 -16987
rect 12345 -16987 12428 -16970
rect 12462 -16970 12478 -16953
rect 12670 -16953 12736 -16937
rect 12670 -16970 12686 -16953
rect 12462 -16987 12545 -16970
rect 12345 -17025 12545 -16987
rect 12603 -16987 12686 -16970
rect 12720 -16970 12736 -16953
rect 12928 -16953 12994 -16937
rect 12928 -16970 12944 -16953
rect 12720 -16987 12803 -16970
rect 12603 -17025 12803 -16987
rect 12861 -16987 12944 -16970
rect 12978 -16970 12994 -16953
rect 13186 -16953 13252 -16937
rect 13186 -16970 13202 -16953
rect 12978 -16987 13061 -16970
rect 12861 -17025 13061 -16987
rect 13119 -16987 13202 -16970
rect 13236 -16970 13252 -16953
rect 13444 -16953 13510 -16937
rect 13444 -16970 13460 -16953
rect 13236 -16987 13319 -16970
rect 13119 -17025 13319 -16987
rect 13377 -16987 13460 -16970
rect 13494 -16970 13510 -16953
rect 13702 -16953 13768 -16937
rect 13702 -16970 13718 -16953
rect 13494 -16987 13577 -16970
rect 13377 -17025 13577 -16987
rect 13635 -16987 13718 -16970
rect 13752 -16970 13768 -16953
rect 14559 -16952 14625 -16936
rect 14559 -16969 14575 -16952
rect 13752 -16987 13835 -16970
rect 13635 -17025 13835 -16987
rect 14492 -16986 14575 -16969
rect 14609 -16969 14625 -16952
rect 14817 -16952 14883 -16936
rect 14817 -16969 14833 -16952
rect 14609 -16986 14692 -16969
rect 14492 -17024 14692 -16986
rect 14750 -16986 14833 -16969
rect 14867 -16969 14883 -16952
rect 15075 -16952 15141 -16936
rect 15075 -16969 15091 -16952
rect 14867 -16986 14950 -16969
rect 14750 -17024 14950 -16986
rect 15008 -16986 15091 -16969
rect 15125 -16969 15141 -16952
rect 15333 -16952 15399 -16936
rect 15333 -16969 15349 -16952
rect 15125 -16986 15208 -16969
rect 15008 -17024 15208 -16986
rect 15266 -16986 15349 -16969
rect 15383 -16969 15399 -16952
rect 15591 -16952 15657 -16936
rect 15591 -16969 15607 -16952
rect 15383 -16986 15466 -16969
rect 15266 -17024 15466 -16986
rect 15524 -16986 15607 -16969
rect 15641 -16969 15657 -16952
rect 15849 -16952 15915 -16936
rect 15849 -16969 15865 -16952
rect 15641 -16986 15724 -16969
rect 15524 -17024 15724 -16986
rect 15782 -16986 15865 -16969
rect 15899 -16969 15915 -16952
rect 16107 -16952 16173 -16936
rect 16107 -16969 16123 -16952
rect 15899 -16986 15982 -16969
rect 15782 -17024 15982 -16986
rect 16040 -16986 16123 -16969
rect 16157 -16969 16173 -16952
rect 16365 -16952 16431 -16936
rect 16365 -16969 16381 -16952
rect 16157 -16986 16240 -16969
rect 16040 -17024 16240 -16986
rect 16298 -16986 16381 -16969
rect 16415 -16969 16431 -16952
rect 16415 -16986 16498 -16969
rect 16298 -17024 16498 -16986
rect 9159 -17263 9359 -17225
rect 9159 -17280 9242 -17263
rect 9226 -17297 9242 -17280
rect 9276 -17280 9359 -17263
rect 9417 -17263 9617 -17225
rect 9417 -17280 9500 -17263
rect 9276 -17297 9292 -17280
rect 9226 -17313 9292 -17297
rect 9484 -17297 9500 -17280
rect 9534 -17280 9617 -17263
rect 9675 -17263 9875 -17225
rect 9675 -17280 9758 -17263
rect 9534 -17297 9550 -17280
rect 9484 -17313 9550 -17297
rect 9742 -17297 9758 -17280
rect 9792 -17280 9875 -17263
rect 9933 -17263 10133 -17225
rect 9933 -17280 10016 -17263
rect 9792 -17297 9808 -17280
rect 9742 -17313 9808 -17297
rect 10000 -17297 10016 -17280
rect 10050 -17280 10133 -17263
rect 10191 -17263 10391 -17225
rect 10191 -17280 10274 -17263
rect 10050 -17297 10066 -17280
rect 10000 -17313 10066 -17297
rect 10258 -17297 10274 -17280
rect 10308 -17280 10391 -17263
rect 10449 -17263 10649 -17225
rect 10449 -17280 10532 -17263
rect 10308 -17297 10324 -17280
rect 10258 -17313 10324 -17297
rect 10516 -17297 10532 -17280
rect 10566 -17280 10649 -17263
rect 10707 -17263 10907 -17225
rect 10707 -17280 10790 -17263
rect 10566 -17297 10582 -17280
rect 10516 -17313 10582 -17297
rect 10774 -17297 10790 -17280
rect 10824 -17280 10907 -17263
rect 10965 -17263 11165 -17225
rect 10965 -17280 11048 -17263
rect 10824 -17297 10840 -17280
rect 10774 -17313 10840 -17297
rect 11032 -17297 11048 -17280
rect 11082 -17280 11165 -17263
rect 11829 -17263 12029 -17225
rect 11829 -17280 11912 -17263
rect 11082 -17297 11098 -17280
rect 11032 -17313 11098 -17297
rect 11896 -17297 11912 -17280
rect 11946 -17280 12029 -17263
rect 12087 -17263 12287 -17225
rect 12087 -17280 12170 -17263
rect 11946 -17297 11962 -17280
rect 11896 -17313 11962 -17297
rect 12154 -17297 12170 -17280
rect 12204 -17280 12287 -17263
rect 12345 -17263 12545 -17225
rect 12345 -17280 12428 -17263
rect 12204 -17297 12220 -17280
rect 12154 -17313 12220 -17297
rect 12412 -17297 12428 -17280
rect 12462 -17280 12545 -17263
rect 12603 -17263 12803 -17225
rect 12603 -17280 12686 -17263
rect 12462 -17297 12478 -17280
rect 12412 -17313 12478 -17297
rect 12670 -17297 12686 -17280
rect 12720 -17280 12803 -17263
rect 12861 -17263 13061 -17225
rect 12861 -17280 12944 -17263
rect 12720 -17297 12736 -17280
rect 12670 -17313 12736 -17297
rect 12928 -17297 12944 -17280
rect 12978 -17280 13061 -17263
rect 13119 -17263 13319 -17225
rect 13119 -17280 13202 -17263
rect 12978 -17297 12994 -17280
rect 12928 -17313 12994 -17297
rect 13186 -17297 13202 -17280
rect 13236 -17280 13319 -17263
rect 13377 -17263 13577 -17225
rect 13377 -17280 13460 -17263
rect 13236 -17297 13252 -17280
rect 13186 -17313 13252 -17297
rect 13444 -17297 13460 -17280
rect 13494 -17280 13577 -17263
rect 13635 -17263 13835 -17225
rect 13635 -17280 13718 -17263
rect 13494 -17297 13510 -17280
rect 13444 -17313 13510 -17297
rect 13702 -17297 13718 -17280
rect 13752 -17280 13835 -17263
rect 14492 -17262 14692 -17224
rect 14492 -17279 14575 -17262
rect 13752 -17297 13768 -17280
rect 13702 -17313 13768 -17297
rect 14559 -17296 14575 -17279
rect 14609 -17279 14692 -17262
rect 14750 -17262 14950 -17224
rect 14750 -17279 14833 -17262
rect 14609 -17296 14625 -17279
rect 14559 -17312 14625 -17296
rect 14817 -17296 14833 -17279
rect 14867 -17279 14950 -17262
rect 15008 -17262 15208 -17224
rect 15008 -17279 15091 -17262
rect 14867 -17296 14883 -17279
rect 14817 -17312 14883 -17296
rect 15075 -17296 15091 -17279
rect 15125 -17279 15208 -17262
rect 15266 -17262 15466 -17224
rect 15266 -17279 15349 -17262
rect 15125 -17296 15141 -17279
rect 15075 -17312 15141 -17296
rect 15333 -17296 15349 -17279
rect 15383 -17279 15466 -17262
rect 15524 -17262 15724 -17224
rect 15524 -17279 15607 -17262
rect 15383 -17296 15399 -17279
rect 15333 -17312 15399 -17296
rect 15591 -17296 15607 -17279
rect 15641 -17279 15724 -17262
rect 15782 -17262 15982 -17224
rect 15782 -17279 15865 -17262
rect 15641 -17296 15657 -17279
rect 15591 -17312 15657 -17296
rect 15849 -17296 15865 -17279
rect 15899 -17279 15982 -17262
rect 16040 -17262 16240 -17224
rect 16040 -17279 16123 -17262
rect 15899 -17296 15915 -17279
rect 15849 -17312 15915 -17296
rect 16107 -17296 16123 -17279
rect 16157 -17279 16240 -17262
rect 16298 -17262 16498 -17224
rect 16298 -17279 16381 -17262
rect 16157 -17296 16173 -17279
rect 16107 -17312 16173 -17296
rect 16365 -17296 16381 -17279
rect 16415 -17279 16498 -17262
rect 16415 -17296 16431 -17279
rect 16365 -17312 16431 -17296
rect 9226 -17371 9292 -17355
rect 9226 -17388 9242 -17371
rect 9159 -17405 9242 -17388
rect 9276 -17388 9292 -17371
rect 9484 -17371 9550 -17355
rect 9484 -17388 9500 -17371
rect 9276 -17405 9359 -17388
rect 9159 -17443 9359 -17405
rect 9417 -17405 9500 -17388
rect 9534 -17388 9550 -17371
rect 9742 -17371 9808 -17355
rect 9742 -17388 9758 -17371
rect 9534 -17405 9617 -17388
rect 9417 -17443 9617 -17405
rect 9675 -17405 9758 -17388
rect 9792 -17388 9808 -17371
rect 10000 -17371 10066 -17355
rect 10000 -17388 10016 -17371
rect 9792 -17405 9875 -17388
rect 9675 -17443 9875 -17405
rect 9933 -17405 10016 -17388
rect 10050 -17388 10066 -17371
rect 10258 -17371 10324 -17355
rect 10258 -17388 10274 -17371
rect 10050 -17405 10133 -17388
rect 9933 -17443 10133 -17405
rect 10191 -17405 10274 -17388
rect 10308 -17388 10324 -17371
rect 10516 -17371 10582 -17355
rect 10516 -17388 10532 -17371
rect 10308 -17405 10391 -17388
rect 10191 -17443 10391 -17405
rect 10449 -17405 10532 -17388
rect 10566 -17388 10582 -17371
rect 10774 -17371 10840 -17355
rect 10774 -17388 10790 -17371
rect 10566 -17405 10649 -17388
rect 10449 -17443 10649 -17405
rect 10707 -17405 10790 -17388
rect 10824 -17388 10840 -17371
rect 11032 -17371 11098 -17355
rect 11032 -17388 11048 -17371
rect 10824 -17405 10907 -17388
rect 10707 -17443 10907 -17405
rect 10965 -17405 11048 -17388
rect 11082 -17388 11098 -17371
rect 11896 -17371 11962 -17355
rect 11896 -17388 11912 -17371
rect 11082 -17405 11165 -17388
rect 10965 -17443 11165 -17405
rect 11829 -17405 11912 -17388
rect 11946 -17388 11962 -17371
rect 12154 -17371 12220 -17355
rect 12154 -17388 12170 -17371
rect 11946 -17405 12029 -17388
rect 11829 -17443 12029 -17405
rect 12087 -17405 12170 -17388
rect 12204 -17388 12220 -17371
rect 12412 -17371 12478 -17355
rect 12412 -17388 12428 -17371
rect 12204 -17405 12287 -17388
rect 12087 -17443 12287 -17405
rect 12345 -17405 12428 -17388
rect 12462 -17388 12478 -17371
rect 12670 -17371 12736 -17355
rect 12670 -17388 12686 -17371
rect 12462 -17405 12545 -17388
rect 12345 -17443 12545 -17405
rect 12603 -17405 12686 -17388
rect 12720 -17388 12736 -17371
rect 12928 -17371 12994 -17355
rect 12928 -17388 12944 -17371
rect 12720 -17405 12803 -17388
rect 12603 -17443 12803 -17405
rect 12861 -17405 12944 -17388
rect 12978 -17388 12994 -17371
rect 13186 -17371 13252 -17355
rect 13186 -17388 13202 -17371
rect 12978 -17405 13061 -17388
rect 12861 -17443 13061 -17405
rect 13119 -17405 13202 -17388
rect 13236 -17388 13252 -17371
rect 13444 -17371 13510 -17355
rect 13444 -17388 13460 -17371
rect 13236 -17405 13319 -17388
rect 13119 -17443 13319 -17405
rect 13377 -17405 13460 -17388
rect 13494 -17388 13510 -17371
rect 13702 -17371 13768 -17355
rect 13702 -17388 13718 -17371
rect 13494 -17405 13577 -17388
rect 13377 -17443 13577 -17405
rect 13635 -17405 13718 -17388
rect 13752 -17388 13768 -17371
rect 14559 -17370 14625 -17354
rect 14559 -17387 14575 -17370
rect 13752 -17405 13835 -17388
rect 13635 -17443 13835 -17405
rect 14492 -17404 14575 -17387
rect 14609 -17387 14625 -17370
rect 14817 -17370 14883 -17354
rect 14817 -17387 14833 -17370
rect 14609 -17404 14692 -17387
rect 14492 -17442 14692 -17404
rect 14750 -17404 14833 -17387
rect 14867 -17387 14883 -17370
rect 15075 -17370 15141 -17354
rect 15075 -17387 15091 -17370
rect 14867 -17404 14950 -17387
rect 14750 -17442 14950 -17404
rect 15008 -17404 15091 -17387
rect 15125 -17387 15141 -17370
rect 15333 -17370 15399 -17354
rect 15333 -17387 15349 -17370
rect 15125 -17404 15208 -17387
rect 15008 -17442 15208 -17404
rect 15266 -17404 15349 -17387
rect 15383 -17387 15399 -17370
rect 15591 -17370 15657 -17354
rect 15591 -17387 15607 -17370
rect 15383 -17404 15466 -17387
rect 15266 -17442 15466 -17404
rect 15524 -17404 15607 -17387
rect 15641 -17387 15657 -17370
rect 15849 -17370 15915 -17354
rect 15849 -17387 15865 -17370
rect 15641 -17404 15724 -17387
rect 15524 -17442 15724 -17404
rect 15782 -17404 15865 -17387
rect 15899 -17387 15915 -17370
rect 16107 -17370 16173 -17354
rect 16107 -17387 16123 -17370
rect 15899 -17404 15982 -17387
rect 15782 -17442 15982 -17404
rect 16040 -17404 16123 -17387
rect 16157 -17387 16173 -17370
rect 16365 -17370 16431 -17354
rect 16365 -17387 16381 -17370
rect 16157 -17404 16240 -17387
rect 16040 -17442 16240 -17404
rect 16298 -17404 16381 -17387
rect 16415 -17387 16431 -17370
rect 16415 -17404 16498 -17387
rect 16298 -17442 16498 -17404
rect 9159 -17681 9359 -17643
rect 9159 -17698 9242 -17681
rect 9226 -17715 9242 -17698
rect 9276 -17698 9359 -17681
rect 9417 -17681 9617 -17643
rect 9417 -17698 9500 -17681
rect 9276 -17715 9292 -17698
rect 9226 -17731 9292 -17715
rect 9484 -17715 9500 -17698
rect 9534 -17698 9617 -17681
rect 9675 -17681 9875 -17643
rect 9675 -17698 9758 -17681
rect 9534 -17715 9550 -17698
rect 9484 -17731 9550 -17715
rect 9742 -17715 9758 -17698
rect 9792 -17698 9875 -17681
rect 9933 -17681 10133 -17643
rect 9933 -17698 10016 -17681
rect 9792 -17715 9808 -17698
rect 9742 -17731 9808 -17715
rect 10000 -17715 10016 -17698
rect 10050 -17698 10133 -17681
rect 10191 -17681 10391 -17643
rect 10191 -17698 10274 -17681
rect 10050 -17715 10066 -17698
rect 10000 -17731 10066 -17715
rect 10258 -17715 10274 -17698
rect 10308 -17698 10391 -17681
rect 10449 -17681 10649 -17643
rect 10449 -17698 10532 -17681
rect 10308 -17715 10324 -17698
rect 10258 -17731 10324 -17715
rect 10516 -17715 10532 -17698
rect 10566 -17698 10649 -17681
rect 10707 -17681 10907 -17643
rect 10707 -17698 10790 -17681
rect 10566 -17715 10582 -17698
rect 10516 -17731 10582 -17715
rect 10774 -17715 10790 -17698
rect 10824 -17698 10907 -17681
rect 10965 -17681 11165 -17643
rect 10965 -17698 11048 -17681
rect 10824 -17715 10840 -17698
rect 10774 -17731 10840 -17715
rect 11032 -17715 11048 -17698
rect 11082 -17698 11165 -17681
rect 11829 -17681 12029 -17643
rect 11829 -17698 11912 -17681
rect 11082 -17715 11098 -17698
rect 11032 -17731 11098 -17715
rect 11896 -17715 11912 -17698
rect 11946 -17698 12029 -17681
rect 12087 -17681 12287 -17643
rect 12087 -17698 12170 -17681
rect 11946 -17715 11962 -17698
rect 11896 -17731 11962 -17715
rect 12154 -17715 12170 -17698
rect 12204 -17698 12287 -17681
rect 12345 -17681 12545 -17643
rect 12345 -17698 12428 -17681
rect 12204 -17715 12220 -17698
rect 12154 -17731 12220 -17715
rect 12412 -17715 12428 -17698
rect 12462 -17698 12545 -17681
rect 12603 -17681 12803 -17643
rect 12603 -17698 12686 -17681
rect 12462 -17715 12478 -17698
rect 12412 -17731 12478 -17715
rect 12670 -17715 12686 -17698
rect 12720 -17698 12803 -17681
rect 12861 -17681 13061 -17643
rect 12861 -17698 12944 -17681
rect 12720 -17715 12736 -17698
rect 12670 -17731 12736 -17715
rect 12928 -17715 12944 -17698
rect 12978 -17698 13061 -17681
rect 13119 -17681 13319 -17643
rect 13119 -17698 13202 -17681
rect 12978 -17715 12994 -17698
rect 12928 -17731 12994 -17715
rect 13186 -17715 13202 -17698
rect 13236 -17698 13319 -17681
rect 13377 -17681 13577 -17643
rect 13377 -17698 13460 -17681
rect 13236 -17715 13252 -17698
rect 13186 -17731 13252 -17715
rect 13444 -17715 13460 -17698
rect 13494 -17698 13577 -17681
rect 13635 -17681 13835 -17643
rect 13635 -17698 13718 -17681
rect 13494 -17715 13510 -17698
rect 13444 -17731 13510 -17715
rect 13702 -17715 13718 -17698
rect 13752 -17698 13835 -17681
rect 14492 -17680 14692 -17642
rect 14492 -17697 14575 -17680
rect 13752 -17715 13768 -17698
rect 13702 -17731 13768 -17715
rect 14559 -17714 14575 -17697
rect 14609 -17697 14692 -17680
rect 14750 -17680 14950 -17642
rect 14750 -17697 14833 -17680
rect 14609 -17714 14625 -17697
rect 14559 -17730 14625 -17714
rect 14817 -17714 14833 -17697
rect 14867 -17697 14950 -17680
rect 15008 -17680 15208 -17642
rect 15008 -17697 15091 -17680
rect 14867 -17714 14883 -17697
rect 14817 -17730 14883 -17714
rect 15075 -17714 15091 -17697
rect 15125 -17697 15208 -17680
rect 15266 -17680 15466 -17642
rect 15266 -17697 15349 -17680
rect 15125 -17714 15141 -17697
rect 15075 -17730 15141 -17714
rect 15333 -17714 15349 -17697
rect 15383 -17697 15466 -17680
rect 15524 -17680 15724 -17642
rect 15524 -17697 15607 -17680
rect 15383 -17714 15399 -17697
rect 15333 -17730 15399 -17714
rect 15591 -17714 15607 -17697
rect 15641 -17697 15724 -17680
rect 15782 -17680 15982 -17642
rect 15782 -17697 15865 -17680
rect 15641 -17714 15657 -17697
rect 15591 -17730 15657 -17714
rect 15849 -17714 15865 -17697
rect 15899 -17697 15982 -17680
rect 16040 -17680 16240 -17642
rect 16040 -17697 16123 -17680
rect 15899 -17714 15915 -17697
rect 15849 -17730 15915 -17714
rect 16107 -17714 16123 -17697
rect 16157 -17697 16240 -17680
rect 16298 -17680 16498 -17642
rect 16298 -17697 16381 -17680
rect 16157 -17714 16173 -17697
rect 16107 -17730 16173 -17714
rect 16365 -17714 16381 -17697
rect 16415 -17697 16498 -17680
rect 16415 -17714 16431 -17697
rect 16365 -17730 16431 -17714
rect 9226 -17789 9292 -17773
rect 9226 -17806 9242 -17789
rect 9159 -17823 9242 -17806
rect 9276 -17806 9292 -17789
rect 9484 -17789 9550 -17773
rect 9484 -17806 9500 -17789
rect 9276 -17823 9359 -17806
rect 9159 -17861 9359 -17823
rect 9417 -17823 9500 -17806
rect 9534 -17806 9550 -17789
rect 9742 -17789 9808 -17773
rect 9742 -17806 9758 -17789
rect 9534 -17823 9617 -17806
rect 9417 -17861 9617 -17823
rect 9675 -17823 9758 -17806
rect 9792 -17806 9808 -17789
rect 10000 -17789 10066 -17773
rect 10000 -17806 10016 -17789
rect 9792 -17823 9875 -17806
rect 9675 -17861 9875 -17823
rect 9933 -17823 10016 -17806
rect 10050 -17806 10066 -17789
rect 10258 -17789 10324 -17773
rect 10258 -17806 10274 -17789
rect 10050 -17823 10133 -17806
rect 9933 -17861 10133 -17823
rect 10191 -17823 10274 -17806
rect 10308 -17806 10324 -17789
rect 10516 -17789 10582 -17773
rect 10516 -17806 10532 -17789
rect 10308 -17823 10391 -17806
rect 10191 -17861 10391 -17823
rect 10449 -17823 10532 -17806
rect 10566 -17806 10582 -17789
rect 10774 -17789 10840 -17773
rect 10774 -17806 10790 -17789
rect 10566 -17823 10649 -17806
rect 10449 -17861 10649 -17823
rect 10707 -17823 10790 -17806
rect 10824 -17806 10840 -17789
rect 11032 -17789 11098 -17773
rect 11032 -17806 11048 -17789
rect 10824 -17823 10907 -17806
rect 10707 -17861 10907 -17823
rect 10965 -17823 11048 -17806
rect 11082 -17806 11098 -17789
rect 11896 -17789 11962 -17773
rect 11896 -17806 11912 -17789
rect 11082 -17823 11165 -17806
rect 10965 -17861 11165 -17823
rect 11829 -17823 11912 -17806
rect 11946 -17806 11962 -17789
rect 12154 -17789 12220 -17773
rect 12154 -17806 12170 -17789
rect 11946 -17823 12029 -17806
rect 11829 -17861 12029 -17823
rect 12087 -17823 12170 -17806
rect 12204 -17806 12220 -17789
rect 12412 -17789 12478 -17773
rect 12412 -17806 12428 -17789
rect 12204 -17823 12287 -17806
rect 12087 -17861 12287 -17823
rect 12345 -17823 12428 -17806
rect 12462 -17806 12478 -17789
rect 12670 -17789 12736 -17773
rect 12670 -17806 12686 -17789
rect 12462 -17823 12545 -17806
rect 12345 -17861 12545 -17823
rect 12603 -17823 12686 -17806
rect 12720 -17806 12736 -17789
rect 12928 -17789 12994 -17773
rect 12928 -17806 12944 -17789
rect 12720 -17823 12803 -17806
rect 12603 -17861 12803 -17823
rect 12861 -17823 12944 -17806
rect 12978 -17806 12994 -17789
rect 13186 -17789 13252 -17773
rect 13186 -17806 13202 -17789
rect 12978 -17823 13061 -17806
rect 12861 -17861 13061 -17823
rect 13119 -17823 13202 -17806
rect 13236 -17806 13252 -17789
rect 13444 -17789 13510 -17773
rect 13444 -17806 13460 -17789
rect 13236 -17823 13319 -17806
rect 13119 -17861 13319 -17823
rect 13377 -17823 13460 -17806
rect 13494 -17806 13510 -17789
rect 13702 -17789 13768 -17773
rect 13702 -17806 13718 -17789
rect 13494 -17823 13577 -17806
rect 13377 -17861 13577 -17823
rect 13635 -17823 13718 -17806
rect 13752 -17806 13768 -17789
rect 14559 -17788 14625 -17772
rect 14559 -17805 14575 -17788
rect 13752 -17823 13835 -17806
rect 13635 -17861 13835 -17823
rect 14492 -17822 14575 -17805
rect 14609 -17805 14625 -17788
rect 14817 -17788 14883 -17772
rect 14817 -17805 14833 -17788
rect 14609 -17822 14692 -17805
rect 14492 -17860 14692 -17822
rect 14750 -17822 14833 -17805
rect 14867 -17805 14883 -17788
rect 15075 -17788 15141 -17772
rect 15075 -17805 15091 -17788
rect 14867 -17822 14950 -17805
rect 14750 -17860 14950 -17822
rect 15008 -17822 15091 -17805
rect 15125 -17805 15141 -17788
rect 15333 -17788 15399 -17772
rect 15333 -17805 15349 -17788
rect 15125 -17822 15208 -17805
rect 15008 -17860 15208 -17822
rect 15266 -17822 15349 -17805
rect 15383 -17805 15399 -17788
rect 15591 -17788 15657 -17772
rect 15591 -17805 15607 -17788
rect 15383 -17822 15466 -17805
rect 15266 -17860 15466 -17822
rect 15524 -17822 15607 -17805
rect 15641 -17805 15657 -17788
rect 15849 -17788 15915 -17772
rect 15849 -17805 15865 -17788
rect 15641 -17822 15724 -17805
rect 15524 -17860 15724 -17822
rect 15782 -17822 15865 -17805
rect 15899 -17805 15915 -17788
rect 16107 -17788 16173 -17772
rect 16107 -17805 16123 -17788
rect 15899 -17822 15982 -17805
rect 15782 -17860 15982 -17822
rect 16040 -17822 16123 -17805
rect 16157 -17805 16173 -17788
rect 16365 -17788 16431 -17772
rect 16365 -17805 16381 -17788
rect 16157 -17822 16240 -17805
rect 16040 -17860 16240 -17822
rect 16298 -17822 16381 -17805
rect 16415 -17805 16431 -17788
rect 16415 -17822 16498 -17805
rect 16298 -17860 16498 -17822
rect 9159 -18099 9359 -18061
rect 9159 -18116 9242 -18099
rect 9226 -18133 9242 -18116
rect 9276 -18116 9359 -18099
rect 9417 -18099 9617 -18061
rect 9417 -18116 9500 -18099
rect 9276 -18133 9292 -18116
rect 9226 -18149 9292 -18133
rect 9484 -18133 9500 -18116
rect 9534 -18116 9617 -18099
rect 9675 -18099 9875 -18061
rect 9675 -18116 9758 -18099
rect 9534 -18133 9550 -18116
rect 9484 -18149 9550 -18133
rect 9742 -18133 9758 -18116
rect 9792 -18116 9875 -18099
rect 9933 -18099 10133 -18061
rect 9933 -18116 10016 -18099
rect 9792 -18133 9808 -18116
rect 9742 -18149 9808 -18133
rect 10000 -18133 10016 -18116
rect 10050 -18116 10133 -18099
rect 10191 -18099 10391 -18061
rect 10191 -18116 10274 -18099
rect 10050 -18133 10066 -18116
rect 10000 -18149 10066 -18133
rect 10258 -18133 10274 -18116
rect 10308 -18116 10391 -18099
rect 10449 -18099 10649 -18061
rect 10449 -18116 10532 -18099
rect 10308 -18133 10324 -18116
rect 10258 -18149 10324 -18133
rect 10516 -18133 10532 -18116
rect 10566 -18116 10649 -18099
rect 10707 -18099 10907 -18061
rect 10707 -18116 10790 -18099
rect 10566 -18133 10582 -18116
rect 10516 -18149 10582 -18133
rect 10774 -18133 10790 -18116
rect 10824 -18116 10907 -18099
rect 10965 -18099 11165 -18061
rect 10965 -18116 11048 -18099
rect 10824 -18133 10840 -18116
rect 10774 -18149 10840 -18133
rect 11032 -18133 11048 -18116
rect 11082 -18116 11165 -18099
rect 11829 -18099 12029 -18061
rect 11829 -18116 11912 -18099
rect 11082 -18133 11098 -18116
rect 11032 -18149 11098 -18133
rect 11896 -18133 11912 -18116
rect 11946 -18116 12029 -18099
rect 12087 -18099 12287 -18061
rect 12087 -18116 12170 -18099
rect 11946 -18133 11962 -18116
rect 11896 -18149 11962 -18133
rect 12154 -18133 12170 -18116
rect 12204 -18116 12287 -18099
rect 12345 -18099 12545 -18061
rect 12345 -18116 12428 -18099
rect 12204 -18133 12220 -18116
rect 12154 -18149 12220 -18133
rect 12412 -18133 12428 -18116
rect 12462 -18116 12545 -18099
rect 12603 -18099 12803 -18061
rect 12603 -18116 12686 -18099
rect 12462 -18133 12478 -18116
rect 12412 -18149 12478 -18133
rect 12670 -18133 12686 -18116
rect 12720 -18116 12803 -18099
rect 12861 -18099 13061 -18061
rect 12861 -18116 12944 -18099
rect 12720 -18133 12736 -18116
rect 12670 -18149 12736 -18133
rect 12928 -18133 12944 -18116
rect 12978 -18116 13061 -18099
rect 13119 -18099 13319 -18061
rect 13119 -18116 13202 -18099
rect 12978 -18133 12994 -18116
rect 12928 -18149 12994 -18133
rect 13186 -18133 13202 -18116
rect 13236 -18116 13319 -18099
rect 13377 -18099 13577 -18061
rect 13377 -18116 13460 -18099
rect 13236 -18133 13252 -18116
rect 13186 -18149 13252 -18133
rect 13444 -18133 13460 -18116
rect 13494 -18116 13577 -18099
rect 13635 -18099 13835 -18061
rect 13635 -18116 13718 -18099
rect 13494 -18133 13510 -18116
rect 13444 -18149 13510 -18133
rect 13702 -18133 13718 -18116
rect 13752 -18116 13835 -18099
rect 14492 -18098 14692 -18060
rect 14492 -18115 14575 -18098
rect 13752 -18133 13768 -18116
rect 13702 -18149 13768 -18133
rect 14559 -18132 14575 -18115
rect 14609 -18115 14692 -18098
rect 14750 -18098 14950 -18060
rect 14750 -18115 14833 -18098
rect 14609 -18132 14625 -18115
rect 14559 -18148 14625 -18132
rect 14817 -18132 14833 -18115
rect 14867 -18115 14950 -18098
rect 15008 -18098 15208 -18060
rect 15008 -18115 15091 -18098
rect 14867 -18132 14883 -18115
rect 14817 -18148 14883 -18132
rect 15075 -18132 15091 -18115
rect 15125 -18115 15208 -18098
rect 15266 -18098 15466 -18060
rect 15266 -18115 15349 -18098
rect 15125 -18132 15141 -18115
rect 15075 -18148 15141 -18132
rect 15333 -18132 15349 -18115
rect 15383 -18115 15466 -18098
rect 15524 -18098 15724 -18060
rect 15524 -18115 15607 -18098
rect 15383 -18132 15399 -18115
rect 15333 -18148 15399 -18132
rect 15591 -18132 15607 -18115
rect 15641 -18115 15724 -18098
rect 15782 -18098 15982 -18060
rect 15782 -18115 15865 -18098
rect 15641 -18132 15657 -18115
rect 15591 -18148 15657 -18132
rect 15849 -18132 15865 -18115
rect 15899 -18115 15982 -18098
rect 16040 -18098 16240 -18060
rect 16040 -18115 16123 -18098
rect 15899 -18132 15915 -18115
rect 15849 -18148 15915 -18132
rect 16107 -18132 16123 -18115
rect 16157 -18115 16240 -18098
rect 16298 -18098 16498 -18060
rect 16298 -18115 16381 -18098
rect 16157 -18132 16173 -18115
rect 16107 -18148 16173 -18132
rect 16365 -18132 16381 -18115
rect 16415 -18115 16498 -18098
rect 16415 -18132 16431 -18115
rect 16365 -18148 16431 -18132
rect 9106 -18441 9172 -18425
rect 9106 -18458 9122 -18441
rect 9039 -18475 9122 -18458
rect 9156 -18458 9172 -18441
rect 9646 -18441 9712 -18425
rect 9646 -18458 9662 -18441
rect 9156 -18475 9239 -18458
rect 9039 -18513 9239 -18475
rect 9579 -18475 9662 -18458
rect 9696 -18458 9712 -18441
rect 10126 -18441 10192 -18425
rect 10126 -18458 10142 -18441
rect 9696 -18475 9779 -18458
rect 9579 -18513 9779 -18475
rect 10059 -18475 10142 -18458
rect 10176 -18458 10192 -18441
rect 10629 -18439 10695 -18423
rect 10629 -18456 10645 -18439
rect 10176 -18475 10259 -18458
rect 10059 -18513 10259 -18475
rect 10562 -18473 10645 -18456
rect 10679 -18456 10695 -18439
rect 11139 -18429 11205 -18413
rect 11139 -18446 11155 -18429
rect 10679 -18473 10762 -18456
rect 10562 -18511 10762 -18473
rect 11072 -18463 11155 -18446
rect 11189 -18446 11205 -18429
rect 11776 -18441 11842 -18425
rect 11189 -18463 11272 -18446
rect 11776 -18458 11792 -18441
rect 11072 -18501 11272 -18463
rect 11709 -18475 11792 -18458
rect 11826 -18458 11842 -18441
rect 12316 -18441 12382 -18425
rect 12316 -18458 12332 -18441
rect 11826 -18475 11909 -18458
rect 11709 -18513 11909 -18475
rect 12249 -18475 12332 -18458
rect 12366 -18458 12382 -18441
rect 12796 -18441 12862 -18425
rect 12796 -18458 12812 -18441
rect 12366 -18475 12449 -18458
rect 12249 -18513 12449 -18475
rect 12729 -18475 12812 -18458
rect 12846 -18458 12862 -18441
rect 13299 -18439 13365 -18423
rect 13299 -18456 13315 -18439
rect 12846 -18475 12929 -18458
rect 12729 -18513 12929 -18475
rect 13232 -18473 13315 -18456
rect 13349 -18456 13365 -18439
rect 13809 -18429 13875 -18413
rect 13809 -18446 13825 -18429
rect 13349 -18473 13432 -18456
rect 13232 -18511 13432 -18473
rect 13742 -18463 13825 -18446
rect 13859 -18446 13875 -18429
rect 14439 -18440 14505 -18424
rect 13859 -18463 13942 -18446
rect 14439 -18457 14455 -18440
rect 13742 -18501 13942 -18463
rect 14372 -18474 14455 -18457
rect 14489 -18457 14505 -18440
rect 14979 -18440 15045 -18424
rect 14979 -18457 14995 -18440
rect 14489 -18474 14572 -18457
rect 9039 -18751 9239 -18713
rect 9039 -18768 9122 -18751
rect 9106 -18785 9122 -18768
rect 9156 -18768 9239 -18751
rect 9579 -18751 9779 -18713
rect 9579 -18768 9662 -18751
rect 9156 -18785 9172 -18768
rect 9106 -18801 9172 -18785
rect 9646 -18785 9662 -18768
rect 9696 -18768 9779 -18751
rect 10059 -18751 10259 -18713
rect 10059 -18768 10142 -18751
rect 9696 -18785 9712 -18768
rect 9646 -18801 9712 -18785
rect 10126 -18785 10142 -18768
rect 10176 -18768 10259 -18751
rect 10562 -18749 10762 -18711
rect 10562 -18766 10645 -18749
rect 10176 -18785 10192 -18768
rect 10126 -18801 10192 -18785
rect 10629 -18783 10645 -18766
rect 10679 -18766 10762 -18749
rect 11072 -18739 11272 -18701
rect 14372 -18512 14572 -18474
rect 14912 -18474 14995 -18457
rect 15029 -18457 15045 -18440
rect 15459 -18440 15525 -18424
rect 15459 -18457 15475 -18440
rect 15029 -18474 15112 -18457
rect 14912 -18512 15112 -18474
rect 15392 -18474 15475 -18457
rect 15509 -18457 15525 -18440
rect 15962 -18438 16028 -18422
rect 15962 -18455 15978 -18438
rect 15509 -18474 15592 -18457
rect 15392 -18512 15592 -18474
rect 15895 -18472 15978 -18455
rect 16012 -18455 16028 -18438
rect 16472 -18428 16538 -18412
rect 16472 -18445 16488 -18428
rect 16012 -18472 16095 -18455
rect 15895 -18510 16095 -18472
rect 16405 -18462 16488 -18445
rect 16522 -18445 16538 -18428
rect 16522 -18462 16605 -18445
rect 16405 -18500 16605 -18462
rect 11072 -18756 11155 -18739
rect 10679 -18783 10695 -18766
rect 10629 -18799 10695 -18783
rect 11139 -18773 11155 -18756
rect 11189 -18756 11272 -18739
rect 11709 -18751 11909 -18713
rect 11189 -18773 11205 -18756
rect 11709 -18768 11792 -18751
rect 11139 -18789 11205 -18773
rect 11776 -18785 11792 -18768
rect 11826 -18768 11909 -18751
rect 12249 -18751 12449 -18713
rect 12249 -18768 12332 -18751
rect 11826 -18785 11842 -18768
rect 11776 -18801 11842 -18785
rect 12316 -18785 12332 -18768
rect 12366 -18768 12449 -18751
rect 12729 -18751 12929 -18713
rect 12729 -18768 12812 -18751
rect 12366 -18785 12382 -18768
rect 12316 -18801 12382 -18785
rect 12796 -18785 12812 -18768
rect 12846 -18768 12929 -18751
rect 13232 -18749 13432 -18711
rect 13232 -18766 13315 -18749
rect 12846 -18785 12862 -18768
rect 12796 -18801 12862 -18785
rect 13299 -18783 13315 -18766
rect 13349 -18766 13432 -18749
rect 13742 -18739 13942 -18701
rect 13742 -18756 13825 -18739
rect 13349 -18783 13365 -18766
rect 13299 -18799 13365 -18783
rect 13809 -18773 13825 -18756
rect 13859 -18756 13942 -18739
rect 14372 -18750 14572 -18712
rect 13859 -18773 13875 -18756
rect 14372 -18767 14455 -18750
rect 13809 -18789 13875 -18773
rect 14439 -18784 14455 -18767
rect 14489 -18767 14572 -18750
rect 14912 -18750 15112 -18712
rect 14912 -18767 14995 -18750
rect 14489 -18784 14505 -18767
rect 14439 -18800 14505 -18784
rect 14979 -18784 14995 -18767
rect 15029 -18767 15112 -18750
rect 15392 -18750 15592 -18712
rect 15392 -18767 15475 -18750
rect 15029 -18784 15045 -18767
rect 14979 -18800 15045 -18784
rect 15459 -18784 15475 -18767
rect 15509 -18767 15592 -18750
rect 15895 -18748 16095 -18710
rect 15895 -18765 15978 -18748
rect 15509 -18784 15525 -18767
rect 15459 -18800 15525 -18784
rect 15962 -18782 15978 -18765
rect 16012 -18765 16095 -18748
rect 16405 -18738 16605 -18700
rect 16405 -18755 16488 -18738
rect 16012 -18782 16028 -18765
rect 15962 -18798 16028 -18782
rect 16472 -18772 16488 -18755
rect 16522 -18755 16605 -18738
rect 16522 -18772 16538 -18755
rect 16472 -18788 16538 -18772
rect 16682 -19541 16748 -19525
rect 16682 -19575 16698 -19541
rect 16732 -19575 16748 -19541
rect 16682 -19591 16748 -19575
rect 16700 -19622 16730 -19591
rect 9429 -20167 9545 -20139
rect 9429 -20205 9453 -20167
rect 9519 -20205 9545 -20167
rect 10044 -20175 10230 -20159
rect 10044 -20192 10060 -20175
rect 9429 -20255 9545 -20205
rect 9737 -20209 10060 -20192
rect 10214 -20192 10230 -20175
rect 10770 -20169 10886 -20141
rect 10214 -20209 10537 -20192
rect 9737 -20256 10537 -20209
rect 10770 -20207 10794 -20169
rect 10860 -20207 10886 -20169
rect 9429 -20429 9545 -20365
rect 10770 -20257 10886 -20207
rect 11140 -20169 11256 -20141
rect 11140 -20207 11164 -20169
rect 11230 -20207 11256 -20169
rect 11140 -20257 11256 -20207
rect 11562 -20169 11678 -20141
rect 11562 -20207 11586 -20169
rect 11652 -20207 11678 -20169
rect 11562 -20257 11678 -20207
rect 11984 -20169 12100 -20141
rect 11984 -20207 12008 -20169
rect 12074 -20207 12100 -20169
rect 12714 -20175 12900 -20159
rect 12714 -20192 12730 -20175
rect 11984 -20257 12100 -20207
rect 12407 -20209 12730 -20192
rect 12884 -20192 12900 -20175
rect 13471 -20169 13587 -20141
rect 12884 -20209 13207 -20192
rect 12407 -20256 13207 -20209
rect 13471 -20207 13495 -20169
rect 13561 -20207 13587 -20169
rect 9737 -20413 10537 -20366
rect 13471 -20257 13587 -20207
rect 13841 -20169 13957 -20141
rect 13841 -20207 13865 -20169
rect 13931 -20207 13957 -20169
rect 13841 -20257 13957 -20207
rect 14263 -20169 14379 -20141
rect 14263 -20207 14287 -20169
rect 14353 -20207 14379 -20169
rect 14263 -20257 14379 -20207
rect 14685 -20169 14801 -20141
rect 14685 -20207 14709 -20169
rect 14775 -20207 14801 -20169
rect 15377 -20174 15563 -20158
rect 15377 -20191 15393 -20174
rect 14685 -20257 14801 -20207
rect 15070 -20208 15393 -20191
rect 15547 -20191 15563 -20174
rect 15547 -20208 15870 -20191
rect 15070 -20255 15870 -20208
rect 9737 -20430 10060 -20413
rect 10044 -20447 10060 -20430
rect 10214 -20430 10537 -20413
rect 10214 -20447 10230 -20430
rect 10770 -20431 10886 -20367
rect 11140 -20431 11256 -20367
rect 11562 -20431 11678 -20367
rect 11984 -20431 12100 -20367
rect 12407 -20413 13207 -20366
rect 12407 -20430 12730 -20413
rect 10044 -20463 10230 -20447
rect 12714 -20447 12730 -20430
rect 12884 -20430 13207 -20413
rect 12884 -20447 12900 -20430
rect 13471 -20431 13587 -20367
rect 13841 -20431 13957 -20367
rect 14263 -20431 14379 -20367
rect 14685 -20431 14801 -20367
rect 15070 -20412 15870 -20365
rect 15070 -20429 15393 -20412
rect 12714 -20463 12900 -20447
rect 15377 -20446 15393 -20429
rect 15547 -20429 15870 -20412
rect 15547 -20446 15563 -20429
rect 15377 -20462 15563 -20446
rect 17072 -19543 17138 -19527
rect 17072 -19577 17088 -19543
rect 17122 -19577 17138 -19543
rect 17072 -19593 17138 -19577
rect 17090 -19624 17120 -19593
rect 16700 -19989 16730 -19958
rect 16682 -20005 16748 -19989
rect 16682 -20039 16698 -20005
rect 16732 -20039 16748 -20005
rect 16682 -20055 16748 -20039
rect 17090 -19991 17120 -19960
rect 17072 -20007 17138 -19991
rect 17072 -20041 17088 -20007
rect 17122 -20041 17138 -20007
rect 17072 -20057 17138 -20041
rect 16686 -20337 16752 -20321
rect 16686 -20371 16702 -20337
rect 16736 -20371 16752 -20337
rect 16686 -20387 16752 -20371
rect 16704 -20409 16734 -20387
rect 17076 -20337 17142 -20321
rect 17076 -20371 17092 -20337
rect 17126 -20371 17142 -20337
rect 17076 -20387 17142 -20371
rect 17094 -20409 17124 -20387
rect 16704 -20515 16734 -20493
rect 16686 -20531 16752 -20515
rect 16686 -20565 16702 -20531
rect 16736 -20565 16752 -20531
rect 16686 -20581 16752 -20565
rect 17094 -20515 17124 -20493
rect 17076 -20531 17142 -20515
rect 17076 -20565 17092 -20531
rect 17126 -20565 17142 -20531
rect 17076 -20581 17142 -20565
rect 9226 -21185 9292 -21169
rect 9226 -21202 9242 -21185
rect 9159 -21219 9242 -21202
rect 9276 -21202 9292 -21185
rect 9484 -21185 9550 -21169
rect 9484 -21202 9500 -21185
rect 9276 -21219 9359 -21202
rect 9159 -21257 9359 -21219
rect 9417 -21219 9500 -21202
rect 9534 -21202 9550 -21185
rect 9742 -21185 9808 -21169
rect 9742 -21202 9758 -21185
rect 9534 -21219 9617 -21202
rect 9417 -21257 9617 -21219
rect 9675 -21219 9758 -21202
rect 9792 -21202 9808 -21185
rect 10000 -21185 10066 -21169
rect 10000 -21202 10016 -21185
rect 9792 -21219 9875 -21202
rect 9675 -21257 9875 -21219
rect 9933 -21219 10016 -21202
rect 10050 -21202 10066 -21185
rect 10258 -21185 10324 -21169
rect 10258 -21202 10274 -21185
rect 10050 -21219 10133 -21202
rect 9933 -21257 10133 -21219
rect 10191 -21219 10274 -21202
rect 10308 -21202 10324 -21185
rect 10516 -21185 10582 -21169
rect 10516 -21202 10532 -21185
rect 10308 -21219 10391 -21202
rect 10191 -21257 10391 -21219
rect 10449 -21219 10532 -21202
rect 10566 -21202 10582 -21185
rect 10774 -21185 10840 -21169
rect 10774 -21202 10790 -21185
rect 10566 -21219 10649 -21202
rect 10449 -21257 10649 -21219
rect 10707 -21219 10790 -21202
rect 10824 -21202 10840 -21185
rect 11032 -21185 11098 -21169
rect 11032 -21202 11048 -21185
rect 10824 -21219 10907 -21202
rect 10707 -21257 10907 -21219
rect 10965 -21219 11048 -21202
rect 11082 -21202 11098 -21185
rect 11896 -21185 11962 -21169
rect 11896 -21202 11912 -21185
rect 11082 -21219 11165 -21202
rect 10965 -21257 11165 -21219
rect 11829 -21219 11912 -21202
rect 11946 -21202 11962 -21185
rect 12154 -21185 12220 -21169
rect 12154 -21202 12170 -21185
rect 11946 -21219 12029 -21202
rect 11829 -21257 12029 -21219
rect 12087 -21219 12170 -21202
rect 12204 -21202 12220 -21185
rect 12412 -21185 12478 -21169
rect 12412 -21202 12428 -21185
rect 12204 -21219 12287 -21202
rect 12087 -21257 12287 -21219
rect 12345 -21219 12428 -21202
rect 12462 -21202 12478 -21185
rect 12670 -21185 12736 -21169
rect 12670 -21202 12686 -21185
rect 12462 -21219 12545 -21202
rect 12345 -21257 12545 -21219
rect 12603 -21219 12686 -21202
rect 12720 -21202 12736 -21185
rect 12928 -21185 12994 -21169
rect 12928 -21202 12944 -21185
rect 12720 -21219 12803 -21202
rect 12603 -21257 12803 -21219
rect 12861 -21219 12944 -21202
rect 12978 -21202 12994 -21185
rect 13186 -21185 13252 -21169
rect 13186 -21202 13202 -21185
rect 12978 -21219 13061 -21202
rect 12861 -21257 13061 -21219
rect 13119 -21219 13202 -21202
rect 13236 -21202 13252 -21185
rect 13444 -21185 13510 -21169
rect 13444 -21202 13460 -21185
rect 13236 -21219 13319 -21202
rect 13119 -21257 13319 -21219
rect 13377 -21219 13460 -21202
rect 13494 -21202 13510 -21185
rect 13702 -21185 13768 -21169
rect 13702 -21202 13718 -21185
rect 13494 -21219 13577 -21202
rect 13377 -21257 13577 -21219
rect 13635 -21219 13718 -21202
rect 13752 -21202 13768 -21185
rect 14559 -21184 14625 -21168
rect 14559 -21201 14575 -21184
rect 13752 -21219 13835 -21202
rect 13635 -21257 13835 -21219
rect 14492 -21218 14575 -21201
rect 14609 -21201 14625 -21184
rect 14817 -21184 14883 -21168
rect 14817 -21201 14833 -21184
rect 14609 -21218 14692 -21201
rect 14492 -21256 14692 -21218
rect 14750 -21218 14833 -21201
rect 14867 -21201 14883 -21184
rect 15075 -21184 15141 -21168
rect 15075 -21201 15091 -21184
rect 14867 -21218 14950 -21201
rect 14750 -21256 14950 -21218
rect 15008 -21218 15091 -21201
rect 15125 -21201 15141 -21184
rect 15333 -21184 15399 -21168
rect 15333 -21201 15349 -21184
rect 15125 -21218 15208 -21201
rect 15008 -21256 15208 -21218
rect 15266 -21218 15349 -21201
rect 15383 -21201 15399 -21184
rect 15591 -21184 15657 -21168
rect 15591 -21201 15607 -21184
rect 15383 -21218 15466 -21201
rect 15266 -21256 15466 -21218
rect 15524 -21218 15607 -21201
rect 15641 -21201 15657 -21184
rect 15849 -21184 15915 -21168
rect 15849 -21201 15865 -21184
rect 15641 -21218 15724 -21201
rect 15524 -21256 15724 -21218
rect 15782 -21218 15865 -21201
rect 15899 -21201 15915 -21184
rect 16107 -21184 16173 -21168
rect 16107 -21201 16123 -21184
rect 15899 -21218 15982 -21201
rect 15782 -21256 15982 -21218
rect 16040 -21218 16123 -21201
rect 16157 -21201 16173 -21184
rect 16365 -21184 16431 -21168
rect 16365 -21201 16381 -21184
rect 16157 -21218 16240 -21201
rect 16040 -21256 16240 -21218
rect 16298 -21218 16381 -21201
rect 16415 -21201 16431 -21184
rect 16415 -21218 16498 -21201
rect 16298 -21256 16498 -21218
rect 9159 -21495 9359 -21457
rect 9159 -21512 9242 -21495
rect 9226 -21529 9242 -21512
rect 9276 -21512 9359 -21495
rect 9417 -21495 9617 -21457
rect 9417 -21512 9500 -21495
rect 9276 -21529 9292 -21512
rect 9226 -21545 9292 -21529
rect 9484 -21529 9500 -21512
rect 9534 -21512 9617 -21495
rect 9675 -21495 9875 -21457
rect 9675 -21512 9758 -21495
rect 9534 -21529 9550 -21512
rect 9484 -21545 9550 -21529
rect 9742 -21529 9758 -21512
rect 9792 -21512 9875 -21495
rect 9933 -21495 10133 -21457
rect 9933 -21512 10016 -21495
rect 9792 -21529 9808 -21512
rect 9742 -21545 9808 -21529
rect 10000 -21529 10016 -21512
rect 10050 -21512 10133 -21495
rect 10191 -21495 10391 -21457
rect 10191 -21512 10274 -21495
rect 10050 -21529 10066 -21512
rect 10000 -21545 10066 -21529
rect 10258 -21529 10274 -21512
rect 10308 -21512 10391 -21495
rect 10449 -21495 10649 -21457
rect 10449 -21512 10532 -21495
rect 10308 -21529 10324 -21512
rect 10258 -21545 10324 -21529
rect 10516 -21529 10532 -21512
rect 10566 -21512 10649 -21495
rect 10707 -21495 10907 -21457
rect 10707 -21512 10790 -21495
rect 10566 -21529 10582 -21512
rect 10516 -21545 10582 -21529
rect 10774 -21529 10790 -21512
rect 10824 -21512 10907 -21495
rect 10965 -21495 11165 -21457
rect 10965 -21512 11048 -21495
rect 10824 -21529 10840 -21512
rect 10774 -21545 10840 -21529
rect 11032 -21529 11048 -21512
rect 11082 -21512 11165 -21495
rect 11829 -21495 12029 -21457
rect 11829 -21512 11912 -21495
rect 11082 -21529 11098 -21512
rect 11032 -21545 11098 -21529
rect 11896 -21529 11912 -21512
rect 11946 -21512 12029 -21495
rect 12087 -21495 12287 -21457
rect 12087 -21512 12170 -21495
rect 11946 -21529 11962 -21512
rect 11896 -21545 11962 -21529
rect 12154 -21529 12170 -21512
rect 12204 -21512 12287 -21495
rect 12345 -21495 12545 -21457
rect 12345 -21512 12428 -21495
rect 12204 -21529 12220 -21512
rect 12154 -21545 12220 -21529
rect 12412 -21529 12428 -21512
rect 12462 -21512 12545 -21495
rect 12603 -21495 12803 -21457
rect 12603 -21512 12686 -21495
rect 12462 -21529 12478 -21512
rect 12412 -21545 12478 -21529
rect 12670 -21529 12686 -21512
rect 12720 -21512 12803 -21495
rect 12861 -21495 13061 -21457
rect 12861 -21512 12944 -21495
rect 12720 -21529 12736 -21512
rect 12670 -21545 12736 -21529
rect 12928 -21529 12944 -21512
rect 12978 -21512 13061 -21495
rect 13119 -21495 13319 -21457
rect 13119 -21512 13202 -21495
rect 12978 -21529 12994 -21512
rect 12928 -21545 12994 -21529
rect 13186 -21529 13202 -21512
rect 13236 -21512 13319 -21495
rect 13377 -21495 13577 -21457
rect 13377 -21512 13460 -21495
rect 13236 -21529 13252 -21512
rect 13186 -21545 13252 -21529
rect 13444 -21529 13460 -21512
rect 13494 -21512 13577 -21495
rect 13635 -21495 13835 -21457
rect 13635 -21512 13718 -21495
rect 13494 -21529 13510 -21512
rect 13444 -21545 13510 -21529
rect 13702 -21529 13718 -21512
rect 13752 -21512 13835 -21495
rect 14492 -21494 14692 -21456
rect 14492 -21511 14575 -21494
rect 13752 -21529 13768 -21512
rect 13702 -21545 13768 -21529
rect 14559 -21528 14575 -21511
rect 14609 -21511 14692 -21494
rect 14750 -21494 14950 -21456
rect 14750 -21511 14833 -21494
rect 14609 -21528 14625 -21511
rect 14559 -21544 14625 -21528
rect 14817 -21528 14833 -21511
rect 14867 -21511 14950 -21494
rect 15008 -21494 15208 -21456
rect 15008 -21511 15091 -21494
rect 14867 -21528 14883 -21511
rect 14817 -21544 14883 -21528
rect 15075 -21528 15091 -21511
rect 15125 -21511 15208 -21494
rect 15266 -21494 15466 -21456
rect 15266 -21511 15349 -21494
rect 15125 -21528 15141 -21511
rect 15075 -21544 15141 -21528
rect 15333 -21528 15349 -21511
rect 15383 -21511 15466 -21494
rect 15524 -21494 15724 -21456
rect 15524 -21511 15607 -21494
rect 15383 -21528 15399 -21511
rect 15333 -21544 15399 -21528
rect 15591 -21528 15607 -21511
rect 15641 -21511 15724 -21494
rect 15782 -21494 15982 -21456
rect 15782 -21511 15865 -21494
rect 15641 -21528 15657 -21511
rect 15591 -21544 15657 -21528
rect 15849 -21528 15865 -21511
rect 15899 -21511 15982 -21494
rect 16040 -21494 16240 -21456
rect 16040 -21511 16123 -21494
rect 15899 -21528 15915 -21511
rect 15849 -21544 15915 -21528
rect 16107 -21528 16123 -21511
rect 16157 -21511 16240 -21494
rect 16298 -21494 16498 -21456
rect 16298 -21511 16381 -21494
rect 16157 -21528 16173 -21511
rect 16107 -21544 16173 -21528
rect 16365 -21528 16381 -21511
rect 16415 -21511 16498 -21494
rect 16415 -21528 16431 -21511
rect 16365 -21544 16431 -21528
rect 9226 -21603 9292 -21587
rect 9226 -21620 9242 -21603
rect 9159 -21637 9242 -21620
rect 9276 -21620 9292 -21603
rect 9484 -21603 9550 -21587
rect 9484 -21620 9500 -21603
rect 9276 -21637 9359 -21620
rect 9159 -21675 9359 -21637
rect 9417 -21637 9500 -21620
rect 9534 -21620 9550 -21603
rect 9742 -21603 9808 -21587
rect 9742 -21620 9758 -21603
rect 9534 -21637 9617 -21620
rect 9417 -21675 9617 -21637
rect 9675 -21637 9758 -21620
rect 9792 -21620 9808 -21603
rect 10000 -21603 10066 -21587
rect 10000 -21620 10016 -21603
rect 9792 -21637 9875 -21620
rect 9675 -21675 9875 -21637
rect 9933 -21637 10016 -21620
rect 10050 -21620 10066 -21603
rect 10258 -21603 10324 -21587
rect 10258 -21620 10274 -21603
rect 10050 -21637 10133 -21620
rect 9933 -21675 10133 -21637
rect 10191 -21637 10274 -21620
rect 10308 -21620 10324 -21603
rect 10516 -21603 10582 -21587
rect 10516 -21620 10532 -21603
rect 10308 -21637 10391 -21620
rect 10191 -21675 10391 -21637
rect 10449 -21637 10532 -21620
rect 10566 -21620 10582 -21603
rect 10774 -21603 10840 -21587
rect 10774 -21620 10790 -21603
rect 10566 -21637 10649 -21620
rect 10449 -21675 10649 -21637
rect 10707 -21637 10790 -21620
rect 10824 -21620 10840 -21603
rect 11032 -21603 11098 -21587
rect 11032 -21620 11048 -21603
rect 10824 -21637 10907 -21620
rect 10707 -21675 10907 -21637
rect 10965 -21637 11048 -21620
rect 11082 -21620 11098 -21603
rect 11896 -21603 11962 -21587
rect 11896 -21620 11912 -21603
rect 11082 -21637 11165 -21620
rect 10965 -21675 11165 -21637
rect 11829 -21637 11912 -21620
rect 11946 -21620 11962 -21603
rect 12154 -21603 12220 -21587
rect 12154 -21620 12170 -21603
rect 11946 -21637 12029 -21620
rect 11829 -21675 12029 -21637
rect 12087 -21637 12170 -21620
rect 12204 -21620 12220 -21603
rect 12412 -21603 12478 -21587
rect 12412 -21620 12428 -21603
rect 12204 -21637 12287 -21620
rect 12087 -21675 12287 -21637
rect 12345 -21637 12428 -21620
rect 12462 -21620 12478 -21603
rect 12670 -21603 12736 -21587
rect 12670 -21620 12686 -21603
rect 12462 -21637 12545 -21620
rect 12345 -21675 12545 -21637
rect 12603 -21637 12686 -21620
rect 12720 -21620 12736 -21603
rect 12928 -21603 12994 -21587
rect 12928 -21620 12944 -21603
rect 12720 -21637 12803 -21620
rect 12603 -21675 12803 -21637
rect 12861 -21637 12944 -21620
rect 12978 -21620 12994 -21603
rect 13186 -21603 13252 -21587
rect 13186 -21620 13202 -21603
rect 12978 -21637 13061 -21620
rect 12861 -21675 13061 -21637
rect 13119 -21637 13202 -21620
rect 13236 -21620 13252 -21603
rect 13444 -21603 13510 -21587
rect 13444 -21620 13460 -21603
rect 13236 -21637 13319 -21620
rect 13119 -21675 13319 -21637
rect 13377 -21637 13460 -21620
rect 13494 -21620 13510 -21603
rect 13702 -21603 13768 -21587
rect 13702 -21620 13718 -21603
rect 13494 -21637 13577 -21620
rect 13377 -21675 13577 -21637
rect 13635 -21637 13718 -21620
rect 13752 -21620 13768 -21603
rect 14559 -21602 14625 -21586
rect 14559 -21619 14575 -21602
rect 13752 -21637 13835 -21620
rect 13635 -21675 13835 -21637
rect 14492 -21636 14575 -21619
rect 14609 -21619 14625 -21602
rect 14817 -21602 14883 -21586
rect 14817 -21619 14833 -21602
rect 14609 -21636 14692 -21619
rect 14492 -21674 14692 -21636
rect 14750 -21636 14833 -21619
rect 14867 -21619 14883 -21602
rect 15075 -21602 15141 -21586
rect 15075 -21619 15091 -21602
rect 14867 -21636 14950 -21619
rect 14750 -21674 14950 -21636
rect 15008 -21636 15091 -21619
rect 15125 -21619 15141 -21602
rect 15333 -21602 15399 -21586
rect 15333 -21619 15349 -21602
rect 15125 -21636 15208 -21619
rect 15008 -21674 15208 -21636
rect 15266 -21636 15349 -21619
rect 15383 -21619 15399 -21602
rect 15591 -21602 15657 -21586
rect 15591 -21619 15607 -21602
rect 15383 -21636 15466 -21619
rect 15266 -21674 15466 -21636
rect 15524 -21636 15607 -21619
rect 15641 -21619 15657 -21602
rect 15849 -21602 15915 -21586
rect 15849 -21619 15865 -21602
rect 15641 -21636 15724 -21619
rect 15524 -21674 15724 -21636
rect 15782 -21636 15865 -21619
rect 15899 -21619 15915 -21602
rect 16107 -21602 16173 -21586
rect 16107 -21619 16123 -21602
rect 15899 -21636 15982 -21619
rect 15782 -21674 15982 -21636
rect 16040 -21636 16123 -21619
rect 16157 -21619 16173 -21602
rect 16365 -21602 16431 -21586
rect 16365 -21619 16381 -21602
rect 16157 -21636 16240 -21619
rect 16040 -21674 16240 -21636
rect 16298 -21636 16381 -21619
rect 16415 -21619 16431 -21602
rect 16415 -21636 16498 -21619
rect 16298 -21674 16498 -21636
rect 9159 -21913 9359 -21875
rect 9159 -21930 9242 -21913
rect 9226 -21947 9242 -21930
rect 9276 -21930 9359 -21913
rect 9417 -21913 9617 -21875
rect 9417 -21930 9500 -21913
rect 9276 -21947 9292 -21930
rect 9226 -21963 9292 -21947
rect 9484 -21947 9500 -21930
rect 9534 -21930 9617 -21913
rect 9675 -21913 9875 -21875
rect 9675 -21930 9758 -21913
rect 9534 -21947 9550 -21930
rect 9484 -21963 9550 -21947
rect 9742 -21947 9758 -21930
rect 9792 -21930 9875 -21913
rect 9933 -21913 10133 -21875
rect 9933 -21930 10016 -21913
rect 9792 -21947 9808 -21930
rect 9742 -21963 9808 -21947
rect 10000 -21947 10016 -21930
rect 10050 -21930 10133 -21913
rect 10191 -21913 10391 -21875
rect 10191 -21930 10274 -21913
rect 10050 -21947 10066 -21930
rect 10000 -21963 10066 -21947
rect 10258 -21947 10274 -21930
rect 10308 -21930 10391 -21913
rect 10449 -21913 10649 -21875
rect 10449 -21930 10532 -21913
rect 10308 -21947 10324 -21930
rect 10258 -21963 10324 -21947
rect 10516 -21947 10532 -21930
rect 10566 -21930 10649 -21913
rect 10707 -21913 10907 -21875
rect 10707 -21930 10790 -21913
rect 10566 -21947 10582 -21930
rect 10516 -21963 10582 -21947
rect 10774 -21947 10790 -21930
rect 10824 -21930 10907 -21913
rect 10965 -21913 11165 -21875
rect 10965 -21930 11048 -21913
rect 10824 -21947 10840 -21930
rect 10774 -21963 10840 -21947
rect 11032 -21947 11048 -21930
rect 11082 -21930 11165 -21913
rect 11829 -21913 12029 -21875
rect 11829 -21930 11912 -21913
rect 11082 -21947 11098 -21930
rect 11032 -21963 11098 -21947
rect 11896 -21947 11912 -21930
rect 11946 -21930 12029 -21913
rect 12087 -21913 12287 -21875
rect 12087 -21930 12170 -21913
rect 11946 -21947 11962 -21930
rect 11896 -21963 11962 -21947
rect 12154 -21947 12170 -21930
rect 12204 -21930 12287 -21913
rect 12345 -21913 12545 -21875
rect 12345 -21930 12428 -21913
rect 12204 -21947 12220 -21930
rect 12154 -21963 12220 -21947
rect 12412 -21947 12428 -21930
rect 12462 -21930 12545 -21913
rect 12603 -21913 12803 -21875
rect 12603 -21930 12686 -21913
rect 12462 -21947 12478 -21930
rect 12412 -21963 12478 -21947
rect 12670 -21947 12686 -21930
rect 12720 -21930 12803 -21913
rect 12861 -21913 13061 -21875
rect 12861 -21930 12944 -21913
rect 12720 -21947 12736 -21930
rect 12670 -21963 12736 -21947
rect 12928 -21947 12944 -21930
rect 12978 -21930 13061 -21913
rect 13119 -21913 13319 -21875
rect 13119 -21930 13202 -21913
rect 12978 -21947 12994 -21930
rect 12928 -21963 12994 -21947
rect 13186 -21947 13202 -21930
rect 13236 -21930 13319 -21913
rect 13377 -21913 13577 -21875
rect 13377 -21930 13460 -21913
rect 13236 -21947 13252 -21930
rect 13186 -21963 13252 -21947
rect 13444 -21947 13460 -21930
rect 13494 -21930 13577 -21913
rect 13635 -21913 13835 -21875
rect 13635 -21930 13718 -21913
rect 13494 -21947 13510 -21930
rect 13444 -21963 13510 -21947
rect 13702 -21947 13718 -21930
rect 13752 -21930 13835 -21913
rect 14492 -21912 14692 -21874
rect 14492 -21929 14575 -21912
rect 13752 -21947 13768 -21930
rect 13702 -21963 13768 -21947
rect 14559 -21946 14575 -21929
rect 14609 -21929 14692 -21912
rect 14750 -21912 14950 -21874
rect 14750 -21929 14833 -21912
rect 14609 -21946 14625 -21929
rect 14559 -21962 14625 -21946
rect 14817 -21946 14833 -21929
rect 14867 -21929 14950 -21912
rect 15008 -21912 15208 -21874
rect 15008 -21929 15091 -21912
rect 14867 -21946 14883 -21929
rect 14817 -21962 14883 -21946
rect 15075 -21946 15091 -21929
rect 15125 -21929 15208 -21912
rect 15266 -21912 15466 -21874
rect 15266 -21929 15349 -21912
rect 15125 -21946 15141 -21929
rect 15075 -21962 15141 -21946
rect 15333 -21946 15349 -21929
rect 15383 -21929 15466 -21912
rect 15524 -21912 15724 -21874
rect 15524 -21929 15607 -21912
rect 15383 -21946 15399 -21929
rect 15333 -21962 15399 -21946
rect 15591 -21946 15607 -21929
rect 15641 -21929 15724 -21912
rect 15782 -21912 15982 -21874
rect 15782 -21929 15865 -21912
rect 15641 -21946 15657 -21929
rect 15591 -21962 15657 -21946
rect 15849 -21946 15865 -21929
rect 15899 -21929 15982 -21912
rect 16040 -21912 16240 -21874
rect 16040 -21929 16123 -21912
rect 15899 -21946 15915 -21929
rect 15849 -21962 15915 -21946
rect 16107 -21946 16123 -21929
rect 16157 -21929 16240 -21912
rect 16298 -21912 16498 -21874
rect 16298 -21929 16381 -21912
rect 16157 -21946 16173 -21929
rect 16107 -21962 16173 -21946
rect 16365 -21946 16381 -21929
rect 16415 -21929 16498 -21912
rect 16415 -21946 16431 -21929
rect 16365 -21962 16431 -21946
rect 9226 -22021 9292 -22005
rect 9226 -22038 9242 -22021
rect 9159 -22055 9242 -22038
rect 9276 -22038 9292 -22021
rect 9484 -22021 9550 -22005
rect 9484 -22038 9500 -22021
rect 9276 -22055 9359 -22038
rect 9159 -22093 9359 -22055
rect 9417 -22055 9500 -22038
rect 9534 -22038 9550 -22021
rect 9742 -22021 9808 -22005
rect 9742 -22038 9758 -22021
rect 9534 -22055 9617 -22038
rect 9417 -22093 9617 -22055
rect 9675 -22055 9758 -22038
rect 9792 -22038 9808 -22021
rect 10000 -22021 10066 -22005
rect 10000 -22038 10016 -22021
rect 9792 -22055 9875 -22038
rect 9675 -22093 9875 -22055
rect 9933 -22055 10016 -22038
rect 10050 -22038 10066 -22021
rect 10258 -22021 10324 -22005
rect 10258 -22038 10274 -22021
rect 10050 -22055 10133 -22038
rect 9933 -22093 10133 -22055
rect 10191 -22055 10274 -22038
rect 10308 -22038 10324 -22021
rect 10516 -22021 10582 -22005
rect 10516 -22038 10532 -22021
rect 10308 -22055 10391 -22038
rect 10191 -22093 10391 -22055
rect 10449 -22055 10532 -22038
rect 10566 -22038 10582 -22021
rect 10774 -22021 10840 -22005
rect 10774 -22038 10790 -22021
rect 10566 -22055 10649 -22038
rect 10449 -22093 10649 -22055
rect 10707 -22055 10790 -22038
rect 10824 -22038 10840 -22021
rect 11032 -22021 11098 -22005
rect 11032 -22038 11048 -22021
rect 10824 -22055 10907 -22038
rect 10707 -22093 10907 -22055
rect 10965 -22055 11048 -22038
rect 11082 -22038 11098 -22021
rect 11896 -22021 11962 -22005
rect 11896 -22038 11912 -22021
rect 11082 -22055 11165 -22038
rect 10965 -22093 11165 -22055
rect 11829 -22055 11912 -22038
rect 11946 -22038 11962 -22021
rect 12154 -22021 12220 -22005
rect 12154 -22038 12170 -22021
rect 11946 -22055 12029 -22038
rect 11829 -22093 12029 -22055
rect 12087 -22055 12170 -22038
rect 12204 -22038 12220 -22021
rect 12412 -22021 12478 -22005
rect 12412 -22038 12428 -22021
rect 12204 -22055 12287 -22038
rect 12087 -22093 12287 -22055
rect 12345 -22055 12428 -22038
rect 12462 -22038 12478 -22021
rect 12670 -22021 12736 -22005
rect 12670 -22038 12686 -22021
rect 12462 -22055 12545 -22038
rect 12345 -22093 12545 -22055
rect 12603 -22055 12686 -22038
rect 12720 -22038 12736 -22021
rect 12928 -22021 12994 -22005
rect 12928 -22038 12944 -22021
rect 12720 -22055 12803 -22038
rect 12603 -22093 12803 -22055
rect 12861 -22055 12944 -22038
rect 12978 -22038 12994 -22021
rect 13186 -22021 13252 -22005
rect 13186 -22038 13202 -22021
rect 12978 -22055 13061 -22038
rect 12861 -22093 13061 -22055
rect 13119 -22055 13202 -22038
rect 13236 -22038 13252 -22021
rect 13444 -22021 13510 -22005
rect 13444 -22038 13460 -22021
rect 13236 -22055 13319 -22038
rect 13119 -22093 13319 -22055
rect 13377 -22055 13460 -22038
rect 13494 -22038 13510 -22021
rect 13702 -22021 13768 -22005
rect 13702 -22038 13718 -22021
rect 13494 -22055 13577 -22038
rect 13377 -22093 13577 -22055
rect 13635 -22055 13718 -22038
rect 13752 -22038 13768 -22021
rect 14559 -22020 14625 -22004
rect 14559 -22037 14575 -22020
rect 13752 -22055 13835 -22038
rect 13635 -22093 13835 -22055
rect 14492 -22054 14575 -22037
rect 14609 -22037 14625 -22020
rect 14817 -22020 14883 -22004
rect 14817 -22037 14833 -22020
rect 14609 -22054 14692 -22037
rect 14492 -22092 14692 -22054
rect 14750 -22054 14833 -22037
rect 14867 -22037 14883 -22020
rect 15075 -22020 15141 -22004
rect 15075 -22037 15091 -22020
rect 14867 -22054 14950 -22037
rect 14750 -22092 14950 -22054
rect 15008 -22054 15091 -22037
rect 15125 -22037 15141 -22020
rect 15333 -22020 15399 -22004
rect 15333 -22037 15349 -22020
rect 15125 -22054 15208 -22037
rect 15008 -22092 15208 -22054
rect 15266 -22054 15349 -22037
rect 15383 -22037 15399 -22020
rect 15591 -22020 15657 -22004
rect 15591 -22037 15607 -22020
rect 15383 -22054 15466 -22037
rect 15266 -22092 15466 -22054
rect 15524 -22054 15607 -22037
rect 15641 -22037 15657 -22020
rect 15849 -22020 15915 -22004
rect 15849 -22037 15865 -22020
rect 15641 -22054 15724 -22037
rect 15524 -22092 15724 -22054
rect 15782 -22054 15865 -22037
rect 15899 -22037 15915 -22020
rect 16107 -22020 16173 -22004
rect 16107 -22037 16123 -22020
rect 15899 -22054 15982 -22037
rect 15782 -22092 15982 -22054
rect 16040 -22054 16123 -22037
rect 16157 -22037 16173 -22020
rect 16365 -22020 16431 -22004
rect 16365 -22037 16381 -22020
rect 16157 -22054 16240 -22037
rect 16040 -22092 16240 -22054
rect 16298 -22054 16381 -22037
rect 16415 -22037 16431 -22020
rect 16415 -22054 16498 -22037
rect 16298 -22092 16498 -22054
rect 9159 -22331 9359 -22293
rect 9159 -22348 9242 -22331
rect 9226 -22365 9242 -22348
rect 9276 -22348 9359 -22331
rect 9417 -22331 9617 -22293
rect 9417 -22348 9500 -22331
rect 9276 -22365 9292 -22348
rect 9226 -22381 9292 -22365
rect 9484 -22365 9500 -22348
rect 9534 -22348 9617 -22331
rect 9675 -22331 9875 -22293
rect 9675 -22348 9758 -22331
rect 9534 -22365 9550 -22348
rect 9484 -22381 9550 -22365
rect 9742 -22365 9758 -22348
rect 9792 -22348 9875 -22331
rect 9933 -22331 10133 -22293
rect 9933 -22348 10016 -22331
rect 9792 -22365 9808 -22348
rect 9742 -22381 9808 -22365
rect 10000 -22365 10016 -22348
rect 10050 -22348 10133 -22331
rect 10191 -22331 10391 -22293
rect 10191 -22348 10274 -22331
rect 10050 -22365 10066 -22348
rect 10000 -22381 10066 -22365
rect 10258 -22365 10274 -22348
rect 10308 -22348 10391 -22331
rect 10449 -22331 10649 -22293
rect 10449 -22348 10532 -22331
rect 10308 -22365 10324 -22348
rect 10258 -22381 10324 -22365
rect 10516 -22365 10532 -22348
rect 10566 -22348 10649 -22331
rect 10707 -22331 10907 -22293
rect 10707 -22348 10790 -22331
rect 10566 -22365 10582 -22348
rect 10516 -22381 10582 -22365
rect 10774 -22365 10790 -22348
rect 10824 -22348 10907 -22331
rect 10965 -22331 11165 -22293
rect 10965 -22348 11048 -22331
rect 10824 -22365 10840 -22348
rect 10774 -22381 10840 -22365
rect 11032 -22365 11048 -22348
rect 11082 -22348 11165 -22331
rect 11829 -22331 12029 -22293
rect 11829 -22348 11912 -22331
rect 11082 -22365 11098 -22348
rect 11032 -22381 11098 -22365
rect 11896 -22365 11912 -22348
rect 11946 -22348 12029 -22331
rect 12087 -22331 12287 -22293
rect 12087 -22348 12170 -22331
rect 11946 -22365 11962 -22348
rect 11896 -22381 11962 -22365
rect 12154 -22365 12170 -22348
rect 12204 -22348 12287 -22331
rect 12345 -22331 12545 -22293
rect 12345 -22348 12428 -22331
rect 12204 -22365 12220 -22348
rect 12154 -22381 12220 -22365
rect 12412 -22365 12428 -22348
rect 12462 -22348 12545 -22331
rect 12603 -22331 12803 -22293
rect 12603 -22348 12686 -22331
rect 12462 -22365 12478 -22348
rect 12412 -22381 12478 -22365
rect 12670 -22365 12686 -22348
rect 12720 -22348 12803 -22331
rect 12861 -22331 13061 -22293
rect 12861 -22348 12944 -22331
rect 12720 -22365 12736 -22348
rect 12670 -22381 12736 -22365
rect 12928 -22365 12944 -22348
rect 12978 -22348 13061 -22331
rect 13119 -22331 13319 -22293
rect 13119 -22348 13202 -22331
rect 12978 -22365 12994 -22348
rect 12928 -22381 12994 -22365
rect 13186 -22365 13202 -22348
rect 13236 -22348 13319 -22331
rect 13377 -22331 13577 -22293
rect 13377 -22348 13460 -22331
rect 13236 -22365 13252 -22348
rect 13186 -22381 13252 -22365
rect 13444 -22365 13460 -22348
rect 13494 -22348 13577 -22331
rect 13635 -22331 13835 -22293
rect 13635 -22348 13718 -22331
rect 13494 -22365 13510 -22348
rect 13444 -22381 13510 -22365
rect 13702 -22365 13718 -22348
rect 13752 -22348 13835 -22331
rect 14492 -22330 14692 -22292
rect 14492 -22347 14575 -22330
rect 13752 -22365 13768 -22348
rect 13702 -22381 13768 -22365
rect 14559 -22364 14575 -22347
rect 14609 -22347 14692 -22330
rect 14750 -22330 14950 -22292
rect 14750 -22347 14833 -22330
rect 14609 -22364 14625 -22347
rect 14559 -22380 14625 -22364
rect 14817 -22364 14833 -22347
rect 14867 -22347 14950 -22330
rect 15008 -22330 15208 -22292
rect 15008 -22347 15091 -22330
rect 14867 -22364 14883 -22347
rect 14817 -22380 14883 -22364
rect 15075 -22364 15091 -22347
rect 15125 -22347 15208 -22330
rect 15266 -22330 15466 -22292
rect 15266 -22347 15349 -22330
rect 15125 -22364 15141 -22347
rect 15075 -22380 15141 -22364
rect 15333 -22364 15349 -22347
rect 15383 -22347 15466 -22330
rect 15524 -22330 15724 -22292
rect 15524 -22347 15607 -22330
rect 15383 -22364 15399 -22347
rect 15333 -22380 15399 -22364
rect 15591 -22364 15607 -22347
rect 15641 -22347 15724 -22330
rect 15782 -22330 15982 -22292
rect 15782 -22347 15865 -22330
rect 15641 -22364 15657 -22347
rect 15591 -22380 15657 -22364
rect 15849 -22364 15865 -22347
rect 15899 -22347 15982 -22330
rect 16040 -22330 16240 -22292
rect 16040 -22347 16123 -22330
rect 15899 -22364 15915 -22347
rect 15849 -22380 15915 -22364
rect 16107 -22364 16123 -22347
rect 16157 -22347 16240 -22330
rect 16298 -22330 16498 -22292
rect 16298 -22347 16381 -22330
rect 16157 -22364 16173 -22347
rect 16107 -22380 16173 -22364
rect 16365 -22364 16381 -22347
rect 16415 -22347 16498 -22330
rect 16415 -22364 16431 -22347
rect 16365 -22380 16431 -22364
rect 9226 -22439 9292 -22423
rect 9226 -22456 9242 -22439
rect 9159 -22473 9242 -22456
rect 9276 -22456 9292 -22439
rect 9484 -22439 9550 -22423
rect 9484 -22456 9500 -22439
rect 9276 -22473 9359 -22456
rect 9159 -22511 9359 -22473
rect 9417 -22473 9500 -22456
rect 9534 -22456 9550 -22439
rect 9742 -22439 9808 -22423
rect 9742 -22456 9758 -22439
rect 9534 -22473 9617 -22456
rect 9417 -22511 9617 -22473
rect 9675 -22473 9758 -22456
rect 9792 -22456 9808 -22439
rect 10000 -22439 10066 -22423
rect 10000 -22456 10016 -22439
rect 9792 -22473 9875 -22456
rect 9675 -22511 9875 -22473
rect 9933 -22473 10016 -22456
rect 10050 -22456 10066 -22439
rect 10258 -22439 10324 -22423
rect 10258 -22456 10274 -22439
rect 10050 -22473 10133 -22456
rect 9933 -22511 10133 -22473
rect 10191 -22473 10274 -22456
rect 10308 -22456 10324 -22439
rect 10516 -22439 10582 -22423
rect 10516 -22456 10532 -22439
rect 10308 -22473 10391 -22456
rect 10191 -22511 10391 -22473
rect 10449 -22473 10532 -22456
rect 10566 -22456 10582 -22439
rect 10774 -22439 10840 -22423
rect 10774 -22456 10790 -22439
rect 10566 -22473 10649 -22456
rect 10449 -22511 10649 -22473
rect 10707 -22473 10790 -22456
rect 10824 -22456 10840 -22439
rect 11032 -22439 11098 -22423
rect 11032 -22456 11048 -22439
rect 10824 -22473 10907 -22456
rect 10707 -22511 10907 -22473
rect 10965 -22473 11048 -22456
rect 11082 -22456 11098 -22439
rect 11896 -22439 11962 -22423
rect 11896 -22456 11912 -22439
rect 11082 -22473 11165 -22456
rect 10965 -22511 11165 -22473
rect 11829 -22473 11912 -22456
rect 11946 -22456 11962 -22439
rect 12154 -22439 12220 -22423
rect 12154 -22456 12170 -22439
rect 11946 -22473 12029 -22456
rect 11829 -22511 12029 -22473
rect 12087 -22473 12170 -22456
rect 12204 -22456 12220 -22439
rect 12412 -22439 12478 -22423
rect 12412 -22456 12428 -22439
rect 12204 -22473 12287 -22456
rect 12087 -22511 12287 -22473
rect 12345 -22473 12428 -22456
rect 12462 -22456 12478 -22439
rect 12670 -22439 12736 -22423
rect 12670 -22456 12686 -22439
rect 12462 -22473 12545 -22456
rect 12345 -22511 12545 -22473
rect 12603 -22473 12686 -22456
rect 12720 -22456 12736 -22439
rect 12928 -22439 12994 -22423
rect 12928 -22456 12944 -22439
rect 12720 -22473 12803 -22456
rect 12603 -22511 12803 -22473
rect 12861 -22473 12944 -22456
rect 12978 -22456 12994 -22439
rect 13186 -22439 13252 -22423
rect 13186 -22456 13202 -22439
rect 12978 -22473 13061 -22456
rect 12861 -22511 13061 -22473
rect 13119 -22473 13202 -22456
rect 13236 -22456 13252 -22439
rect 13444 -22439 13510 -22423
rect 13444 -22456 13460 -22439
rect 13236 -22473 13319 -22456
rect 13119 -22511 13319 -22473
rect 13377 -22473 13460 -22456
rect 13494 -22456 13510 -22439
rect 13702 -22439 13768 -22423
rect 13702 -22456 13718 -22439
rect 13494 -22473 13577 -22456
rect 13377 -22511 13577 -22473
rect 13635 -22473 13718 -22456
rect 13752 -22456 13768 -22439
rect 14559 -22438 14625 -22422
rect 14559 -22455 14575 -22438
rect 13752 -22473 13835 -22456
rect 13635 -22511 13835 -22473
rect 14492 -22472 14575 -22455
rect 14609 -22455 14625 -22438
rect 14817 -22438 14883 -22422
rect 14817 -22455 14833 -22438
rect 14609 -22472 14692 -22455
rect 14492 -22510 14692 -22472
rect 14750 -22472 14833 -22455
rect 14867 -22455 14883 -22438
rect 15075 -22438 15141 -22422
rect 15075 -22455 15091 -22438
rect 14867 -22472 14950 -22455
rect 14750 -22510 14950 -22472
rect 15008 -22472 15091 -22455
rect 15125 -22455 15141 -22438
rect 15333 -22438 15399 -22422
rect 15333 -22455 15349 -22438
rect 15125 -22472 15208 -22455
rect 15008 -22510 15208 -22472
rect 15266 -22472 15349 -22455
rect 15383 -22455 15399 -22438
rect 15591 -22438 15657 -22422
rect 15591 -22455 15607 -22438
rect 15383 -22472 15466 -22455
rect 15266 -22510 15466 -22472
rect 15524 -22472 15607 -22455
rect 15641 -22455 15657 -22438
rect 15849 -22438 15915 -22422
rect 15849 -22455 15865 -22438
rect 15641 -22472 15724 -22455
rect 15524 -22510 15724 -22472
rect 15782 -22472 15865 -22455
rect 15899 -22455 15915 -22438
rect 16107 -22438 16173 -22422
rect 16107 -22455 16123 -22438
rect 15899 -22472 15982 -22455
rect 15782 -22510 15982 -22472
rect 16040 -22472 16123 -22455
rect 16157 -22455 16173 -22438
rect 16365 -22438 16431 -22422
rect 16365 -22455 16381 -22438
rect 16157 -22472 16240 -22455
rect 16040 -22510 16240 -22472
rect 16298 -22472 16381 -22455
rect 16415 -22455 16431 -22438
rect 16415 -22472 16498 -22455
rect 16298 -22510 16498 -22472
rect 9159 -22749 9359 -22711
rect 9159 -22766 9242 -22749
rect 9226 -22783 9242 -22766
rect 9276 -22766 9359 -22749
rect 9417 -22749 9617 -22711
rect 9417 -22766 9500 -22749
rect 9276 -22783 9292 -22766
rect 9226 -22799 9292 -22783
rect 9484 -22783 9500 -22766
rect 9534 -22766 9617 -22749
rect 9675 -22749 9875 -22711
rect 9675 -22766 9758 -22749
rect 9534 -22783 9550 -22766
rect 9484 -22799 9550 -22783
rect 9742 -22783 9758 -22766
rect 9792 -22766 9875 -22749
rect 9933 -22749 10133 -22711
rect 9933 -22766 10016 -22749
rect 9792 -22783 9808 -22766
rect 9742 -22799 9808 -22783
rect 10000 -22783 10016 -22766
rect 10050 -22766 10133 -22749
rect 10191 -22749 10391 -22711
rect 10191 -22766 10274 -22749
rect 10050 -22783 10066 -22766
rect 10000 -22799 10066 -22783
rect 10258 -22783 10274 -22766
rect 10308 -22766 10391 -22749
rect 10449 -22749 10649 -22711
rect 10449 -22766 10532 -22749
rect 10308 -22783 10324 -22766
rect 10258 -22799 10324 -22783
rect 10516 -22783 10532 -22766
rect 10566 -22766 10649 -22749
rect 10707 -22749 10907 -22711
rect 10707 -22766 10790 -22749
rect 10566 -22783 10582 -22766
rect 10516 -22799 10582 -22783
rect 10774 -22783 10790 -22766
rect 10824 -22766 10907 -22749
rect 10965 -22749 11165 -22711
rect 10965 -22766 11048 -22749
rect 10824 -22783 10840 -22766
rect 10774 -22799 10840 -22783
rect 11032 -22783 11048 -22766
rect 11082 -22766 11165 -22749
rect 11829 -22749 12029 -22711
rect 11829 -22766 11912 -22749
rect 11082 -22783 11098 -22766
rect 11032 -22799 11098 -22783
rect 11896 -22783 11912 -22766
rect 11946 -22766 12029 -22749
rect 12087 -22749 12287 -22711
rect 12087 -22766 12170 -22749
rect 11946 -22783 11962 -22766
rect 11896 -22799 11962 -22783
rect 12154 -22783 12170 -22766
rect 12204 -22766 12287 -22749
rect 12345 -22749 12545 -22711
rect 12345 -22766 12428 -22749
rect 12204 -22783 12220 -22766
rect 12154 -22799 12220 -22783
rect 12412 -22783 12428 -22766
rect 12462 -22766 12545 -22749
rect 12603 -22749 12803 -22711
rect 12603 -22766 12686 -22749
rect 12462 -22783 12478 -22766
rect 12412 -22799 12478 -22783
rect 12670 -22783 12686 -22766
rect 12720 -22766 12803 -22749
rect 12861 -22749 13061 -22711
rect 12861 -22766 12944 -22749
rect 12720 -22783 12736 -22766
rect 12670 -22799 12736 -22783
rect 12928 -22783 12944 -22766
rect 12978 -22766 13061 -22749
rect 13119 -22749 13319 -22711
rect 13119 -22766 13202 -22749
rect 12978 -22783 12994 -22766
rect 12928 -22799 12994 -22783
rect 13186 -22783 13202 -22766
rect 13236 -22766 13319 -22749
rect 13377 -22749 13577 -22711
rect 13377 -22766 13460 -22749
rect 13236 -22783 13252 -22766
rect 13186 -22799 13252 -22783
rect 13444 -22783 13460 -22766
rect 13494 -22766 13577 -22749
rect 13635 -22749 13835 -22711
rect 13635 -22766 13718 -22749
rect 13494 -22783 13510 -22766
rect 13444 -22799 13510 -22783
rect 13702 -22783 13718 -22766
rect 13752 -22766 13835 -22749
rect 14492 -22748 14692 -22710
rect 14492 -22765 14575 -22748
rect 13752 -22783 13768 -22766
rect 13702 -22799 13768 -22783
rect 14559 -22782 14575 -22765
rect 14609 -22765 14692 -22748
rect 14750 -22748 14950 -22710
rect 14750 -22765 14833 -22748
rect 14609 -22782 14625 -22765
rect 14559 -22798 14625 -22782
rect 14817 -22782 14833 -22765
rect 14867 -22765 14950 -22748
rect 15008 -22748 15208 -22710
rect 15008 -22765 15091 -22748
rect 14867 -22782 14883 -22765
rect 14817 -22798 14883 -22782
rect 15075 -22782 15091 -22765
rect 15125 -22765 15208 -22748
rect 15266 -22748 15466 -22710
rect 15266 -22765 15349 -22748
rect 15125 -22782 15141 -22765
rect 15075 -22798 15141 -22782
rect 15333 -22782 15349 -22765
rect 15383 -22765 15466 -22748
rect 15524 -22748 15724 -22710
rect 15524 -22765 15607 -22748
rect 15383 -22782 15399 -22765
rect 15333 -22798 15399 -22782
rect 15591 -22782 15607 -22765
rect 15641 -22765 15724 -22748
rect 15782 -22748 15982 -22710
rect 15782 -22765 15865 -22748
rect 15641 -22782 15657 -22765
rect 15591 -22798 15657 -22782
rect 15849 -22782 15865 -22765
rect 15899 -22765 15982 -22748
rect 16040 -22748 16240 -22710
rect 16040 -22765 16123 -22748
rect 15899 -22782 15915 -22765
rect 15849 -22798 15915 -22782
rect 16107 -22782 16123 -22765
rect 16157 -22765 16240 -22748
rect 16298 -22748 16498 -22710
rect 16298 -22765 16381 -22748
rect 16157 -22782 16173 -22765
rect 16107 -22798 16173 -22782
rect 16365 -22782 16381 -22765
rect 16415 -22765 16498 -22748
rect 16415 -22782 16431 -22765
rect 16365 -22798 16431 -22782
rect 9226 -22857 9292 -22841
rect 9226 -22874 9242 -22857
rect 9159 -22891 9242 -22874
rect 9276 -22874 9292 -22857
rect 9484 -22857 9550 -22841
rect 9484 -22874 9500 -22857
rect 9276 -22891 9359 -22874
rect 9159 -22929 9359 -22891
rect 9417 -22891 9500 -22874
rect 9534 -22874 9550 -22857
rect 9742 -22857 9808 -22841
rect 9742 -22874 9758 -22857
rect 9534 -22891 9617 -22874
rect 9417 -22929 9617 -22891
rect 9675 -22891 9758 -22874
rect 9792 -22874 9808 -22857
rect 10000 -22857 10066 -22841
rect 10000 -22874 10016 -22857
rect 9792 -22891 9875 -22874
rect 9675 -22929 9875 -22891
rect 9933 -22891 10016 -22874
rect 10050 -22874 10066 -22857
rect 10258 -22857 10324 -22841
rect 10258 -22874 10274 -22857
rect 10050 -22891 10133 -22874
rect 9933 -22929 10133 -22891
rect 10191 -22891 10274 -22874
rect 10308 -22874 10324 -22857
rect 10516 -22857 10582 -22841
rect 10516 -22874 10532 -22857
rect 10308 -22891 10391 -22874
rect 10191 -22929 10391 -22891
rect 10449 -22891 10532 -22874
rect 10566 -22874 10582 -22857
rect 10774 -22857 10840 -22841
rect 10774 -22874 10790 -22857
rect 10566 -22891 10649 -22874
rect 10449 -22929 10649 -22891
rect 10707 -22891 10790 -22874
rect 10824 -22874 10840 -22857
rect 11032 -22857 11098 -22841
rect 11032 -22874 11048 -22857
rect 10824 -22891 10907 -22874
rect 10707 -22929 10907 -22891
rect 10965 -22891 11048 -22874
rect 11082 -22874 11098 -22857
rect 11896 -22857 11962 -22841
rect 11896 -22874 11912 -22857
rect 11082 -22891 11165 -22874
rect 10965 -22929 11165 -22891
rect 11829 -22891 11912 -22874
rect 11946 -22874 11962 -22857
rect 12154 -22857 12220 -22841
rect 12154 -22874 12170 -22857
rect 11946 -22891 12029 -22874
rect 11829 -22929 12029 -22891
rect 12087 -22891 12170 -22874
rect 12204 -22874 12220 -22857
rect 12412 -22857 12478 -22841
rect 12412 -22874 12428 -22857
rect 12204 -22891 12287 -22874
rect 12087 -22929 12287 -22891
rect 12345 -22891 12428 -22874
rect 12462 -22874 12478 -22857
rect 12670 -22857 12736 -22841
rect 12670 -22874 12686 -22857
rect 12462 -22891 12545 -22874
rect 12345 -22929 12545 -22891
rect 12603 -22891 12686 -22874
rect 12720 -22874 12736 -22857
rect 12928 -22857 12994 -22841
rect 12928 -22874 12944 -22857
rect 12720 -22891 12803 -22874
rect 12603 -22929 12803 -22891
rect 12861 -22891 12944 -22874
rect 12978 -22874 12994 -22857
rect 13186 -22857 13252 -22841
rect 13186 -22874 13202 -22857
rect 12978 -22891 13061 -22874
rect 12861 -22929 13061 -22891
rect 13119 -22891 13202 -22874
rect 13236 -22874 13252 -22857
rect 13444 -22857 13510 -22841
rect 13444 -22874 13460 -22857
rect 13236 -22891 13319 -22874
rect 13119 -22929 13319 -22891
rect 13377 -22891 13460 -22874
rect 13494 -22874 13510 -22857
rect 13702 -22857 13768 -22841
rect 13702 -22874 13718 -22857
rect 13494 -22891 13577 -22874
rect 13377 -22929 13577 -22891
rect 13635 -22891 13718 -22874
rect 13752 -22874 13768 -22857
rect 14559 -22856 14625 -22840
rect 14559 -22873 14575 -22856
rect 13752 -22891 13835 -22874
rect 13635 -22929 13835 -22891
rect 14492 -22890 14575 -22873
rect 14609 -22873 14625 -22856
rect 14817 -22856 14883 -22840
rect 14817 -22873 14833 -22856
rect 14609 -22890 14692 -22873
rect 14492 -22928 14692 -22890
rect 14750 -22890 14833 -22873
rect 14867 -22873 14883 -22856
rect 15075 -22856 15141 -22840
rect 15075 -22873 15091 -22856
rect 14867 -22890 14950 -22873
rect 14750 -22928 14950 -22890
rect 15008 -22890 15091 -22873
rect 15125 -22873 15141 -22856
rect 15333 -22856 15399 -22840
rect 15333 -22873 15349 -22856
rect 15125 -22890 15208 -22873
rect 15008 -22928 15208 -22890
rect 15266 -22890 15349 -22873
rect 15383 -22873 15399 -22856
rect 15591 -22856 15657 -22840
rect 15591 -22873 15607 -22856
rect 15383 -22890 15466 -22873
rect 15266 -22928 15466 -22890
rect 15524 -22890 15607 -22873
rect 15641 -22873 15657 -22856
rect 15849 -22856 15915 -22840
rect 15849 -22873 15865 -22856
rect 15641 -22890 15724 -22873
rect 15524 -22928 15724 -22890
rect 15782 -22890 15865 -22873
rect 15899 -22873 15915 -22856
rect 16107 -22856 16173 -22840
rect 16107 -22873 16123 -22856
rect 15899 -22890 15982 -22873
rect 15782 -22928 15982 -22890
rect 16040 -22890 16123 -22873
rect 16157 -22873 16173 -22856
rect 16365 -22856 16431 -22840
rect 16365 -22873 16381 -22856
rect 16157 -22890 16240 -22873
rect 16040 -22928 16240 -22890
rect 16298 -22890 16381 -22873
rect 16415 -22873 16431 -22856
rect 16415 -22890 16498 -22873
rect 16298 -22928 16498 -22890
rect 9159 -23167 9359 -23129
rect 9159 -23184 9242 -23167
rect 9226 -23201 9242 -23184
rect 9276 -23184 9359 -23167
rect 9417 -23167 9617 -23129
rect 9417 -23184 9500 -23167
rect 9276 -23201 9292 -23184
rect 9226 -23217 9292 -23201
rect 9484 -23201 9500 -23184
rect 9534 -23184 9617 -23167
rect 9675 -23167 9875 -23129
rect 9675 -23184 9758 -23167
rect 9534 -23201 9550 -23184
rect 9484 -23217 9550 -23201
rect 9742 -23201 9758 -23184
rect 9792 -23184 9875 -23167
rect 9933 -23167 10133 -23129
rect 9933 -23184 10016 -23167
rect 9792 -23201 9808 -23184
rect 9742 -23217 9808 -23201
rect 10000 -23201 10016 -23184
rect 10050 -23184 10133 -23167
rect 10191 -23167 10391 -23129
rect 10191 -23184 10274 -23167
rect 10050 -23201 10066 -23184
rect 10000 -23217 10066 -23201
rect 10258 -23201 10274 -23184
rect 10308 -23184 10391 -23167
rect 10449 -23167 10649 -23129
rect 10449 -23184 10532 -23167
rect 10308 -23201 10324 -23184
rect 10258 -23217 10324 -23201
rect 10516 -23201 10532 -23184
rect 10566 -23184 10649 -23167
rect 10707 -23167 10907 -23129
rect 10707 -23184 10790 -23167
rect 10566 -23201 10582 -23184
rect 10516 -23217 10582 -23201
rect 10774 -23201 10790 -23184
rect 10824 -23184 10907 -23167
rect 10965 -23167 11165 -23129
rect 10965 -23184 11048 -23167
rect 10824 -23201 10840 -23184
rect 10774 -23217 10840 -23201
rect 11032 -23201 11048 -23184
rect 11082 -23184 11165 -23167
rect 11829 -23167 12029 -23129
rect 11829 -23184 11912 -23167
rect 11082 -23201 11098 -23184
rect 11032 -23217 11098 -23201
rect 11896 -23201 11912 -23184
rect 11946 -23184 12029 -23167
rect 12087 -23167 12287 -23129
rect 12087 -23184 12170 -23167
rect 11946 -23201 11962 -23184
rect 11896 -23217 11962 -23201
rect 12154 -23201 12170 -23184
rect 12204 -23184 12287 -23167
rect 12345 -23167 12545 -23129
rect 12345 -23184 12428 -23167
rect 12204 -23201 12220 -23184
rect 12154 -23217 12220 -23201
rect 12412 -23201 12428 -23184
rect 12462 -23184 12545 -23167
rect 12603 -23167 12803 -23129
rect 12603 -23184 12686 -23167
rect 12462 -23201 12478 -23184
rect 12412 -23217 12478 -23201
rect 12670 -23201 12686 -23184
rect 12720 -23184 12803 -23167
rect 12861 -23167 13061 -23129
rect 12861 -23184 12944 -23167
rect 12720 -23201 12736 -23184
rect 12670 -23217 12736 -23201
rect 12928 -23201 12944 -23184
rect 12978 -23184 13061 -23167
rect 13119 -23167 13319 -23129
rect 13119 -23184 13202 -23167
rect 12978 -23201 12994 -23184
rect 12928 -23217 12994 -23201
rect 13186 -23201 13202 -23184
rect 13236 -23184 13319 -23167
rect 13377 -23167 13577 -23129
rect 13377 -23184 13460 -23167
rect 13236 -23201 13252 -23184
rect 13186 -23217 13252 -23201
rect 13444 -23201 13460 -23184
rect 13494 -23184 13577 -23167
rect 13635 -23167 13835 -23129
rect 13635 -23184 13718 -23167
rect 13494 -23201 13510 -23184
rect 13444 -23217 13510 -23201
rect 13702 -23201 13718 -23184
rect 13752 -23184 13835 -23167
rect 14492 -23166 14692 -23128
rect 14492 -23183 14575 -23166
rect 13752 -23201 13768 -23184
rect 13702 -23217 13768 -23201
rect 14559 -23200 14575 -23183
rect 14609 -23183 14692 -23166
rect 14750 -23166 14950 -23128
rect 14750 -23183 14833 -23166
rect 14609 -23200 14625 -23183
rect 14559 -23216 14625 -23200
rect 14817 -23200 14833 -23183
rect 14867 -23183 14950 -23166
rect 15008 -23166 15208 -23128
rect 15008 -23183 15091 -23166
rect 14867 -23200 14883 -23183
rect 14817 -23216 14883 -23200
rect 15075 -23200 15091 -23183
rect 15125 -23183 15208 -23166
rect 15266 -23166 15466 -23128
rect 15266 -23183 15349 -23166
rect 15125 -23200 15141 -23183
rect 15075 -23216 15141 -23200
rect 15333 -23200 15349 -23183
rect 15383 -23183 15466 -23166
rect 15524 -23166 15724 -23128
rect 15524 -23183 15607 -23166
rect 15383 -23200 15399 -23183
rect 15333 -23216 15399 -23200
rect 15591 -23200 15607 -23183
rect 15641 -23183 15724 -23166
rect 15782 -23166 15982 -23128
rect 15782 -23183 15865 -23166
rect 15641 -23200 15657 -23183
rect 15591 -23216 15657 -23200
rect 15849 -23200 15865 -23183
rect 15899 -23183 15982 -23166
rect 16040 -23166 16240 -23128
rect 16040 -23183 16123 -23166
rect 15899 -23200 15915 -23183
rect 15849 -23216 15915 -23200
rect 16107 -23200 16123 -23183
rect 16157 -23183 16240 -23166
rect 16298 -23166 16498 -23128
rect 16298 -23183 16381 -23166
rect 16157 -23200 16173 -23183
rect 16107 -23216 16173 -23200
rect 16365 -23200 16381 -23183
rect 16415 -23183 16498 -23166
rect 16415 -23200 16431 -23183
rect 16365 -23216 16431 -23200
rect 9226 -23275 9292 -23259
rect 9226 -23292 9242 -23275
rect 9159 -23309 9242 -23292
rect 9276 -23292 9292 -23275
rect 9484 -23275 9550 -23259
rect 9484 -23292 9500 -23275
rect 9276 -23309 9359 -23292
rect 9159 -23347 9359 -23309
rect 9417 -23309 9500 -23292
rect 9534 -23292 9550 -23275
rect 9742 -23275 9808 -23259
rect 9742 -23292 9758 -23275
rect 9534 -23309 9617 -23292
rect 9417 -23347 9617 -23309
rect 9675 -23309 9758 -23292
rect 9792 -23292 9808 -23275
rect 10000 -23275 10066 -23259
rect 10000 -23292 10016 -23275
rect 9792 -23309 9875 -23292
rect 9675 -23347 9875 -23309
rect 9933 -23309 10016 -23292
rect 10050 -23292 10066 -23275
rect 10258 -23275 10324 -23259
rect 10258 -23292 10274 -23275
rect 10050 -23309 10133 -23292
rect 9933 -23347 10133 -23309
rect 10191 -23309 10274 -23292
rect 10308 -23292 10324 -23275
rect 10516 -23275 10582 -23259
rect 10516 -23292 10532 -23275
rect 10308 -23309 10391 -23292
rect 10191 -23347 10391 -23309
rect 10449 -23309 10532 -23292
rect 10566 -23292 10582 -23275
rect 10774 -23275 10840 -23259
rect 10774 -23292 10790 -23275
rect 10566 -23309 10649 -23292
rect 10449 -23347 10649 -23309
rect 10707 -23309 10790 -23292
rect 10824 -23292 10840 -23275
rect 11032 -23275 11098 -23259
rect 11032 -23292 11048 -23275
rect 10824 -23309 10907 -23292
rect 10707 -23347 10907 -23309
rect 10965 -23309 11048 -23292
rect 11082 -23292 11098 -23275
rect 11896 -23275 11962 -23259
rect 11896 -23292 11912 -23275
rect 11082 -23309 11165 -23292
rect 10965 -23347 11165 -23309
rect 11829 -23309 11912 -23292
rect 11946 -23292 11962 -23275
rect 12154 -23275 12220 -23259
rect 12154 -23292 12170 -23275
rect 11946 -23309 12029 -23292
rect 11829 -23347 12029 -23309
rect 12087 -23309 12170 -23292
rect 12204 -23292 12220 -23275
rect 12412 -23275 12478 -23259
rect 12412 -23292 12428 -23275
rect 12204 -23309 12287 -23292
rect 12087 -23347 12287 -23309
rect 12345 -23309 12428 -23292
rect 12462 -23292 12478 -23275
rect 12670 -23275 12736 -23259
rect 12670 -23292 12686 -23275
rect 12462 -23309 12545 -23292
rect 12345 -23347 12545 -23309
rect 12603 -23309 12686 -23292
rect 12720 -23292 12736 -23275
rect 12928 -23275 12994 -23259
rect 12928 -23292 12944 -23275
rect 12720 -23309 12803 -23292
rect 12603 -23347 12803 -23309
rect 12861 -23309 12944 -23292
rect 12978 -23292 12994 -23275
rect 13186 -23275 13252 -23259
rect 13186 -23292 13202 -23275
rect 12978 -23309 13061 -23292
rect 12861 -23347 13061 -23309
rect 13119 -23309 13202 -23292
rect 13236 -23292 13252 -23275
rect 13444 -23275 13510 -23259
rect 13444 -23292 13460 -23275
rect 13236 -23309 13319 -23292
rect 13119 -23347 13319 -23309
rect 13377 -23309 13460 -23292
rect 13494 -23292 13510 -23275
rect 13702 -23275 13768 -23259
rect 13702 -23292 13718 -23275
rect 13494 -23309 13577 -23292
rect 13377 -23347 13577 -23309
rect 13635 -23309 13718 -23292
rect 13752 -23292 13768 -23275
rect 14559 -23274 14625 -23258
rect 14559 -23291 14575 -23274
rect 13752 -23309 13835 -23292
rect 13635 -23347 13835 -23309
rect 14492 -23308 14575 -23291
rect 14609 -23291 14625 -23274
rect 14817 -23274 14883 -23258
rect 14817 -23291 14833 -23274
rect 14609 -23308 14692 -23291
rect 14492 -23346 14692 -23308
rect 14750 -23308 14833 -23291
rect 14867 -23291 14883 -23274
rect 15075 -23274 15141 -23258
rect 15075 -23291 15091 -23274
rect 14867 -23308 14950 -23291
rect 14750 -23346 14950 -23308
rect 15008 -23308 15091 -23291
rect 15125 -23291 15141 -23274
rect 15333 -23274 15399 -23258
rect 15333 -23291 15349 -23274
rect 15125 -23308 15208 -23291
rect 15008 -23346 15208 -23308
rect 15266 -23308 15349 -23291
rect 15383 -23291 15399 -23274
rect 15591 -23274 15657 -23258
rect 15591 -23291 15607 -23274
rect 15383 -23308 15466 -23291
rect 15266 -23346 15466 -23308
rect 15524 -23308 15607 -23291
rect 15641 -23291 15657 -23274
rect 15849 -23274 15915 -23258
rect 15849 -23291 15865 -23274
rect 15641 -23308 15724 -23291
rect 15524 -23346 15724 -23308
rect 15782 -23308 15865 -23291
rect 15899 -23291 15915 -23274
rect 16107 -23274 16173 -23258
rect 16107 -23291 16123 -23274
rect 15899 -23308 15982 -23291
rect 15782 -23346 15982 -23308
rect 16040 -23308 16123 -23291
rect 16157 -23291 16173 -23274
rect 16365 -23274 16431 -23258
rect 16365 -23291 16381 -23274
rect 16157 -23308 16240 -23291
rect 16040 -23346 16240 -23308
rect 16298 -23308 16381 -23291
rect 16415 -23291 16431 -23274
rect 16415 -23308 16498 -23291
rect 16298 -23346 16498 -23308
rect 9159 -23585 9359 -23547
rect 9159 -23602 9242 -23585
rect 9226 -23619 9242 -23602
rect 9276 -23602 9359 -23585
rect 9417 -23585 9617 -23547
rect 9417 -23602 9500 -23585
rect 9276 -23619 9292 -23602
rect 9226 -23635 9292 -23619
rect 9484 -23619 9500 -23602
rect 9534 -23602 9617 -23585
rect 9675 -23585 9875 -23547
rect 9675 -23602 9758 -23585
rect 9534 -23619 9550 -23602
rect 9484 -23635 9550 -23619
rect 9742 -23619 9758 -23602
rect 9792 -23602 9875 -23585
rect 9933 -23585 10133 -23547
rect 9933 -23602 10016 -23585
rect 9792 -23619 9808 -23602
rect 9742 -23635 9808 -23619
rect 10000 -23619 10016 -23602
rect 10050 -23602 10133 -23585
rect 10191 -23585 10391 -23547
rect 10191 -23602 10274 -23585
rect 10050 -23619 10066 -23602
rect 10000 -23635 10066 -23619
rect 10258 -23619 10274 -23602
rect 10308 -23602 10391 -23585
rect 10449 -23585 10649 -23547
rect 10449 -23602 10532 -23585
rect 10308 -23619 10324 -23602
rect 10258 -23635 10324 -23619
rect 10516 -23619 10532 -23602
rect 10566 -23602 10649 -23585
rect 10707 -23585 10907 -23547
rect 10707 -23602 10790 -23585
rect 10566 -23619 10582 -23602
rect 10516 -23635 10582 -23619
rect 10774 -23619 10790 -23602
rect 10824 -23602 10907 -23585
rect 10965 -23585 11165 -23547
rect 10965 -23602 11048 -23585
rect 10824 -23619 10840 -23602
rect 10774 -23635 10840 -23619
rect 11032 -23619 11048 -23602
rect 11082 -23602 11165 -23585
rect 11829 -23585 12029 -23547
rect 11829 -23602 11912 -23585
rect 11082 -23619 11098 -23602
rect 11032 -23635 11098 -23619
rect 11896 -23619 11912 -23602
rect 11946 -23602 12029 -23585
rect 12087 -23585 12287 -23547
rect 12087 -23602 12170 -23585
rect 11946 -23619 11962 -23602
rect 11896 -23635 11962 -23619
rect 12154 -23619 12170 -23602
rect 12204 -23602 12287 -23585
rect 12345 -23585 12545 -23547
rect 12345 -23602 12428 -23585
rect 12204 -23619 12220 -23602
rect 12154 -23635 12220 -23619
rect 12412 -23619 12428 -23602
rect 12462 -23602 12545 -23585
rect 12603 -23585 12803 -23547
rect 12603 -23602 12686 -23585
rect 12462 -23619 12478 -23602
rect 12412 -23635 12478 -23619
rect 12670 -23619 12686 -23602
rect 12720 -23602 12803 -23585
rect 12861 -23585 13061 -23547
rect 12861 -23602 12944 -23585
rect 12720 -23619 12736 -23602
rect 12670 -23635 12736 -23619
rect 12928 -23619 12944 -23602
rect 12978 -23602 13061 -23585
rect 13119 -23585 13319 -23547
rect 13119 -23602 13202 -23585
rect 12978 -23619 12994 -23602
rect 12928 -23635 12994 -23619
rect 13186 -23619 13202 -23602
rect 13236 -23602 13319 -23585
rect 13377 -23585 13577 -23547
rect 13377 -23602 13460 -23585
rect 13236 -23619 13252 -23602
rect 13186 -23635 13252 -23619
rect 13444 -23619 13460 -23602
rect 13494 -23602 13577 -23585
rect 13635 -23585 13835 -23547
rect 13635 -23602 13718 -23585
rect 13494 -23619 13510 -23602
rect 13444 -23635 13510 -23619
rect 13702 -23619 13718 -23602
rect 13752 -23602 13835 -23585
rect 14492 -23584 14692 -23546
rect 14492 -23601 14575 -23584
rect 13752 -23619 13768 -23602
rect 13702 -23635 13768 -23619
rect 14559 -23618 14575 -23601
rect 14609 -23601 14692 -23584
rect 14750 -23584 14950 -23546
rect 14750 -23601 14833 -23584
rect 14609 -23618 14625 -23601
rect 14559 -23634 14625 -23618
rect 14817 -23618 14833 -23601
rect 14867 -23601 14950 -23584
rect 15008 -23584 15208 -23546
rect 15008 -23601 15091 -23584
rect 14867 -23618 14883 -23601
rect 14817 -23634 14883 -23618
rect 15075 -23618 15091 -23601
rect 15125 -23601 15208 -23584
rect 15266 -23584 15466 -23546
rect 15266 -23601 15349 -23584
rect 15125 -23618 15141 -23601
rect 15075 -23634 15141 -23618
rect 15333 -23618 15349 -23601
rect 15383 -23601 15466 -23584
rect 15524 -23584 15724 -23546
rect 15524 -23601 15607 -23584
rect 15383 -23618 15399 -23601
rect 15333 -23634 15399 -23618
rect 15591 -23618 15607 -23601
rect 15641 -23601 15724 -23584
rect 15782 -23584 15982 -23546
rect 15782 -23601 15865 -23584
rect 15641 -23618 15657 -23601
rect 15591 -23634 15657 -23618
rect 15849 -23618 15865 -23601
rect 15899 -23601 15982 -23584
rect 16040 -23584 16240 -23546
rect 16040 -23601 16123 -23584
rect 15899 -23618 15915 -23601
rect 15849 -23634 15915 -23618
rect 16107 -23618 16123 -23601
rect 16157 -23601 16240 -23584
rect 16298 -23584 16498 -23546
rect 16298 -23601 16381 -23584
rect 16157 -23618 16173 -23601
rect 16107 -23634 16173 -23618
rect 16365 -23618 16381 -23601
rect 16415 -23601 16498 -23584
rect 16415 -23618 16431 -23601
rect 16365 -23634 16431 -23618
rect 9226 -23693 9292 -23677
rect 9226 -23710 9242 -23693
rect 9159 -23727 9242 -23710
rect 9276 -23710 9292 -23693
rect 9484 -23693 9550 -23677
rect 9484 -23710 9500 -23693
rect 9276 -23727 9359 -23710
rect 9159 -23765 9359 -23727
rect 9417 -23727 9500 -23710
rect 9534 -23710 9550 -23693
rect 9742 -23693 9808 -23677
rect 9742 -23710 9758 -23693
rect 9534 -23727 9617 -23710
rect 9417 -23765 9617 -23727
rect 9675 -23727 9758 -23710
rect 9792 -23710 9808 -23693
rect 10000 -23693 10066 -23677
rect 10000 -23710 10016 -23693
rect 9792 -23727 9875 -23710
rect 9675 -23765 9875 -23727
rect 9933 -23727 10016 -23710
rect 10050 -23710 10066 -23693
rect 10258 -23693 10324 -23677
rect 10258 -23710 10274 -23693
rect 10050 -23727 10133 -23710
rect 9933 -23765 10133 -23727
rect 10191 -23727 10274 -23710
rect 10308 -23710 10324 -23693
rect 10516 -23693 10582 -23677
rect 10516 -23710 10532 -23693
rect 10308 -23727 10391 -23710
rect 10191 -23765 10391 -23727
rect 10449 -23727 10532 -23710
rect 10566 -23710 10582 -23693
rect 10774 -23693 10840 -23677
rect 10774 -23710 10790 -23693
rect 10566 -23727 10649 -23710
rect 10449 -23765 10649 -23727
rect 10707 -23727 10790 -23710
rect 10824 -23710 10840 -23693
rect 11032 -23693 11098 -23677
rect 11032 -23710 11048 -23693
rect 10824 -23727 10907 -23710
rect 10707 -23765 10907 -23727
rect 10965 -23727 11048 -23710
rect 11082 -23710 11098 -23693
rect 11896 -23693 11962 -23677
rect 11896 -23710 11912 -23693
rect 11082 -23727 11165 -23710
rect 10965 -23765 11165 -23727
rect 11829 -23727 11912 -23710
rect 11946 -23710 11962 -23693
rect 12154 -23693 12220 -23677
rect 12154 -23710 12170 -23693
rect 11946 -23727 12029 -23710
rect 11829 -23765 12029 -23727
rect 12087 -23727 12170 -23710
rect 12204 -23710 12220 -23693
rect 12412 -23693 12478 -23677
rect 12412 -23710 12428 -23693
rect 12204 -23727 12287 -23710
rect 12087 -23765 12287 -23727
rect 12345 -23727 12428 -23710
rect 12462 -23710 12478 -23693
rect 12670 -23693 12736 -23677
rect 12670 -23710 12686 -23693
rect 12462 -23727 12545 -23710
rect 12345 -23765 12545 -23727
rect 12603 -23727 12686 -23710
rect 12720 -23710 12736 -23693
rect 12928 -23693 12994 -23677
rect 12928 -23710 12944 -23693
rect 12720 -23727 12803 -23710
rect 12603 -23765 12803 -23727
rect 12861 -23727 12944 -23710
rect 12978 -23710 12994 -23693
rect 13186 -23693 13252 -23677
rect 13186 -23710 13202 -23693
rect 12978 -23727 13061 -23710
rect 12861 -23765 13061 -23727
rect 13119 -23727 13202 -23710
rect 13236 -23710 13252 -23693
rect 13444 -23693 13510 -23677
rect 13444 -23710 13460 -23693
rect 13236 -23727 13319 -23710
rect 13119 -23765 13319 -23727
rect 13377 -23727 13460 -23710
rect 13494 -23710 13510 -23693
rect 13702 -23693 13768 -23677
rect 13702 -23710 13718 -23693
rect 13494 -23727 13577 -23710
rect 13377 -23765 13577 -23727
rect 13635 -23727 13718 -23710
rect 13752 -23710 13768 -23693
rect 14559 -23692 14625 -23676
rect 14559 -23709 14575 -23692
rect 13752 -23727 13835 -23710
rect 13635 -23765 13835 -23727
rect 14492 -23726 14575 -23709
rect 14609 -23709 14625 -23692
rect 14817 -23692 14883 -23676
rect 14817 -23709 14833 -23692
rect 14609 -23726 14692 -23709
rect 14492 -23764 14692 -23726
rect 14750 -23726 14833 -23709
rect 14867 -23709 14883 -23692
rect 15075 -23692 15141 -23676
rect 15075 -23709 15091 -23692
rect 14867 -23726 14950 -23709
rect 14750 -23764 14950 -23726
rect 15008 -23726 15091 -23709
rect 15125 -23709 15141 -23692
rect 15333 -23692 15399 -23676
rect 15333 -23709 15349 -23692
rect 15125 -23726 15208 -23709
rect 15008 -23764 15208 -23726
rect 15266 -23726 15349 -23709
rect 15383 -23709 15399 -23692
rect 15591 -23692 15657 -23676
rect 15591 -23709 15607 -23692
rect 15383 -23726 15466 -23709
rect 15266 -23764 15466 -23726
rect 15524 -23726 15607 -23709
rect 15641 -23709 15657 -23692
rect 15849 -23692 15915 -23676
rect 15849 -23709 15865 -23692
rect 15641 -23726 15724 -23709
rect 15524 -23764 15724 -23726
rect 15782 -23726 15865 -23709
rect 15899 -23709 15915 -23692
rect 16107 -23692 16173 -23676
rect 16107 -23709 16123 -23692
rect 15899 -23726 15982 -23709
rect 15782 -23764 15982 -23726
rect 16040 -23726 16123 -23709
rect 16157 -23709 16173 -23692
rect 16365 -23692 16431 -23676
rect 16365 -23709 16381 -23692
rect 16157 -23726 16240 -23709
rect 16040 -23764 16240 -23726
rect 16298 -23726 16381 -23709
rect 16415 -23709 16431 -23692
rect 16415 -23726 16498 -23709
rect 16298 -23764 16498 -23726
rect 9159 -24003 9359 -23965
rect 9159 -24020 9242 -24003
rect 9226 -24037 9242 -24020
rect 9276 -24020 9359 -24003
rect 9417 -24003 9617 -23965
rect 9417 -24020 9500 -24003
rect 9276 -24037 9292 -24020
rect 9226 -24053 9292 -24037
rect 9484 -24037 9500 -24020
rect 9534 -24020 9617 -24003
rect 9675 -24003 9875 -23965
rect 9675 -24020 9758 -24003
rect 9534 -24037 9550 -24020
rect 9484 -24053 9550 -24037
rect 9742 -24037 9758 -24020
rect 9792 -24020 9875 -24003
rect 9933 -24003 10133 -23965
rect 9933 -24020 10016 -24003
rect 9792 -24037 9808 -24020
rect 9742 -24053 9808 -24037
rect 10000 -24037 10016 -24020
rect 10050 -24020 10133 -24003
rect 10191 -24003 10391 -23965
rect 10191 -24020 10274 -24003
rect 10050 -24037 10066 -24020
rect 10000 -24053 10066 -24037
rect 10258 -24037 10274 -24020
rect 10308 -24020 10391 -24003
rect 10449 -24003 10649 -23965
rect 10449 -24020 10532 -24003
rect 10308 -24037 10324 -24020
rect 10258 -24053 10324 -24037
rect 10516 -24037 10532 -24020
rect 10566 -24020 10649 -24003
rect 10707 -24003 10907 -23965
rect 10707 -24020 10790 -24003
rect 10566 -24037 10582 -24020
rect 10516 -24053 10582 -24037
rect 10774 -24037 10790 -24020
rect 10824 -24020 10907 -24003
rect 10965 -24003 11165 -23965
rect 10965 -24020 11048 -24003
rect 10824 -24037 10840 -24020
rect 10774 -24053 10840 -24037
rect 11032 -24037 11048 -24020
rect 11082 -24020 11165 -24003
rect 11829 -24003 12029 -23965
rect 11829 -24020 11912 -24003
rect 11082 -24037 11098 -24020
rect 11032 -24053 11098 -24037
rect 11896 -24037 11912 -24020
rect 11946 -24020 12029 -24003
rect 12087 -24003 12287 -23965
rect 12087 -24020 12170 -24003
rect 11946 -24037 11962 -24020
rect 11896 -24053 11962 -24037
rect 12154 -24037 12170 -24020
rect 12204 -24020 12287 -24003
rect 12345 -24003 12545 -23965
rect 12345 -24020 12428 -24003
rect 12204 -24037 12220 -24020
rect 12154 -24053 12220 -24037
rect 12412 -24037 12428 -24020
rect 12462 -24020 12545 -24003
rect 12603 -24003 12803 -23965
rect 12603 -24020 12686 -24003
rect 12462 -24037 12478 -24020
rect 12412 -24053 12478 -24037
rect 12670 -24037 12686 -24020
rect 12720 -24020 12803 -24003
rect 12861 -24003 13061 -23965
rect 12861 -24020 12944 -24003
rect 12720 -24037 12736 -24020
rect 12670 -24053 12736 -24037
rect 12928 -24037 12944 -24020
rect 12978 -24020 13061 -24003
rect 13119 -24003 13319 -23965
rect 13119 -24020 13202 -24003
rect 12978 -24037 12994 -24020
rect 12928 -24053 12994 -24037
rect 13186 -24037 13202 -24020
rect 13236 -24020 13319 -24003
rect 13377 -24003 13577 -23965
rect 13377 -24020 13460 -24003
rect 13236 -24037 13252 -24020
rect 13186 -24053 13252 -24037
rect 13444 -24037 13460 -24020
rect 13494 -24020 13577 -24003
rect 13635 -24003 13835 -23965
rect 13635 -24020 13718 -24003
rect 13494 -24037 13510 -24020
rect 13444 -24053 13510 -24037
rect 13702 -24037 13718 -24020
rect 13752 -24020 13835 -24003
rect 14492 -24002 14692 -23964
rect 14492 -24019 14575 -24002
rect 13752 -24037 13768 -24020
rect 13702 -24053 13768 -24037
rect 14559 -24036 14575 -24019
rect 14609 -24019 14692 -24002
rect 14750 -24002 14950 -23964
rect 14750 -24019 14833 -24002
rect 14609 -24036 14625 -24019
rect 14559 -24052 14625 -24036
rect 14817 -24036 14833 -24019
rect 14867 -24019 14950 -24002
rect 15008 -24002 15208 -23964
rect 15008 -24019 15091 -24002
rect 14867 -24036 14883 -24019
rect 14817 -24052 14883 -24036
rect 15075 -24036 15091 -24019
rect 15125 -24019 15208 -24002
rect 15266 -24002 15466 -23964
rect 15266 -24019 15349 -24002
rect 15125 -24036 15141 -24019
rect 15075 -24052 15141 -24036
rect 15333 -24036 15349 -24019
rect 15383 -24019 15466 -24002
rect 15524 -24002 15724 -23964
rect 15524 -24019 15607 -24002
rect 15383 -24036 15399 -24019
rect 15333 -24052 15399 -24036
rect 15591 -24036 15607 -24019
rect 15641 -24019 15724 -24002
rect 15782 -24002 15982 -23964
rect 15782 -24019 15865 -24002
rect 15641 -24036 15657 -24019
rect 15591 -24052 15657 -24036
rect 15849 -24036 15865 -24019
rect 15899 -24019 15982 -24002
rect 16040 -24002 16240 -23964
rect 16040 -24019 16123 -24002
rect 15899 -24036 15915 -24019
rect 15849 -24052 15915 -24036
rect 16107 -24036 16123 -24019
rect 16157 -24019 16240 -24002
rect 16298 -24002 16498 -23964
rect 16298 -24019 16381 -24002
rect 16157 -24036 16173 -24019
rect 16107 -24052 16173 -24036
rect 16365 -24036 16381 -24019
rect 16415 -24019 16498 -24002
rect 16415 -24036 16431 -24019
rect 16365 -24052 16431 -24036
rect 9106 -24345 9172 -24329
rect 9106 -24362 9122 -24345
rect 9039 -24379 9122 -24362
rect 9156 -24362 9172 -24345
rect 9646 -24345 9712 -24329
rect 9646 -24362 9662 -24345
rect 9156 -24379 9239 -24362
rect 9039 -24417 9239 -24379
rect 9579 -24379 9662 -24362
rect 9696 -24362 9712 -24345
rect 10126 -24345 10192 -24329
rect 10126 -24362 10142 -24345
rect 9696 -24379 9779 -24362
rect 9579 -24417 9779 -24379
rect 10059 -24379 10142 -24362
rect 10176 -24362 10192 -24345
rect 10629 -24343 10695 -24327
rect 10629 -24360 10645 -24343
rect 10176 -24379 10259 -24362
rect 10059 -24417 10259 -24379
rect 10562 -24377 10645 -24360
rect 10679 -24360 10695 -24343
rect 11139 -24333 11205 -24317
rect 11139 -24350 11155 -24333
rect 10679 -24377 10762 -24360
rect 10562 -24415 10762 -24377
rect 11072 -24367 11155 -24350
rect 11189 -24350 11205 -24333
rect 11776 -24345 11842 -24329
rect 11189 -24367 11272 -24350
rect 11776 -24362 11792 -24345
rect 11072 -24405 11272 -24367
rect 11709 -24379 11792 -24362
rect 11826 -24362 11842 -24345
rect 12316 -24345 12382 -24329
rect 12316 -24362 12332 -24345
rect 11826 -24379 11909 -24362
rect 11709 -24417 11909 -24379
rect 12249 -24379 12332 -24362
rect 12366 -24362 12382 -24345
rect 12796 -24345 12862 -24329
rect 12796 -24362 12812 -24345
rect 12366 -24379 12449 -24362
rect 12249 -24417 12449 -24379
rect 12729 -24379 12812 -24362
rect 12846 -24362 12862 -24345
rect 13299 -24343 13365 -24327
rect 13299 -24360 13315 -24343
rect 12846 -24379 12929 -24362
rect 12729 -24417 12929 -24379
rect 13232 -24377 13315 -24360
rect 13349 -24360 13365 -24343
rect 13809 -24333 13875 -24317
rect 13809 -24350 13825 -24333
rect 13349 -24377 13432 -24360
rect 13232 -24415 13432 -24377
rect 13742 -24367 13825 -24350
rect 13859 -24350 13875 -24333
rect 14439 -24344 14505 -24328
rect 13859 -24367 13942 -24350
rect 14439 -24361 14455 -24344
rect 13742 -24405 13942 -24367
rect 14372 -24378 14455 -24361
rect 14489 -24361 14505 -24344
rect 14979 -24344 15045 -24328
rect 14979 -24361 14995 -24344
rect 14489 -24378 14572 -24361
rect 9039 -24655 9239 -24617
rect 9039 -24672 9122 -24655
rect 9106 -24689 9122 -24672
rect 9156 -24672 9239 -24655
rect 9579 -24655 9779 -24617
rect 9579 -24672 9662 -24655
rect 9156 -24689 9172 -24672
rect 9106 -24705 9172 -24689
rect 9646 -24689 9662 -24672
rect 9696 -24672 9779 -24655
rect 10059 -24655 10259 -24617
rect 10059 -24672 10142 -24655
rect 9696 -24689 9712 -24672
rect 9646 -24705 9712 -24689
rect 10126 -24689 10142 -24672
rect 10176 -24672 10259 -24655
rect 10562 -24653 10762 -24615
rect 10562 -24670 10645 -24653
rect 10176 -24689 10192 -24672
rect 10126 -24705 10192 -24689
rect 10629 -24687 10645 -24670
rect 10679 -24670 10762 -24653
rect 11072 -24643 11272 -24605
rect 14372 -24416 14572 -24378
rect 14912 -24378 14995 -24361
rect 15029 -24361 15045 -24344
rect 15459 -24344 15525 -24328
rect 15459 -24361 15475 -24344
rect 15029 -24378 15112 -24361
rect 14912 -24416 15112 -24378
rect 15392 -24378 15475 -24361
rect 15509 -24361 15525 -24344
rect 15962 -24342 16028 -24326
rect 15962 -24359 15978 -24342
rect 15509 -24378 15592 -24361
rect 15392 -24416 15592 -24378
rect 15895 -24376 15978 -24359
rect 16012 -24359 16028 -24342
rect 16472 -24332 16538 -24316
rect 16472 -24349 16488 -24332
rect 16012 -24376 16095 -24359
rect 15895 -24414 16095 -24376
rect 16405 -24366 16488 -24349
rect 16522 -24349 16538 -24332
rect 16522 -24366 16605 -24349
rect 16405 -24404 16605 -24366
rect 11072 -24660 11155 -24643
rect 10679 -24687 10695 -24670
rect 10629 -24703 10695 -24687
rect 11139 -24677 11155 -24660
rect 11189 -24660 11272 -24643
rect 11709 -24655 11909 -24617
rect 11189 -24677 11205 -24660
rect 11709 -24672 11792 -24655
rect 11139 -24693 11205 -24677
rect 11776 -24689 11792 -24672
rect 11826 -24672 11909 -24655
rect 12249 -24655 12449 -24617
rect 12249 -24672 12332 -24655
rect 11826 -24689 11842 -24672
rect 11776 -24705 11842 -24689
rect 12316 -24689 12332 -24672
rect 12366 -24672 12449 -24655
rect 12729 -24655 12929 -24617
rect 12729 -24672 12812 -24655
rect 12366 -24689 12382 -24672
rect 12316 -24705 12382 -24689
rect 12796 -24689 12812 -24672
rect 12846 -24672 12929 -24655
rect 13232 -24653 13432 -24615
rect 13232 -24670 13315 -24653
rect 12846 -24689 12862 -24672
rect 12796 -24705 12862 -24689
rect 13299 -24687 13315 -24670
rect 13349 -24670 13432 -24653
rect 13742 -24643 13942 -24605
rect 13742 -24660 13825 -24643
rect 13349 -24687 13365 -24670
rect 13299 -24703 13365 -24687
rect 13809 -24677 13825 -24660
rect 13859 -24660 13942 -24643
rect 14372 -24654 14572 -24616
rect 13859 -24677 13875 -24660
rect 14372 -24671 14455 -24654
rect 13809 -24693 13875 -24677
rect 14439 -24688 14455 -24671
rect 14489 -24671 14572 -24654
rect 14912 -24654 15112 -24616
rect 14912 -24671 14995 -24654
rect 14489 -24688 14505 -24671
rect 14439 -24704 14505 -24688
rect 14979 -24688 14995 -24671
rect 15029 -24671 15112 -24654
rect 15392 -24654 15592 -24616
rect 15392 -24671 15475 -24654
rect 15029 -24688 15045 -24671
rect 14979 -24704 15045 -24688
rect 15459 -24688 15475 -24671
rect 15509 -24671 15592 -24654
rect 15895 -24652 16095 -24614
rect 15895 -24669 15978 -24652
rect 15509 -24688 15525 -24671
rect 15459 -24704 15525 -24688
rect 15962 -24686 15978 -24669
rect 16012 -24669 16095 -24652
rect 16405 -24642 16605 -24604
rect 16405 -24659 16488 -24642
rect 16012 -24686 16028 -24669
rect 15962 -24702 16028 -24686
rect 16472 -24676 16488 -24659
rect 16522 -24659 16605 -24642
rect 16522 -24676 16538 -24659
rect 16472 -24692 16538 -24676
rect 18036 -7550 19636 -7534
rect 18036 -7584 18052 -7550
rect 19420 -7584 19636 -7550
rect 18036 -7622 19636 -7584
rect 19694 -7550 21294 -7534
rect 19694 -7584 19913 -7550
rect 21278 -7584 21294 -7550
rect 19694 -7622 21294 -7584
rect 18036 -9060 19636 -9022
rect 18036 -9094 18052 -9060
rect 19420 -9094 19636 -9060
rect 18036 -9132 19636 -9094
rect 19694 -9060 21294 -9022
rect 19694 -9094 19913 -9060
rect 21278 -9094 21294 -9060
rect 19694 -9132 21294 -9094
rect 18036 -10570 19636 -10532
rect 18036 -10604 18052 -10570
rect 19420 -10604 19636 -10570
rect 18036 -10642 19636 -10604
rect 19694 -10570 21294 -10532
rect 19694 -10604 19913 -10570
rect 21278 -10604 21294 -10570
rect 19694 -10642 21294 -10604
rect 18036 -12080 19636 -12042
rect 18036 -12114 18052 -12080
rect 19420 -12114 19636 -12080
rect 18036 -12152 19636 -12114
rect 19694 -12080 21294 -12042
rect 19694 -12114 19913 -12080
rect 21278 -12114 21294 -12080
rect 19694 -12152 21294 -12114
rect 18036 -13590 19636 -13552
rect 18036 -13624 18052 -13590
rect 19420 -13624 19636 -13590
rect 18036 -13662 19636 -13624
rect 19694 -13590 21294 -13552
rect 19694 -13624 19913 -13590
rect 21278 -13624 21294 -13590
rect 19694 -13662 21294 -13624
rect 18036 -15100 19636 -15062
rect 18036 -15134 18052 -15100
rect 19420 -15134 19636 -15100
rect 18036 -15172 19636 -15134
rect 19694 -15100 21294 -15062
rect 19694 -15134 19913 -15100
rect 21278 -15134 21294 -15100
rect 19694 -15172 21294 -15134
rect 18036 -16610 19636 -16572
rect 18036 -16644 18052 -16610
rect 19420 -16644 19636 -16610
rect 18036 -16682 19636 -16644
rect 19694 -16610 21294 -16572
rect 19694 -16644 19913 -16610
rect 21278 -16644 21294 -16610
rect 19694 -16682 21294 -16644
rect 18036 -18120 19636 -18082
rect 18036 -18154 18052 -18120
rect 19420 -18154 19636 -18120
rect 18036 -18192 19636 -18154
rect 19694 -18120 21294 -18082
rect 19694 -18154 19913 -18120
rect 21278 -18154 21294 -18120
rect 19694 -18192 21294 -18154
rect 18036 -19630 19636 -19592
rect 18036 -19664 18052 -19630
rect 19420 -19664 19636 -19630
rect 18036 -19702 19636 -19664
rect 19694 -19630 21294 -19592
rect 19694 -19664 19913 -19630
rect 21278 -19664 21294 -19630
rect 19694 -19702 21294 -19664
rect 18036 -21140 19636 -21102
rect 18036 -21174 18052 -21140
rect 19420 -21174 19636 -21140
rect 18036 -21212 19636 -21174
rect 19694 -21140 21294 -21102
rect 19694 -21174 19913 -21140
rect 21278 -21174 21294 -21140
rect 19694 -21212 21294 -21174
rect 18036 -22650 19636 -22612
rect 18036 -22684 18052 -22650
rect 19420 -22684 19636 -22650
rect 18036 -22722 19636 -22684
rect 19694 -22650 21294 -22612
rect 19694 -22684 19913 -22650
rect 21278 -22684 21294 -22650
rect 19694 -22722 21294 -22684
rect 18036 -24160 19636 -24122
rect 18036 -24194 18052 -24160
rect 19420 -24194 19636 -24160
rect 18036 -24232 19636 -24194
rect 19694 -24160 21294 -24122
rect 19694 -24194 19913 -24160
rect 21278 -24194 21294 -24160
rect 19694 -24232 21294 -24194
rect 18036 -25670 19636 -25632
rect 18036 -25704 18052 -25670
rect 19420 -25704 19636 -25670
rect 18036 -25720 19636 -25704
rect 19694 -25670 21294 -25632
rect 19694 -25704 19913 -25670
rect 21278 -25704 21294 -25670
rect 19694 -25720 21294 -25704
<< polycont >>
rect -94156 20615 -93372 20649
rect -92498 20615 -91714 20649
rect -90840 20615 -90056 20649
rect -89182 20615 -88398 20649
rect -87524 20615 -86740 20649
rect -85866 20615 -85082 20649
rect -84208 20615 -83424 20649
rect -82550 20615 -81766 20649
rect -80892 20615 -80108 20649
rect -79234 20615 -78450 20649
rect -77576 20615 -76792 20649
rect -75918 20615 -75134 20649
rect -74260 20615 -73476 20649
rect -72602 20615 -71818 20649
rect -70944 20615 -70160 20649
rect -69286 20615 -68502 20649
rect -67628 20615 -66844 20649
rect -65970 20615 -65186 20649
rect -64312 20615 -63528 20649
rect -62654 20615 -61870 20649
rect -60996 20615 -60212 20649
rect -59338 20615 -58554 20649
rect -57680 20615 -56896 20649
rect -56022 20615 -55238 20649
rect -54364 20615 -53580 20649
rect -52706 20615 -51922 20649
rect -51048 20615 -50264 20649
rect -49390 20615 -48606 20649
rect -47732 20615 -46948 20649
rect -46074 20615 -45290 20649
rect -44416 20615 -43632 20649
rect -42758 20615 -41974 20649
rect -41100 20615 -40316 20649
rect -39442 20615 -38658 20649
rect -37784 20615 -37000 20649
rect -36126 20615 -35342 20649
rect -34468 20615 -33684 20649
rect -32810 20615 -32026 20649
rect -31152 20615 -30368 20649
rect -29494 20615 -28710 20649
rect -94156 19087 -93372 19121
rect -92498 19087 -91714 19121
rect -90840 19087 -90056 19121
rect -89182 19087 -88398 19121
rect -87524 19087 -86740 19121
rect -85866 19087 -85082 19121
rect -84208 19087 -83424 19121
rect -82550 19087 -81766 19121
rect -80892 19087 -80108 19121
rect -79234 19087 -78450 19121
rect -77576 19087 -76792 19121
rect -75918 19087 -75134 19121
rect -74260 19087 -73476 19121
rect -72602 19087 -71818 19121
rect -70944 19087 -70160 19121
rect -69286 19087 -68502 19121
rect -67628 19087 -66844 19121
rect -65970 19087 -65186 19121
rect -64312 19087 -63528 19121
rect -62654 19087 -61870 19121
rect -60996 19087 -60212 19121
rect -59338 19087 -58554 19121
rect -57680 19087 -56896 19121
rect -56022 19087 -55238 19121
rect -54364 19087 -53580 19121
rect -52706 19087 -51922 19121
rect -51048 19087 -50264 19121
rect -49390 19087 -48606 19121
rect -47732 19087 -46948 19121
rect -46074 19087 -45290 19121
rect -44416 19087 -43632 19121
rect -42758 19087 -41974 19121
rect -41100 19087 -40316 19121
rect -39442 19087 -38658 19121
rect -37784 19087 -37000 19121
rect -36126 19087 -35342 19121
rect -34468 19087 -33684 19121
rect -32810 19087 -32026 19121
rect -31152 19087 -30368 19121
rect -29494 19087 -28710 19121
rect -94156 18979 -93372 19013
rect -92498 18979 -91714 19013
rect -90840 18979 -90056 19013
rect -89182 18979 -88398 19013
rect -87524 18979 -86740 19013
rect -85866 18979 -85082 19013
rect -84208 18979 -83424 19013
rect -82550 18979 -81766 19013
rect -80892 18979 -80108 19013
rect -79234 18979 -78450 19013
rect -77576 18979 -76792 19013
rect -75918 18979 -75134 19013
rect -74260 18979 -73476 19013
rect -72602 18979 -71818 19013
rect -70944 18979 -70160 19013
rect -69286 18979 -68502 19013
rect -67628 18979 -66844 19013
rect -65970 18979 -65186 19013
rect -64312 18979 -63528 19013
rect -62654 18979 -61870 19013
rect -60996 18979 -60212 19013
rect -59338 18979 -58554 19013
rect -57680 18979 -56896 19013
rect -56022 18979 -55238 19013
rect -54364 18979 -53580 19013
rect -52706 18979 -51922 19013
rect -51048 18979 -50264 19013
rect -49390 18979 -48606 19013
rect -47732 18979 -46948 19013
rect -46074 18979 -45290 19013
rect -44416 18979 -43632 19013
rect -42758 18979 -41974 19013
rect -41100 18979 -40316 19013
rect -39442 18979 -38658 19013
rect -37784 18979 -37000 19013
rect -36126 18979 -35342 19013
rect -34468 18979 -33684 19013
rect -32810 18979 -32026 19013
rect -31152 18979 -30368 19013
rect -29494 18979 -28710 19013
rect -94156 17451 -93372 17485
rect -92498 17451 -91714 17485
rect -90840 17451 -90056 17485
rect -89182 17451 -88398 17485
rect -87524 17451 -86740 17485
rect -85866 17451 -85082 17485
rect -84208 17451 -83424 17485
rect -82550 17451 -81766 17485
rect -80892 17451 -80108 17485
rect -79234 17451 -78450 17485
rect -77576 17451 -76792 17485
rect -75918 17451 -75134 17485
rect -74260 17451 -73476 17485
rect -72602 17451 -71818 17485
rect -70944 17451 -70160 17485
rect -69286 17451 -68502 17485
rect -67628 17451 -66844 17485
rect -65970 17451 -65186 17485
rect -64312 17451 -63528 17485
rect -62654 17451 -61870 17485
rect -60996 17451 -60212 17485
rect -59338 17451 -58554 17485
rect -57680 17451 -56896 17485
rect -56022 17451 -55238 17485
rect -54364 17451 -53580 17485
rect -52706 17451 -51922 17485
rect -51048 17451 -50264 17485
rect -49390 17451 -48606 17485
rect -47732 17451 -46948 17485
rect -46074 17451 -45290 17485
rect -44416 17451 -43632 17485
rect -42758 17451 -41974 17485
rect -41100 17451 -40316 17485
rect -39442 17451 -38658 17485
rect -37784 17451 -37000 17485
rect -36126 17451 -35342 17485
rect -34468 17451 -33684 17485
rect -32810 17451 -32026 17485
rect -31152 17451 -30368 17485
rect -29494 17451 -28710 17485
rect -94154 17233 -93370 17267
rect -92496 17233 -91712 17267
rect -90838 17233 -90054 17267
rect -89180 17233 -88396 17267
rect -87522 17233 -86738 17267
rect -85864 17233 -85080 17267
rect -84206 17233 -83422 17267
rect -82548 17233 -81764 17267
rect -80890 17233 -80106 17267
rect -79232 17233 -78448 17267
rect -77574 17233 -76790 17267
rect -75916 17233 -75132 17267
rect -74258 17233 -73474 17267
rect -72600 17233 -71816 17267
rect -70942 17233 -70158 17267
rect -69284 17233 -68500 17267
rect -67626 17233 -66842 17267
rect -65968 17233 -65184 17267
rect -64310 17233 -63526 17267
rect -62652 17233 -61868 17267
rect -60994 17233 -60210 17267
rect -59336 17233 -58552 17267
rect -57678 17233 -56894 17267
rect -56020 17233 -55236 17267
rect -54362 17233 -53578 17267
rect -52704 17233 -51920 17267
rect -51046 17233 -50262 17267
rect -49388 17233 -48604 17267
rect -47730 17233 -46946 17267
rect -46072 17233 -45288 17267
rect -44414 17233 -43630 17267
rect -42756 17233 -41972 17267
rect -41098 17233 -40314 17267
rect -39440 17233 -38656 17267
rect -37782 17233 -36998 17267
rect -36124 17233 -35340 17267
rect -34466 17233 -33682 17267
rect -32808 17233 -32024 17267
rect -31150 17233 -30366 17267
rect -29492 17233 -28708 17267
rect -94154 15705 -93370 15739
rect -92496 15705 -91712 15739
rect -90838 15705 -90054 15739
rect -89180 15705 -88396 15739
rect -87522 15705 -86738 15739
rect -85864 15705 -85080 15739
rect -84206 15705 -83422 15739
rect -82548 15705 -81764 15739
rect -80890 15705 -80106 15739
rect -79232 15705 -78448 15739
rect -77574 15705 -76790 15739
rect -75916 15705 -75132 15739
rect -74258 15705 -73474 15739
rect -72600 15705 -71816 15739
rect -70942 15705 -70158 15739
rect -69284 15705 -68500 15739
rect -67626 15705 -66842 15739
rect -65968 15705 -65184 15739
rect -64310 15705 -63526 15739
rect -62652 15705 -61868 15739
rect -60994 15705 -60210 15739
rect -59336 15705 -58552 15739
rect -57678 15705 -56894 15739
rect -56020 15705 -55236 15739
rect -54362 15705 -53578 15739
rect -52704 15705 -51920 15739
rect -51046 15705 -50262 15739
rect -49388 15705 -48604 15739
rect -47730 15705 -46946 15739
rect -46072 15705 -45288 15739
rect -44414 15705 -43630 15739
rect -42756 15705 -41972 15739
rect -41098 15705 -40314 15739
rect -39440 15705 -38656 15739
rect -37782 15705 -36998 15739
rect -36124 15705 -35340 15739
rect -34466 15705 -33682 15739
rect -32808 15705 -32024 15739
rect -31150 15705 -30366 15739
rect -29492 15705 -28708 15739
rect -94154 15597 -93370 15631
rect -92496 15597 -91712 15631
rect -90838 15597 -90054 15631
rect -89180 15597 -88396 15631
rect -87522 15597 -86738 15631
rect -85864 15597 -85080 15631
rect -84206 15597 -83422 15631
rect -82548 15597 -81764 15631
rect -80890 15597 -80106 15631
rect -79232 15597 -78448 15631
rect -77574 15597 -76790 15631
rect -75916 15597 -75132 15631
rect -74258 15597 -73474 15631
rect -72600 15597 -71816 15631
rect -70942 15597 -70158 15631
rect -69284 15597 -68500 15631
rect -67626 15597 -66842 15631
rect -65968 15597 -65184 15631
rect -64310 15597 -63526 15631
rect -62652 15597 -61868 15631
rect -60994 15597 -60210 15631
rect -59336 15597 -58552 15631
rect -57678 15597 -56894 15631
rect -56020 15597 -55236 15631
rect -54362 15597 -53578 15631
rect -52704 15597 -51920 15631
rect -51046 15597 -50262 15631
rect -49388 15597 -48604 15631
rect -47730 15597 -46946 15631
rect -46072 15597 -45288 15631
rect -44414 15597 -43630 15631
rect -42756 15597 -41972 15631
rect -41098 15597 -40314 15631
rect -39440 15597 -38656 15631
rect -37782 15597 -36998 15631
rect -36124 15597 -35340 15631
rect -34466 15597 -33682 15631
rect -32808 15597 -32024 15631
rect -31150 15597 -30366 15631
rect -29492 15597 -28708 15631
rect -94154 14069 -93370 14103
rect -92496 14069 -91712 14103
rect -90838 14069 -90054 14103
rect -89180 14069 -88396 14103
rect -87522 14069 -86738 14103
rect -85864 14069 -85080 14103
rect -84206 14069 -83422 14103
rect -82548 14069 -81764 14103
rect -80890 14069 -80106 14103
rect -79232 14069 -78448 14103
rect -77574 14069 -76790 14103
rect -75916 14069 -75132 14103
rect -74258 14069 -73474 14103
rect -72600 14069 -71816 14103
rect -70942 14069 -70158 14103
rect -69284 14069 -68500 14103
rect -67626 14069 -66842 14103
rect -65968 14069 -65184 14103
rect -64310 14069 -63526 14103
rect -62652 14069 -61868 14103
rect -60994 14069 -60210 14103
rect -59336 14069 -58552 14103
rect -57678 14069 -56894 14103
rect -56020 14069 -55236 14103
rect -54362 14069 -53578 14103
rect -52704 14069 -51920 14103
rect -51046 14069 -50262 14103
rect -49388 14069 -48604 14103
rect -47730 14069 -46946 14103
rect -46072 14069 -45288 14103
rect -44414 14069 -43630 14103
rect -42756 14069 -41972 14103
rect -41098 14069 -40314 14103
rect -39440 14069 -38656 14103
rect -37782 14069 -36998 14103
rect -36124 14069 -35340 14103
rect -34466 14069 -33682 14103
rect -32808 14069 -32024 14103
rect -31150 14069 -30366 14103
rect -29492 14069 -28708 14103
rect -94154 13961 -93370 13995
rect -92496 13961 -91712 13995
rect -90838 13961 -90054 13995
rect -89180 13961 -88396 13995
rect -87522 13961 -86738 13995
rect -85864 13961 -85080 13995
rect -84206 13961 -83422 13995
rect -82548 13961 -81764 13995
rect -80890 13961 -80106 13995
rect -79232 13961 -78448 13995
rect -77574 13961 -76790 13995
rect -75916 13961 -75132 13995
rect -74258 13961 -73474 13995
rect -72600 13961 -71816 13995
rect -70942 13961 -70158 13995
rect -69284 13961 -68500 13995
rect -67626 13961 -66842 13995
rect -65968 13961 -65184 13995
rect -64310 13961 -63526 13995
rect -62652 13961 -61868 13995
rect -60994 13961 -60210 13995
rect -59336 13961 -58552 13995
rect -57678 13961 -56894 13995
rect -56020 13961 -55236 13995
rect -54362 13961 -53578 13995
rect -52704 13961 -51920 13995
rect -51046 13961 -50262 13995
rect -49388 13961 -48604 13995
rect -47730 13961 -46946 13995
rect -46072 13961 -45288 13995
rect -44414 13961 -43630 13995
rect -42756 13961 -41972 13995
rect -41098 13961 -40314 13995
rect -39440 13961 -38656 13995
rect -37782 13961 -36998 13995
rect -36124 13961 -35340 13995
rect -34466 13961 -33682 13995
rect -32808 13961 -32024 13995
rect -31150 13961 -30366 13995
rect -29492 13961 -28708 13995
rect -94154 12433 -93370 12467
rect -92496 12433 -91712 12467
rect -90838 12433 -90054 12467
rect -89180 12433 -88396 12467
rect -87522 12433 -86738 12467
rect -85864 12433 -85080 12467
rect -84206 12433 -83422 12467
rect -82548 12433 -81764 12467
rect -80890 12433 -80106 12467
rect -79232 12433 -78448 12467
rect -77574 12433 -76790 12467
rect -75916 12433 -75132 12467
rect -74258 12433 -73474 12467
rect -72600 12433 -71816 12467
rect -70942 12433 -70158 12467
rect -69284 12433 -68500 12467
rect -67626 12433 -66842 12467
rect -65968 12433 -65184 12467
rect -64310 12433 -63526 12467
rect -62652 12433 -61868 12467
rect -60994 12433 -60210 12467
rect -59336 12433 -58552 12467
rect -57678 12433 -56894 12467
rect -56020 12433 -55236 12467
rect -54362 12433 -53578 12467
rect -52704 12433 -51920 12467
rect -51046 12433 -50262 12467
rect -49388 12433 -48604 12467
rect -47730 12433 -46946 12467
rect -46072 12433 -45288 12467
rect -44414 12433 -43630 12467
rect -42756 12433 -41972 12467
rect -41098 12433 -40314 12467
rect -39440 12433 -38656 12467
rect -37782 12433 -36998 12467
rect -36124 12433 -35340 12467
rect -34466 12433 -33682 12467
rect -32808 12433 -32024 12467
rect -31150 12433 -30366 12467
rect -29492 12433 -28708 12467
rect -94154 12325 -93370 12359
rect -92496 12325 -91712 12359
rect -90838 12325 -90054 12359
rect -89180 12325 -88396 12359
rect -87522 12325 -86738 12359
rect -85864 12325 -85080 12359
rect -84206 12325 -83422 12359
rect -82548 12325 -81764 12359
rect -80890 12325 -80106 12359
rect -79232 12325 -78448 12359
rect -77574 12325 -76790 12359
rect -75916 12325 -75132 12359
rect -74258 12325 -73474 12359
rect -72600 12325 -71816 12359
rect -70942 12325 -70158 12359
rect -69284 12325 -68500 12359
rect -67626 12325 -66842 12359
rect -65968 12325 -65184 12359
rect -64310 12325 -63526 12359
rect -62652 12325 -61868 12359
rect -60994 12325 -60210 12359
rect -59336 12325 -58552 12359
rect -57678 12325 -56894 12359
rect -56020 12325 -55236 12359
rect -54362 12325 -53578 12359
rect -52704 12325 -51920 12359
rect -51046 12325 -50262 12359
rect -49388 12325 -48604 12359
rect -47730 12325 -46946 12359
rect -46072 12325 -45288 12359
rect -44414 12325 -43630 12359
rect -42756 12325 -41972 12359
rect -41098 12325 -40314 12359
rect -39440 12325 -38656 12359
rect -37782 12325 -36998 12359
rect -36124 12325 -35340 12359
rect -34466 12325 -33682 12359
rect -32808 12325 -32024 12359
rect -31150 12325 -30366 12359
rect -29492 12325 -28708 12359
rect -94154 10797 -93370 10831
rect -92496 10797 -91712 10831
rect -90838 10797 -90054 10831
rect -89180 10797 -88396 10831
rect -87522 10797 -86738 10831
rect -85864 10797 -85080 10831
rect -84206 10797 -83422 10831
rect -82548 10797 -81764 10831
rect -80890 10797 -80106 10831
rect -79232 10797 -78448 10831
rect -77574 10797 -76790 10831
rect -75916 10797 -75132 10831
rect -74258 10797 -73474 10831
rect -72600 10797 -71816 10831
rect -70942 10797 -70158 10831
rect -69284 10797 -68500 10831
rect -67626 10797 -66842 10831
rect -65968 10797 -65184 10831
rect -64310 10797 -63526 10831
rect -62652 10797 -61868 10831
rect -60994 10797 -60210 10831
rect -59336 10797 -58552 10831
rect -57678 10797 -56894 10831
rect -56020 10797 -55236 10831
rect -54362 10797 -53578 10831
rect -52704 10797 -51920 10831
rect -51046 10797 -50262 10831
rect -49388 10797 -48604 10831
rect -47730 10797 -46946 10831
rect -46072 10797 -45288 10831
rect -44414 10797 -43630 10831
rect -42756 10797 -41972 10831
rect -41098 10797 -40314 10831
rect -39440 10797 -38656 10831
rect -37782 10797 -36998 10831
rect -36124 10797 -35340 10831
rect -34466 10797 -33682 10831
rect -32808 10797 -32024 10831
rect -31150 10797 -30366 10831
rect -29492 10797 -28708 10831
rect -94154 10687 -93370 10721
rect -92496 10687 -91712 10721
rect -90838 10687 -90054 10721
rect -89180 10687 -88396 10721
rect -87522 10687 -86738 10721
rect -85864 10687 -85080 10721
rect -84206 10687 -83422 10721
rect -82548 10687 -81764 10721
rect -80890 10687 -80106 10721
rect -79232 10687 -78448 10721
rect -77574 10687 -76790 10721
rect -75916 10687 -75132 10721
rect -74258 10687 -73474 10721
rect -72600 10687 -71816 10721
rect -70942 10687 -70158 10721
rect -69284 10687 -68500 10721
rect -67626 10687 -66842 10721
rect -65968 10687 -65184 10721
rect -64310 10687 -63526 10721
rect -62652 10687 -61868 10721
rect -60994 10687 -60210 10721
rect -59336 10687 -58552 10721
rect -57678 10687 -56894 10721
rect -56020 10687 -55236 10721
rect -54362 10687 -53578 10721
rect -52704 10687 -51920 10721
rect -51046 10687 -50262 10721
rect -49388 10687 -48604 10721
rect -47730 10687 -46946 10721
rect -46072 10687 -45288 10721
rect -44414 10687 -43630 10721
rect -42756 10687 -41972 10721
rect -41098 10687 -40314 10721
rect -39440 10687 -38656 10721
rect -37782 10687 -36998 10721
rect -36124 10687 -35340 10721
rect -34466 10687 -33682 10721
rect -32808 10687 -32024 10721
rect -31150 10687 -30366 10721
rect -29492 10687 -28708 10721
rect -94154 9159 -93370 9193
rect -92496 9159 -91712 9193
rect -90838 9159 -90054 9193
rect -89180 9159 -88396 9193
rect -87522 9159 -86738 9193
rect -85864 9159 -85080 9193
rect -84206 9159 -83422 9193
rect -82548 9159 -81764 9193
rect -80890 9159 -80106 9193
rect -79232 9159 -78448 9193
rect -77574 9159 -76790 9193
rect -75916 9159 -75132 9193
rect -74258 9159 -73474 9193
rect -72600 9159 -71816 9193
rect -70942 9159 -70158 9193
rect -69284 9159 -68500 9193
rect -67626 9159 -66842 9193
rect -65968 9159 -65184 9193
rect -64310 9159 -63526 9193
rect -62652 9159 -61868 9193
rect -60994 9159 -60210 9193
rect -59336 9159 -58552 9193
rect -57678 9159 -56894 9193
rect -56020 9159 -55236 9193
rect -54362 9159 -53578 9193
rect -52704 9159 -51920 9193
rect -51046 9159 -50262 9193
rect -49388 9159 -48604 9193
rect -47730 9159 -46946 9193
rect -46072 9159 -45288 9193
rect -44414 9159 -43630 9193
rect -42756 9159 -41972 9193
rect -41098 9159 -40314 9193
rect -39440 9159 -38656 9193
rect -37782 9159 -36998 9193
rect -36124 9159 -35340 9193
rect -34466 9159 -33682 9193
rect -32808 9159 -32024 9193
rect -31150 9159 -30366 9193
rect -29492 9159 -28708 9193
rect -94154 9051 -93370 9085
rect -92496 9051 -91712 9085
rect -90838 9051 -90054 9085
rect -89180 9051 -88396 9085
rect -87522 9051 -86738 9085
rect -85864 9051 -85080 9085
rect -84206 9051 -83422 9085
rect -82548 9051 -81764 9085
rect -80890 9051 -80106 9085
rect -79232 9051 -78448 9085
rect -77574 9051 -76790 9085
rect -75916 9051 -75132 9085
rect -74258 9051 -73474 9085
rect -72600 9051 -71816 9085
rect -70942 9051 -70158 9085
rect -69284 9051 -68500 9085
rect -67626 9051 -66842 9085
rect -65968 9051 -65184 9085
rect -64310 9051 -63526 9085
rect -62652 9051 -61868 9085
rect -60994 9051 -60210 9085
rect -59336 9051 -58552 9085
rect -57678 9051 -56894 9085
rect -56020 9051 -55236 9085
rect -54362 9051 -53578 9085
rect -52704 9051 -51920 9085
rect -51046 9051 -50262 9085
rect -49388 9051 -48604 9085
rect -47730 9051 -46946 9085
rect -46072 9051 -45288 9085
rect -44414 9051 -43630 9085
rect -42756 9051 -41972 9085
rect -41098 9051 -40314 9085
rect -39440 9051 -38656 9085
rect -37782 9051 -36998 9085
rect -36124 9051 -35340 9085
rect -34466 9051 -33682 9085
rect -32808 9051 -32024 9085
rect -31150 9051 -30366 9085
rect -29492 9051 -28708 9085
rect -94154 7523 -93370 7557
rect -92496 7523 -91712 7557
rect -90838 7523 -90054 7557
rect -89180 7523 -88396 7557
rect -87522 7523 -86738 7557
rect -85864 7523 -85080 7557
rect -84206 7523 -83422 7557
rect -82548 7523 -81764 7557
rect -80890 7523 -80106 7557
rect -79232 7523 -78448 7557
rect -77574 7523 -76790 7557
rect -75916 7523 -75132 7557
rect -74258 7523 -73474 7557
rect -72600 7523 -71816 7557
rect -70942 7523 -70158 7557
rect -69284 7523 -68500 7557
rect -67626 7523 -66842 7557
rect -65968 7523 -65184 7557
rect -64310 7523 -63526 7557
rect -62652 7523 -61868 7557
rect -60994 7523 -60210 7557
rect -59336 7523 -58552 7557
rect -57678 7523 -56894 7557
rect -56020 7523 -55236 7557
rect -54362 7523 -53578 7557
rect -52704 7523 -51920 7557
rect -51046 7523 -50262 7557
rect -49388 7523 -48604 7557
rect -47730 7523 -46946 7557
rect -46072 7523 -45288 7557
rect -44414 7523 -43630 7557
rect -42756 7523 -41972 7557
rect -41098 7523 -40314 7557
rect -39440 7523 -38656 7557
rect -37782 7523 -36998 7557
rect -36124 7523 -35340 7557
rect -34466 7523 -33682 7557
rect -32808 7523 -32024 7557
rect -31150 7523 -30366 7557
rect -29492 7523 -28708 7557
rect -94154 7415 -93370 7449
rect -92496 7415 -91712 7449
rect -90838 7415 -90054 7449
rect -89180 7415 -88396 7449
rect -87522 7415 -86738 7449
rect -85864 7415 -85080 7449
rect -84206 7415 -83422 7449
rect -82548 7415 -81764 7449
rect -80890 7415 -80106 7449
rect -79232 7415 -78448 7449
rect -77574 7415 -76790 7449
rect -75916 7415 -75132 7449
rect -74258 7415 -73474 7449
rect -72600 7415 -71816 7449
rect -70942 7415 -70158 7449
rect -69284 7415 -68500 7449
rect -67626 7415 -66842 7449
rect -65968 7415 -65184 7449
rect -64310 7415 -63526 7449
rect -62652 7415 -61868 7449
rect -60994 7415 -60210 7449
rect -59336 7415 -58552 7449
rect -57678 7415 -56894 7449
rect -56020 7415 -55236 7449
rect -54362 7415 -53578 7449
rect -52704 7415 -51920 7449
rect -51046 7415 -50262 7449
rect -49388 7415 -48604 7449
rect -47730 7415 -46946 7449
rect -46072 7415 -45288 7449
rect -44414 7415 -43630 7449
rect -42756 7415 -41972 7449
rect -41098 7415 -40314 7449
rect -39440 7415 -38656 7449
rect -37782 7415 -36998 7449
rect -36124 7415 -35340 7449
rect -34466 7415 -33682 7449
rect -32808 7415 -32024 7449
rect -31150 7415 -30366 7449
rect -29492 7415 -28708 7449
rect -94154 5887 -93370 5921
rect -92496 5887 -91712 5921
rect -90838 5887 -90054 5921
rect -89180 5887 -88396 5921
rect -87522 5887 -86738 5921
rect -85864 5887 -85080 5921
rect -84206 5887 -83422 5921
rect -82548 5887 -81764 5921
rect -80890 5887 -80106 5921
rect -79232 5887 -78448 5921
rect -77574 5887 -76790 5921
rect -75916 5887 -75132 5921
rect -74258 5887 -73474 5921
rect -72600 5887 -71816 5921
rect -70942 5887 -70158 5921
rect -69284 5887 -68500 5921
rect -67626 5887 -66842 5921
rect -65968 5887 -65184 5921
rect -64310 5887 -63526 5921
rect -62652 5887 -61868 5921
rect -60994 5887 -60210 5921
rect -59336 5887 -58552 5921
rect -57678 5887 -56894 5921
rect -56020 5887 -55236 5921
rect -54362 5887 -53578 5921
rect -52704 5887 -51920 5921
rect -51046 5887 -50262 5921
rect -49388 5887 -48604 5921
rect -47730 5887 -46946 5921
rect -46072 5887 -45288 5921
rect -44414 5887 -43630 5921
rect -42756 5887 -41972 5921
rect -41098 5887 -40314 5921
rect -39440 5887 -38656 5921
rect -37782 5887 -36998 5921
rect -36124 5887 -35340 5921
rect -34466 5887 -33682 5921
rect -32808 5887 -32024 5921
rect -31150 5887 -30366 5921
rect -29492 5887 -28708 5921
rect -94154 5779 -93370 5813
rect -92496 5779 -91712 5813
rect -90838 5779 -90054 5813
rect -89180 5779 -88396 5813
rect -87522 5779 -86738 5813
rect -85864 5779 -85080 5813
rect -84206 5779 -83422 5813
rect -82548 5779 -81764 5813
rect -80890 5779 -80106 5813
rect -79232 5779 -78448 5813
rect -77574 5779 -76790 5813
rect -75916 5779 -75132 5813
rect -74258 5779 -73474 5813
rect -72600 5779 -71816 5813
rect -70942 5779 -70158 5813
rect -69284 5779 -68500 5813
rect -67626 5779 -66842 5813
rect -65968 5779 -65184 5813
rect -64310 5779 -63526 5813
rect -62652 5779 -61868 5813
rect -60994 5779 -60210 5813
rect -59336 5779 -58552 5813
rect -57678 5779 -56894 5813
rect -56020 5779 -55236 5813
rect -54362 5779 -53578 5813
rect -52704 5779 -51920 5813
rect -51046 5779 -50262 5813
rect -49388 5779 -48604 5813
rect -47730 5779 -46946 5813
rect -46072 5779 -45288 5813
rect -44414 5779 -43630 5813
rect -42756 5779 -41972 5813
rect -41098 5779 -40314 5813
rect -39440 5779 -38656 5813
rect -37782 5779 -36998 5813
rect -36124 5779 -35340 5813
rect -34466 5779 -33682 5813
rect -32808 5779 -32024 5813
rect -31150 5779 -30366 5813
rect -29492 5779 -28708 5813
rect 2724 5963 2808 5997
rect 3380 5971 3464 6005
rect 3638 5971 3722 6005
rect 4380 5971 4464 6005
rect 4638 5971 4722 6005
rect 5286 5975 5370 6009
rect -94154 4251 -93370 4285
rect -92496 4251 -91712 4285
rect -90838 4251 -90054 4285
rect -89180 4251 -88396 4285
rect -87522 4251 -86738 4285
rect -85864 4251 -85080 4285
rect -84206 4251 -83422 4285
rect -82548 4251 -81764 4285
rect -80890 4251 -80106 4285
rect -79232 4251 -78448 4285
rect -77574 4251 -76790 4285
rect -75916 4251 -75132 4285
rect -74258 4251 -73474 4285
rect -72600 4251 -71816 4285
rect -70942 4251 -70158 4285
rect -69284 4251 -68500 4285
rect -67626 4251 -66842 4285
rect -65968 4251 -65184 4285
rect -64310 4251 -63526 4285
rect -62652 4251 -61868 4285
rect -60994 4251 -60210 4285
rect -59336 4251 -58552 4285
rect -57678 4251 -56894 4285
rect -56020 4251 -55236 4285
rect -54362 4251 -53578 4285
rect -52704 4251 -51920 4285
rect -51046 4251 -50262 4285
rect -49388 4251 -48604 4285
rect -47730 4251 -46946 4285
rect -46072 4251 -45288 4285
rect -44414 4251 -43630 4285
rect -42756 4251 -41972 4285
rect -41098 4251 -40314 4285
rect -39440 4251 -38656 4285
rect -37782 4251 -36998 4285
rect -36124 4251 -35340 4285
rect -34466 4251 -33682 4285
rect -32808 4251 -32024 4285
rect -31150 4251 -30366 4285
rect -29492 4251 -28708 4285
rect -61626 3937 -61592 3971
rect -61434 3937 -61400 3971
rect 1118 5085 1152 5119
rect 1350 5083 1384 5117
rect 1578 5081 1612 5115
rect 1796 5083 1830 5117
rect 8660 5703 8744 5737
rect 9139 5695 9223 5729
rect 6304 5103 6338 5137
rect 6536 5101 6570 5135
rect 6764 5099 6798 5133
rect 6982 5101 7016 5135
rect 1118 4557 1152 4591
rect 9397 5695 9481 5729
rect 9797 5697 9881 5731
rect 10055 5697 10139 5731
rect 10454 5677 10538 5711
rect 1350 4555 1384 4589
rect 1578 4553 1612 4587
rect 1796 4555 1830 4589
rect 6304 4575 6338 4609
rect 6536 4573 6570 4607
rect 6764 4571 6798 4605
rect 13934 5575 14018 5609
rect 14378 5557 14562 5591
rect 11480 5115 11514 5149
rect 11712 5113 11746 5147
rect 11940 5111 11974 5145
rect 12158 5113 12192 5147
rect 6982 4573 7016 4607
rect 11480 4587 11514 4621
rect 11712 4585 11746 4619
rect 11940 4583 11974 4617
rect 12158 4585 12192 4619
rect 14950 5557 15134 5591
rect 15522 5587 15606 5621
rect 1142 4438 1176 4472
rect 1358 4440 1392 4474
rect 1576 4440 1610 4474
rect 1798 4438 1832 4472
rect 6328 4456 6362 4490
rect 6544 4458 6578 4492
rect 6762 4458 6796 4492
rect 6984 4456 7018 4490
rect 11504 4468 11538 4502
rect 11720 4470 11754 4504
rect 11938 4470 11972 4504
rect 17136 4907 17170 4941
rect 17368 4905 17402 4939
rect 17596 4903 17630 4937
rect 12160 4468 12194 4502
rect 17814 4905 17848 4939
rect 1142 4128 1176 4162
rect 1358 4130 1392 4164
rect 1576 4130 1610 4164
rect 1798 4128 1832 4162
rect 6328 4146 6362 4180
rect 6544 4148 6578 4182
rect 17136 4379 17170 4413
rect 17368 4377 17402 4411
rect 17596 4375 17630 4409
rect 17814 4377 17848 4411
rect 17160 4260 17194 4294
rect 17376 4262 17410 4296
rect 17594 4262 17628 4296
rect 17816 4260 17850 4294
rect 6762 4148 6796 4182
rect 6984 4146 7018 4180
rect 11504 4158 11538 4192
rect 11720 4160 11754 4194
rect 11938 4160 11972 4194
rect 12160 4158 12194 4192
rect 17160 3950 17194 3984
rect 17376 3952 17410 3986
rect 17594 3952 17628 3986
rect 17816 3950 17850 3984
rect -61722 3409 -61688 3443
rect -61530 3409 -61496 3443
rect -61674 3284 -61640 3318
rect -61482 3284 -61448 3318
rect 8898 3722 8966 3756
rect 9156 3722 9224 3756
rect 9414 3722 9482 3756
rect 9912 3722 9980 3756
rect 10170 3722 10238 3756
rect 10428 3722 10496 3756
rect 8898 3166 8966 3200
rect 9156 3166 9224 3200
rect 9414 3166 9482 3200
rect 9912 3166 9980 3200
rect 10170 3166 10238 3200
rect 10428 3166 10496 3200
rect 13422 3152 13506 3186
rect -61770 2974 -61736 3008
rect -61578 2974 -61544 3008
rect 2730 2570 2814 2604
rect 3356 2572 3740 2606
rect 4328 2572 4712 2606
rect 5264 2570 5348 2604
rect 9261 1922 9445 1956
rect 9856 1922 10040 1956
rect 16020 3102 16104 3136
rect 13972 3018 14056 3052
rect 14230 3018 14314 3052
rect 14488 3018 14572 3052
rect 14972 3018 15056 3052
rect 15230 3018 15314 3052
rect 15488 3018 15572 3052
rect 13972 2062 14056 2096
rect 14230 2062 14314 2096
rect 14488 2062 14572 2096
rect 14972 2062 15056 2096
rect 15230 2062 15314 2096
rect 15488 2062 15572 2096
rect 13972 1106 14056 1140
rect 14230 1106 14314 1140
rect 14488 1106 14572 1140
rect 14972 1106 15056 1140
rect 15230 1106 15314 1140
rect 15488 1106 15572 1140
rect 26930 2853 26964 2887
rect 27542 2861 27576 2895
rect 28120 2857 28154 2891
rect 28694 2865 28728 2899
rect 29272 2865 29306 2899
rect 27134 2427 27168 2461
rect 29850 2865 29884 2899
rect 27746 2435 27780 2469
rect 28324 2431 28358 2465
rect 30432 2869 30466 2903
rect 28898 2439 28932 2473
rect 31008 2865 31042 2899
rect 29476 2439 29510 2473
rect 31578 2861 31612 2895
rect 30054 2439 30088 2473
rect 30636 2443 30670 2477
rect 31212 2439 31246 2473
rect 31782 2435 31816 2469
rect 27030 2246 27064 2280
rect 27642 2254 27676 2288
rect 28220 2250 28254 2284
rect 28794 2258 28828 2292
rect 29372 2258 29406 2292
rect 29950 2258 29984 2292
rect 30532 2262 30566 2296
rect 31108 2258 31142 2292
rect 26934 1988 26968 2022
rect 31678 2254 31712 2288
rect 27546 1996 27580 2030
rect 28124 1992 28158 2026
rect 28698 2000 28732 2034
rect 29276 2000 29310 2034
rect 29854 2000 29888 2034
rect 30436 2004 30470 2038
rect 31012 2000 31046 2034
rect 31582 1996 31616 2030
rect 28324 799 28358 833
rect 28726 797 28760 831
rect 28524 373 28558 407
rect 29088 408 29122 442
rect 29280 408 29314 442
rect 29472 408 29506 442
rect 29664 408 29698 442
rect 28324 293 28358 327
rect 28724 293 28758 327
rect 28524 -133 28558 -99
rect 28324 -215 28358 -181
rect 28724 -215 28758 -181
rect 28992 -350 29026 -316
rect 29184 -350 29218 -316
rect 29376 -350 29410 -316
rect 29568 -350 29602 -316
rect 29760 -350 29794 -316
rect 28524 -641 28558 -607
rect 8766 -1304 8800 -1270
rect 8868 -1289 8902 -1255
rect 9256 -1188 9290 -1154
rect 9075 -1243 9109 -1209
rect 9505 -1214 9539 -1180
rect 9234 -1350 9268 -1316
rect 9336 -1356 9370 -1322
rect 9591 -1350 9625 -1316
rect 9687 -1302 9721 -1268
rect 9970 -1188 10004 -1154
rect 9835 -1362 9869 -1328
rect 9931 -1314 9965 -1280
rect 10248 -1204 10282 -1170
rect 10075 -1340 10109 -1306
rect 10171 -1312 10205 -1278
rect 10371 -1304 10405 -1270
rect 10711 -1304 10745 -1270
rect 11232 -1304 11266 -1270
rect 11334 -1289 11368 -1255
rect 11722 -1188 11756 -1154
rect 11541 -1243 11575 -1209
rect 11971 -1214 12005 -1180
rect 11700 -1350 11734 -1316
rect 11802 -1356 11836 -1322
rect 12057 -1350 12091 -1316
rect 12153 -1302 12187 -1268
rect 12436 -1188 12470 -1154
rect 12301 -1362 12335 -1328
rect 12397 -1314 12431 -1280
rect 12714 -1204 12748 -1170
rect 12541 -1340 12575 -1306
rect 12637 -1312 12671 -1278
rect 12837 -1304 12871 -1270
rect 13177 -1304 13211 -1270
rect 10189 -2106 10223 -2072
rect 11232 -2106 11266 -2072
rect 11334 -2091 11368 -2057
rect 11722 -1990 11756 -1956
rect 11541 -2045 11575 -2011
rect 11971 -2016 12005 -1982
rect 11700 -2152 11734 -2118
rect 11802 -2158 11836 -2124
rect 12057 -2152 12091 -2118
rect 12153 -2104 12187 -2070
rect 12436 -1990 12470 -1956
rect 12301 -2164 12335 -2130
rect 12397 -2116 12431 -2082
rect 12714 -2006 12748 -1972
rect 12541 -2142 12575 -2108
rect 12637 -2114 12671 -2080
rect 12837 -2106 12871 -2072
rect 13177 -2106 13211 -2072
rect -9126 -4574 -9092 -4540
rect -9024 -4559 -8990 -4525
rect -8636 -4458 -8602 -4424
rect -8817 -4513 -8783 -4479
rect -8387 -4484 -8353 -4450
rect -8658 -4620 -8624 -4586
rect -8556 -4626 -8522 -4592
rect -8301 -4620 -8267 -4586
rect -8205 -4572 -8171 -4538
rect -7922 -4458 -7888 -4424
rect -8057 -4632 -8023 -4598
rect -7961 -4584 -7927 -4550
rect -7644 -4474 -7610 -4440
rect -7817 -4610 -7783 -4576
rect -7721 -4582 -7687 -4548
rect -7521 -4574 -7487 -4540
rect -7181 -4574 -7147 -4540
rect -7010 -4574 -6976 -4540
rect -6908 -4559 -6874 -4525
rect -6520 -4458 -6486 -4424
rect -6701 -4513 -6667 -4479
rect -6271 -4484 -6237 -4450
rect -6542 -4620 -6508 -4586
rect -6440 -4626 -6406 -4592
rect -6185 -4620 -6151 -4586
rect -6089 -4572 -6055 -4538
rect -5806 -4458 -5772 -4424
rect -5941 -4632 -5907 -4598
rect -5845 -4584 -5811 -4550
rect -5528 -4474 -5494 -4440
rect -5701 -4610 -5667 -4576
rect -5605 -4582 -5571 -4548
rect -5405 -4574 -5371 -4540
rect -5065 -4574 -5031 -4540
rect -4894 -4574 -4860 -4540
rect -4792 -4559 -4758 -4525
rect -4404 -4458 -4370 -4424
rect -4585 -4513 -4551 -4479
rect -4155 -4484 -4121 -4450
rect -4426 -4620 -4392 -4586
rect -4324 -4626 -4290 -4592
rect -4069 -4620 -4035 -4586
rect -3973 -4572 -3939 -4538
rect -3690 -4458 -3656 -4424
rect -3825 -4632 -3791 -4598
rect -3729 -4584 -3695 -4550
rect -3412 -4474 -3378 -4440
rect -3585 -4610 -3551 -4576
rect -3489 -4582 -3455 -4548
rect -3289 -4574 -3255 -4540
rect -2949 -4574 -2915 -4540
rect -2778 -4574 -2744 -4540
rect -2676 -4559 -2642 -4525
rect -2288 -4458 -2254 -4424
rect -2469 -4513 -2435 -4479
rect -2039 -4484 -2005 -4450
rect -2310 -4620 -2276 -4586
rect -2208 -4626 -2174 -4592
rect -1953 -4620 -1919 -4586
rect -1857 -4572 -1823 -4538
rect -1574 -4458 -1540 -4424
rect -1709 -4632 -1675 -4598
rect -1613 -4584 -1579 -4550
rect -1296 -4474 -1262 -4440
rect -1469 -4610 -1435 -4576
rect -1373 -4582 -1339 -4548
rect -1173 -4574 -1139 -4540
rect -833 -4574 -799 -4540
rect -662 -4574 -628 -4540
rect -560 -4559 -526 -4525
rect -172 -4458 -138 -4424
rect -353 -4513 -319 -4479
rect 77 -4484 111 -4450
rect -194 -4620 -160 -4586
rect -92 -4626 -58 -4592
rect 163 -4620 197 -4586
rect 259 -4572 293 -4538
rect 542 -4458 576 -4424
rect 407 -4632 441 -4598
rect 503 -4584 537 -4550
rect 820 -4474 854 -4440
rect 647 -4610 681 -4576
rect 743 -4582 777 -4548
rect 943 -4574 977 -4540
rect 1283 -4574 1317 -4540
rect 1454 -4574 1488 -4540
rect 1556 -4559 1590 -4525
rect 1944 -4458 1978 -4424
rect 1763 -4513 1797 -4479
rect 2193 -4484 2227 -4450
rect 1922 -4620 1956 -4586
rect 2024 -4626 2058 -4592
rect 2279 -4620 2313 -4586
rect 2375 -4572 2409 -4538
rect 2658 -4458 2692 -4424
rect 2523 -4632 2557 -4598
rect 2619 -4584 2653 -4550
rect 2936 -4474 2970 -4440
rect 2763 -4610 2797 -4576
rect 2859 -4582 2893 -4548
rect 3059 -4574 3093 -4540
rect 3399 -4574 3433 -4540
rect 3570 -4574 3604 -4540
rect 3672 -4559 3706 -4525
rect 4060 -4458 4094 -4424
rect 3879 -4513 3913 -4479
rect 4309 -4484 4343 -4450
rect 4038 -4620 4072 -4586
rect 4140 -4626 4174 -4592
rect 4395 -4620 4429 -4586
rect 4491 -4572 4525 -4538
rect 4774 -4458 4808 -4424
rect 4639 -4632 4673 -4598
rect 4735 -4584 4769 -4550
rect 5052 -4474 5086 -4440
rect 4879 -4610 4913 -4576
rect 4975 -4582 5009 -4548
rect 5175 -4574 5209 -4540
rect 5515 -4574 5549 -4540
rect 5686 -4574 5720 -4540
rect 5788 -4559 5822 -4525
rect 6176 -4458 6210 -4424
rect 5995 -4513 6029 -4479
rect 6425 -4484 6459 -4450
rect 6154 -4620 6188 -4586
rect 6256 -4626 6290 -4592
rect 6511 -4620 6545 -4586
rect 6607 -4572 6641 -4538
rect 6890 -4458 6924 -4424
rect 6755 -4632 6789 -4598
rect 6851 -4584 6885 -4550
rect 7168 -4474 7202 -4440
rect 6995 -4610 7029 -4576
rect 7091 -4582 7125 -4548
rect 7291 -4574 7325 -4540
rect 7631 -4574 7665 -4540
rect 7802 -4574 7836 -4540
rect 7904 -4559 7938 -4525
rect 8292 -4458 8326 -4424
rect 8111 -4513 8145 -4479
rect 8541 -4484 8575 -4450
rect 8270 -4620 8304 -4586
rect 8372 -4626 8406 -4592
rect 8627 -4620 8661 -4586
rect 8723 -4572 8757 -4538
rect 9006 -4458 9040 -4424
rect 8871 -4632 8905 -4598
rect 8967 -4584 9001 -4550
rect 9284 -4474 9318 -4440
rect 9111 -4610 9145 -4576
rect 9207 -4582 9241 -4548
rect 9407 -4574 9441 -4540
rect 9747 -4574 9781 -4540
rect 9918 -4574 9952 -4540
rect 10020 -4559 10054 -4525
rect 10408 -4458 10442 -4424
rect 10227 -4513 10261 -4479
rect 10657 -4484 10691 -4450
rect 10386 -4620 10420 -4586
rect 10488 -4626 10522 -4592
rect 10743 -4620 10777 -4586
rect 10839 -4572 10873 -4538
rect 11122 -4458 11156 -4424
rect 10987 -4632 11021 -4598
rect 11083 -4584 11117 -4550
rect 11400 -4474 11434 -4440
rect 11227 -4610 11261 -4576
rect 11323 -4582 11357 -4548
rect 11523 -4574 11557 -4540
rect 11863 -4574 11897 -4540
rect 12034 -4574 12068 -4540
rect 12136 -4559 12170 -4525
rect 12524 -4458 12558 -4424
rect 12343 -4513 12377 -4479
rect 12773 -4484 12807 -4450
rect 12502 -4620 12536 -4586
rect 12604 -4626 12638 -4592
rect 12859 -4620 12893 -4586
rect 12955 -4572 12989 -4538
rect 13238 -4458 13272 -4424
rect 13103 -4632 13137 -4598
rect 13199 -4584 13233 -4550
rect 13516 -4474 13550 -4440
rect 13343 -4610 13377 -4576
rect 13439 -4582 13473 -4548
rect 13639 -4574 13673 -4540
rect 13979 -4574 14013 -4540
rect 14150 -4574 14184 -4540
rect 14252 -4559 14286 -4525
rect 14640 -4458 14674 -4424
rect 14459 -4513 14493 -4479
rect 14889 -4484 14923 -4450
rect 14618 -4620 14652 -4586
rect 14720 -4626 14754 -4592
rect 14975 -4620 15009 -4586
rect 15071 -4572 15105 -4538
rect 15354 -4458 15388 -4424
rect 15219 -4632 15253 -4598
rect 15315 -4584 15349 -4550
rect 15632 -4474 15666 -4440
rect 15459 -4610 15493 -4576
rect 15555 -4582 15589 -4548
rect 15755 -4574 15789 -4540
rect 16095 -4574 16129 -4540
rect 16266 -4574 16300 -4540
rect 16368 -4559 16402 -4525
rect 16756 -4458 16790 -4424
rect 16575 -4513 16609 -4479
rect 17005 -4484 17039 -4450
rect 16734 -4620 16768 -4586
rect 16836 -4626 16870 -4592
rect 17091 -4620 17125 -4586
rect 17187 -4572 17221 -4538
rect 17470 -4458 17504 -4424
rect 17335 -4632 17369 -4598
rect 17431 -4584 17465 -4550
rect 17748 -4474 17782 -4440
rect 17575 -4610 17609 -4576
rect 17671 -4582 17705 -4548
rect 17871 -4574 17905 -4540
rect 18211 -4574 18245 -4540
rect 18382 -4574 18416 -4540
rect 18484 -4559 18518 -4525
rect 18872 -4458 18906 -4424
rect 18691 -4513 18725 -4479
rect 19121 -4484 19155 -4450
rect 18850 -4620 18884 -4586
rect 18952 -4626 18986 -4592
rect 19207 -4620 19241 -4586
rect 19303 -4572 19337 -4538
rect 19586 -4458 19620 -4424
rect 19451 -4632 19485 -4598
rect 19547 -4584 19581 -4550
rect 19864 -4474 19898 -4440
rect 19691 -4610 19725 -4576
rect 19787 -4582 19821 -4548
rect 19987 -4574 20021 -4540
rect 20327 -4574 20361 -4540
rect 20498 -4574 20532 -4540
rect 20600 -4559 20634 -4525
rect 20988 -4458 21022 -4424
rect 20807 -4513 20841 -4479
rect 21237 -4484 21271 -4450
rect 20966 -4620 21000 -4586
rect 21068 -4626 21102 -4592
rect 21323 -4620 21357 -4586
rect 21419 -4572 21453 -4538
rect 21702 -4458 21736 -4424
rect 21567 -4632 21601 -4598
rect 21663 -4584 21697 -4550
rect 21980 -4474 22014 -4440
rect 21807 -4610 21841 -4576
rect 21903 -4582 21937 -4548
rect 22103 -4574 22137 -4540
rect 22443 -4574 22477 -4540
rect 22614 -4574 22648 -4540
rect 22716 -4559 22750 -4525
rect 23104 -4458 23138 -4424
rect 22923 -4513 22957 -4479
rect 23353 -4484 23387 -4450
rect 23082 -4620 23116 -4586
rect 23184 -4626 23218 -4592
rect 23439 -4620 23473 -4586
rect 23535 -4572 23569 -4538
rect 23818 -4458 23852 -4424
rect 23683 -4632 23717 -4598
rect 23779 -4584 23813 -4550
rect 24096 -4474 24130 -4440
rect 23923 -4610 23957 -4576
rect 24019 -4582 24053 -4548
rect 24219 -4574 24253 -4540
rect 24559 -4574 24593 -4540
rect 24730 -4574 24764 -4540
rect 24832 -4559 24866 -4525
rect 25220 -4458 25254 -4424
rect 25039 -4513 25073 -4479
rect 25469 -4484 25503 -4450
rect 25198 -4620 25232 -4586
rect 25300 -4626 25334 -4592
rect 25555 -4620 25589 -4586
rect 25651 -4572 25685 -4538
rect 25934 -4458 25968 -4424
rect 25799 -4632 25833 -4598
rect 25895 -4584 25929 -4550
rect 26212 -4474 26246 -4440
rect 26039 -4610 26073 -4576
rect 26135 -4582 26169 -4548
rect 26335 -4574 26369 -4540
rect 26675 -4574 26709 -4540
rect 26846 -4574 26880 -4540
rect 26948 -4559 26982 -4525
rect 27336 -4458 27370 -4424
rect 27155 -4513 27189 -4479
rect 27585 -4484 27619 -4450
rect 27314 -4620 27348 -4586
rect 27416 -4626 27450 -4592
rect 27671 -4620 27705 -4586
rect 27767 -4572 27801 -4538
rect 28050 -4458 28084 -4424
rect 27915 -4632 27949 -4598
rect 28011 -4584 28045 -4550
rect 28328 -4474 28362 -4440
rect 28155 -4610 28189 -4576
rect 28251 -4582 28285 -4548
rect 28451 -4574 28485 -4540
rect 28791 -4574 28825 -4540
rect 28962 -4574 28996 -4540
rect 29064 -4559 29098 -4525
rect 29452 -4458 29486 -4424
rect 29271 -4513 29305 -4479
rect 29701 -4484 29735 -4450
rect 29430 -4620 29464 -4586
rect 29532 -4626 29566 -4592
rect 29787 -4620 29821 -4586
rect 29883 -4572 29917 -4538
rect 30166 -4458 30200 -4424
rect 30031 -4632 30065 -4598
rect 30127 -4584 30161 -4550
rect 30444 -4474 30478 -4440
rect 30271 -4610 30305 -4576
rect 30367 -4582 30401 -4548
rect 30567 -4574 30601 -4540
rect 30907 -4574 30941 -4540
rect 31078 -4574 31112 -4540
rect 31180 -4559 31214 -4525
rect 31568 -4458 31602 -4424
rect 31387 -4513 31421 -4479
rect 31817 -4484 31851 -4450
rect 31546 -4620 31580 -4586
rect 31648 -4626 31682 -4592
rect 31903 -4620 31937 -4586
rect 31999 -4572 32033 -4538
rect 32282 -4458 32316 -4424
rect 32147 -4632 32181 -4598
rect 32243 -4584 32277 -4550
rect 32560 -4474 32594 -4440
rect 32387 -4610 32421 -4576
rect 32483 -4582 32517 -4548
rect 32683 -4574 32717 -4540
rect 33023 -4574 33057 -4540
rect 4431 -7585 5796 -7551
rect 6290 -7585 7657 -7551
rect 4431 -9095 5796 -9061
rect 6290 -9095 7657 -9061
rect 4431 -10605 5796 -10571
rect 6290 -10605 7657 -10571
rect 4431 -12115 5796 -12081
rect 6290 -12115 7657 -12081
rect 4431 -13625 5796 -13591
rect 6290 -13625 7657 -13591
rect 4431 -15135 5796 -15101
rect 6290 -15135 7657 -15101
rect 4431 -16645 5796 -16611
rect 6290 -16645 7657 -16611
rect 4431 -18155 5796 -18121
rect 6290 -18155 7657 -18121
rect 4431 -19665 5796 -19631
rect 6290 -19665 7657 -19631
rect 4431 -21175 5796 -21141
rect 6290 -21175 7657 -21141
rect 4431 -22685 5796 -22651
rect 6290 -22685 7657 -22651
rect 4431 -24195 5796 -24161
rect 6290 -24195 7657 -24161
rect 4431 -25705 5796 -25671
rect 6290 -25705 7657 -25671
rect 9516 -7628 9550 -7594
rect 10176 -7628 10210 -7594
rect 10646 -7628 10680 -7594
rect 11249 -7629 11283 -7595
rect 11507 -7629 11541 -7595
rect 11765 -7629 11799 -7595
rect 12023 -7629 12057 -7595
rect 12281 -7629 12315 -7595
rect 13064 -7629 13098 -7595
rect 13322 -7629 13356 -7595
rect 13580 -7629 13614 -7595
rect 13838 -7629 13872 -7595
rect 14096 -7629 14130 -7595
rect 14870 -7629 14904 -7595
rect 15128 -7629 15162 -7595
rect 15386 -7629 15420 -7595
rect 15644 -7629 15678 -7595
rect 15902 -7629 15936 -7595
rect 9516 -7956 9550 -7922
rect 10176 -7956 10210 -7922
rect 10646 -7956 10680 -7922
rect 11249 -7957 11283 -7923
rect 11507 -7957 11541 -7923
rect 11765 -7957 11799 -7923
rect 12023 -7957 12057 -7923
rect 12281 -7957 12315 -7923
rect 13064 -7957 13098 -7923
rect 13322 -7957 13356 -7923
rect 13580 -7957 13614 -7923
rect 13838 -7957 13872 -7923
rect 14096 -7957 14130 -7923
rect 14870 -7957 14904 -7923
rect 15128 -7957 15162 -7923
rect 15386 -7957 15420 -7923
rect 15644 -7957 15678 -7923
rect 15902 -7957 15936 -7923
rect 9408 -8599 9474 -8561
rect 10060 -8602 10214 -8568
rect 10794 -8599 10860 -8561
rect 11164 -8599 11230 -8561
rect 11586 -8599 11652 -8561
rect 12008 -8599 12074 -8561
rect 12730 -8602 12884 -8568
rect 13508 -8599 13574 -8561
rect 13878 -8599 13944 -8561
rect 14300 -8599 14366 -8561
rect 14722 -8599 14788 -8561
rect 15393 -8601 15547 -8567
rect 16162 -8599 16228 -8561
rect 10060 -8840 10214 -8806
rect 12730 -8840 12884 -8806
rect 15393 -8839 15547 -8805
rect 9242 -9598 9276 -9564
rect 9500 -9598 9534 -9564
rect 9758 -9598 9792 -9564
rect 10016 -9598 10050 -9564
rect 10274 -9598 10308 -9564
rect 10532 -9598 10566 -9564
rect 10790 -9598 10824 -9564
rect 11048 -9598 11082 -9564
rect 11912 -9598 11946 -9564
rect 12170 -9598 12204 -9564
rect 12428 -9598 12462 -9564
rect 12686 -9598 12720 -9564
rect 12944 -9598 12978 -9564
rect 13202 -9598 13236 -9564
rect 13460 -9598 13494 -9564
rect 13718 -9598 13752 -9564
rect 14575 -9597 14609 -9563
rect 14833 -9597 14867 -9563
rect 15091 -9597 15125 -9563
rect 15349 -9597 15383 -9563
rect 15607 -9597 15641 -9563
rect 15865 -9597 15899 -9563
rect 16123 -9597 16157 -9563
rect 16381 -9597 16415 -9563
rect 9242 -9908 9276 -9874
rect 9500 -9908 9534 -9874
rect 9758 -9908 9792 -9874
rect 10016 -9908 10050 -9874
rect 10274 -9908 10308 -9874
rect 10532 -9908 10566 -9874
rect 10790 -9908 10824 -9874
rect 11048 -9908 11082 -9874
rect 11912 -9908 11946 -9874
rect 12170 -9908 12204 -9874
rect 12428 -9908 12462 -9874
rect 12686 -9908 12720 -9874
rect 12944 -9908 12978 -9874
rect 13202 -9908 13236 -9874
rect 13460 -9908 13494 -9874
rect 13718 -9908 13752 -9874
rect 14575 -9907 14609 -9873
rect 14833 -9907 14867 -9873
rect 15091 -9907 15125 -9873
rect 15349 -9907 15383 -9873
rect 15607 -9907 15641 -9873
rect 15865 -9907 15899 -9873
rect 16123 -9907 16157 -9873
rect 16381 -9907 16415 -9873
rect 9242 -10016 9276 -9982
rect 9500 -10016 9534 -9982
rect 9758 -10016 9792 -9982
rect 10016 -10016 10050 -9982
rect 10274 -10016 10308 -9982
rect 10532 -10016 10566 -9982
rect 10790 -10016 10824 -9982
rect 11048 -10016 11082 -9982
rect 11912 -10016 11946 -9982
rect 12170 -10016 12204 -9982
rect 12428 -10016 12462 -9982
rect 12686 -10016 12720 -9982
rect 12944 -10016 12978 -9982
rect 13202 -10016 13236 -9982
rect 13460 -10016 13494 -9982
rect 13718 -10016 13752 -9982
rect 14575 -10015 14609 -9981
rect 14833 -10015 14867 -9981
rect 15091 -10015 15125 -9981
rect 15349 -10015 15383 -9981
rect 15607 -10015 15641 -9981
rect 15865 -10015 15899 -9981
rect 16123 -10015 16157 -9981
rect 16381 -10015 16415 -9981
rect 9242 -10326 9276 -10292
rect 9500 -10326 9534 -10292
rect 9758 -10326 9792 -10292
rect 10016 -10326 10050 -10292
rect 10274 -10326 10308 -10292
rect 10532 -10326 10566 -10292
rect 10790 -10326 10824 -10292
rect 11048 -10326 11082 -10292
rect 11912 -10326 11946 -10292
rect 12170 -10326 12204 -10292
rect 12428 -10326 12462 -10292
rect 12686 -10326 12720 -10292
rect 12944 -10326 12978 -10292
rect 13202 -10326 13236 -10292
rect 13460 -10326 13494 -10292
rect 13718 -10326 13752 -10292
rect 14575 -10325 14609 -10291
rect 14833 -10325 14867 -10291
rect 15091 -10325 15125 -10291
rect 15349 -10325 15383 -10291
rect 15607 -10325 15641 -10291
rect 15865 -10325 15899 -10291
rect 16123 -10325 16157 -10291
rect 16381 -10325 16415 -10291
rect 9242 -10434 9276 -10400
rect 9500 -10434 9534 -10400
rect 9758 -10434 9792 -10400
rect 10016 -10434 10050 -10400
rect 10274 -10434 10308 -10400
rect 10532 -10434 10566 -10400
rect 10790 -10434 10824 -10400
rect 11048 -10434 11082 -10400
rect 11912 -10434 11946 -10400
rect 12170 -10434 12204 -10400
rect 12428 -10434 12462 -10400
rect 12686 -10434 12720 -10400
rect 12944 -10434 12978 -10400
rect 13202 -10434 13236 -10400
rect 13460 -10434 13494 -10400
rect 13718 -10434 13752 -10400
rect 14575 -10433 14609 -10399
rect 14833 -10433 14867 -10399
rect 15091 -10433 15125 -10399
rect 15349 -10433 15383 -10399
rect 15607 -10433 15641 -10399
rect 15865 -10433 15899 -10399
rect 16123 -10433 16157 -10399
rect 16381 -10433 16415 -10399
rect 9242 -10744 9276 -10710
rect 9500 -10744 9534 -10710
rect 9758 -10744 9792 -10710
rect 10016 -10744 10050 -10710
rect 10274 -10744 10308 -10710
rect 10532 -10744 10566 -10710
rect 10790 -10744 10824 -10710
rect 11048 -10744 11082 -10710
rect 11912 -10744 11946 -10710
rect 12170 -10744 12204 -10710
rect 12428 -10744 12462 -10710
rect 12686 -10744 12720 -10710
rect 12944 -10744 12978 -10710
rect 13202 -10744 13236 -10710
rect 13460 -10744 13494 -10710
rect 13718 -10744 13752 -10710
rect 14575 -10743 14609 -10709
rect 14833 -10743 14867 -10709
rect 15091 -10743 15125 -10709
rect 15349 -10743 15383 -10709
rect 15607 -10743 15641 -10709
rect 15865 -10743 15899 -10709
rect 16123 -10743 16157 -10709
rect 16381 -10743 16415 -10709
rect 9242 -10852 9276 -10818
rect 9500 -10852 9534 -10818
rect 9758 -10852 9792 -10818
rect 10016 -10852 10050 -10818
rect 10274 -10852 10308 -10818
rect 10532 -10852 10566 -10818
rect 10790 -10852 10824 -10818
rect 11048 -10852 11082 -10818
rect 11912 -10852 11946 -10818
rect 12170 -10852 12204 -10818
rect 12428 -10852 12462 -10818
rect 12686 -10852 12720 -10818
rect 12944 -10852 12978 -10818
rect 13202 -10852 13236 -10818
rect 13460 -10852 13494 -10818
rect 13718 -10852 13752 -10818
rect 14575 -10851 14609 -10817
rect 14833 -10851 14867 -10817
rect 15091 -10851 15125 -10817
rect 15349 -10851 15383 -10817
rect 15607 -10851 15641 -10817
rect 15865 -10851 15899 -10817
rect 16123 -10851 16157 -10817
rect 16381 -10851 16415 -10817
rect 9242 -11162 9276 -11128
rect 9500 -11162 9534 -11128
rect 9758 -11162 9792 -11128
rect 10016 -11162 10050 -11128
rect 10274 -11162 10308 -11128
rect 10532 -11162 10566 -11128
rect 10790 -11162 10824 -11128
rect 11048 -11162 11082 -11128
rect 11912 -11162 11946 -11128
rect 12170 -11162 12204 -11128
rect 12428 -11162 12462 -11128
rect 12686 -11162 12720 -11128
rect 12944 -11162 12978 -11128
rect 13202 -11162 13236 -11128
rect 13460 -11162 13494 -11128
rect 13718 -11162 13752 -11128
rect 14575 -11161 14609 -11127
rect 14833 -11161 14867 -11127
rect 15091 -11161 15125 -11127
rect 15349 -11161 15383 -11127
rect 15607 -11161 15641 -11127
rect 15865 -11161 15899 -11127
rect 16123 -11161 16157 -11127
rect 16381 -11161 16415 -11127
rect 9242 -11270 9276 -11236
rect 9500 -11270 9534 -11236
rect 9758 -11270 9792 -11236
rect 10016 -11270 10050 -11236
rect 10274 -11270 10308 -11236
rect 10532 -11270 10566 -11236
rect 10790 -11270 10824 -11236
rect 11048 -11270 11082 -11236
rect 11912 -11270 11946 -11236
rect 12170 -11270 12204 -11236
rect 12428 -11270 12462 -11236
rect 12686 -11270 12720 -11236
rect 12944 -11270 12978 -11236
rect 13202 -11270 13236 -11236
rect 13460 -11270 13494 -11236
rect 13718 -11270 13752 -11236
rect 14575 -11269 14609 -11235
rect 14833 -11269 14867 -11235
rect 15091 -11269 15125 -11235
rect 15349 -11269 15383 -11235
rect 15607 -11269 15641 -11235
rect 15865 -11269 15899 -11235
rect 16123 -11269 16157 -11235
rect 16381 -11269 16415 -11235
rect 9242 -11580 9276 -11546
rect 9500 -11580 9534 -11546
rect 9758 -11580 9792 -11546
rect 10016 -11580 10050 -11546
rect 10274 -11580 10308 -11546
rect 10532 -11580 10566 -11546
rect 10790 -11580 10824 -11546
rect 11048 -11580 11082 -11546
rect 11912 -11580 11946 -11546
rect 12170 -11580 12204 -11546
rect 12428 -11580 12462 -11546
rect 12686 -11580 12720 -11546
rect 12944 -11580 12978 -11546
rect 13202 -11580 13236 -11546
rect 13460 -11580 13494 -11546
rect 13718 -11580 13752 -11546
rect 14575 -11579 14609 -11545
rect 14833 -11579 14867 -11545
rect 15091 -11579 15125 -11545
rect 15349 -11579 15383 -11545
rect 15607 -11579 15641 -11545
rect 15865 -11579 15899 -11545
rect 16123 -11579 16157 -11545
rect 16381 -11579 16415 -11545
rect 9242 -11688 9276 -11654
rect 9500 -11688 9534 -11654
rect 9758 -11688 9792 -11654
rect 10016 -11688 10050 -11654
rect 10274 -11688 10308 -11654
rect 10532 -11688 10566 -11654
rect 10790 -11688 10824 -11654
rect 11048 -11688 11082 -11654
rect 11912 -11688 11946 -11654
rect 12170 -11688 12204 -11654
rect 12428 -11688 12462 -11654
rect 12686 -11688 12720 -11654
rect 12944 -11688 12978 -11654
rect 13202 -11688 13236 -11654
rect 13460 -11688 13494 -11654
rect 13718 -11688 13752 -11654
rect 14575 -11687 14609 -11653
rect 14833 -11687 14867 -11653
rect 15091 -11687 15125 -11653
rect 15349 -11687 15383 -11653
rect 15607 -11687 15641 -11653
rect 15865 -11687 15899 -11653
rect 16123 -11687 16157 -11653
rect 16381 -11687 16415 -11653
rect 9242 -11998 9276 -11964
rect 9500 -11998 9534 -11964
rect 9758 -11998 9792 -11964
rect 10016 -11998 10050 -11964
rect 10274 -11998 10308 -11964
rect 10532 -11998 10566 -11964
rect 10790 -11998 10824 -11964
rect 11048 -11998 11082 -11964
rect 11912 -11998 11946 -11964
rect 12170 -11998 12204 -11964
rect 12428 -11998 12462 -11964
rect 12686 -11998 12720 -11964
rect 12944 -11998 12978 -11964
rect 13202 -11998 13236 -11964
rect 13460 -11998 13494 -11964
rect 13718 -11998 13752 -11964
rect 14575 -11997 14609 -11963
rect 14833 -11997 14867 -11963
rect 15091 -11997 15125 -11963
rect 15349 -11997 15383 -11963
rect 15607 -11997 15641 -11963
rect 15865 -11997 15899 -11963
rect 16123 -11997 16157 -11963
rect 16381 -11997 16415 -11963
rect 9242 -12106 9276 -12072
rect 9500 -12106 9534 -12072
rect 9758 -12106 9792 -12072
rect 10016 -12106 10050 -12072
rect 10274 -12106 10308 -12072
rect 10532 -12106 10566 -12072
rect 10790 -12106 10824 -12072
rect 11048 -12106 11082 -12072
rect 11912 -12106 11946 -12072
rect 12170 -12106 12204 -12072
rect 12428 -12106 12462 -12072
rect 12686 -12106 12720 -12072
rect 12944 -12106 12978 -12072
rect 13202 -12106 13236 -12072
rect 13460 -12106 13494 -12072
rect 13718 -12106 13752 -12072
rect 14575 -12105 14609 -12071
rect 14833 -12105 14867 -12071
rect 15091 -12105 15125 -12071
rect 15349 -12105 15383 -12071
rect 15607 -12105 15641 -12071
rect 15865 -12105 15899 -12071
rect 16123 -12105 16157 -12071
rect 16381 -12105 16415 -12071
rect 9242 -12416 9276 -12382
rect 9500 -12416 9534 -12382
rect 9758 -12416 9792 -12382
rect 10016 -12416 10050 -12382
rect 10274 -12416 10308 -12382
rect 10532 -12416 10566 -12382
rect 10790 -12416 10824 -12382
rect 11048 -12416 11082 -12382
rect 11912 -12416 11946 -12382
rect 12170 -12416 12204 -12382
rect 12428 -12416 12462 -12382
rect 12686 -12416 12720 -12382
rect 12944 -12416 12978 -12382
rect 13202 -12416 13236 -12382
rect 13460 -12416 13494 -12382
rect 13718 -12416 13752 -12382
rect 14575 -12415 14609 -12381
rect 14833 -12415 14867 -12381
rect 15091 -12415 15125 -12381
rect 15349 -12415 15383 -12381
rect 15607 -12415 15641 -12381
rect 15865 -12415 15899 -12381
rect 16123 -12415 16157 -12381
rect 16381 -12415 16415 -12381
rect 9122 -12758 9156 -12724
rect 9662 -12758 9696 -12724
rect 10142 -12758 10176 -12724
rect 10645 -12756 10679 -12722
rect 11155 -12746 11189 -12712
rect 11792 -12758 11826 -12724
rect 12332 -12758 12366 -12724
rect 12812 -12758 12846 -12724
rect 13315 -12756 13349 -12722
rect 13825 -12746 13859 -12712
rect 14455 -12757 14489 -12723
rect 9122 -13068 9156 -13034
rect 9662 -13068 9696 -13034
rect 10142 -13068 10176 -13034
rect 10645 -13066 10679 -13032
rect 14995 -12757 15029 -12723
rect 15475 -12757 15509 -12723
rect 15978 -12755 16012 -12721
rect 16488 -12745 16522 -12711
rect 11155 -13056 11189 -13022
rect 11792 -13068 11826 -13034
rect 12332 -13068 12366 -13034
rect 12812 -13068 12846 -13034
rect 13315 -13066 13349 -13032
rect 13825 -13056 13859 -13022
rect 14455 -13067 14489 -13033
rect 14995 -13067 15029 -13033
rect 15475 -13067 15509 -13033
rect 15978 -13065 16012 -13031
rect 16488 -13055 16522 -13021
rect 9408 -14281 9474 -14243
rect 10052 -14284 10206 -14250
rect 10794 -14282 10860 -14244
rect 11164 -14282 11230 -14244
rect 11586 -14282 11652 -14244
rect 12008 -14282 12074 -14244
rect 12729 -14284 12883 -14250
rect 13508 -14278 13574 -14240
rect 13878 -14278 13944 -14240
rect 14300 -14278 14366 -14240
rect 14722 -14278 14788 -14240
rect 15393 -14283 15547 -14249
rect 16106 -14281 16172 -14243
rect 10052 -14522 10206 -14488
rect 12729 -14522 12883 -14488
rect 15393 -14521 15547 -14487
rect 9242 -15315 9276 -15281
rect 9500 -15315 9534 -15281
rect 9758 -15315 9792 -15281
rect 10016 -15315 10050 -15281
rect 10274 -15315 10308 -15281
rect 10532 -15315 10566 -15281
rect 10790 -15315 10824 -15281
rect 11048 -15315 11082 -15281
rect 11912 -15315 11946 -15281
rect 12170 -15315 12204 -15281
rect 12428 -15315 12462 -15281
rect 12686 -15315 12720 -15281
rect 12944 -15315 12978 -15281
rect 13202 -15315 13236 -15281
rect 13460 -15315 13494 -15281
rect 13718 -15315 13752 -15281
rect 14575 -15314 14609 -15280
rect 14833 -15314 14867 -15280
rect 15091 -15314 15125 -15280
rect 15349 -15314 15383 -15280
rect 15607 -15314 15641 -15280
rect 15865 -15314 15899 -15280
rect 16123 -15314 16157 -15280
rect 16381 -15314 16415 -15280
rect 9242 -15625 9276 -15591
rect 9500 -15625 9534 -15591
rect 9758 -15625 9792 -15591
rect 10016 -15625 10050 -15591
rect 10274 -15625 10308 -15591
rect 10532 -15625 10566 -15591
rect 10790 -15625 10824 -15591
rect 11048 -15625 11082 -15591
rect 11912 -15625 11946 -15591
rect 12170 -15625 12204 -15591
rect 12428 -15625 12462 -15591
rect 12686 -15625 12720 -15591
rect 12944 -15625 12978 -15591
rect 13202 -15625 13236 -15591
rect 13460 -15625 13494 -15591
rect 13718 -15625 13752 -15591
rect 14575 -15624 14609 -15590
rect 14833 -15624 14867 -15590
rect 15091 -15624 15125 -15590
rect 15349 -15624 15383 -15590
rect 15607 -15624 15641 -15590
rect 15865 -15624 15899 -15590
rect 16123 -15624 16157 -15590
rect 16381 -15624 16415 -15590
rect 9242 -15733 9276 -15699
rect 9500 -15733 9534 -15699
rect 9758 -15733 9792 -15699
rect 10016 -15733 10050 -15699
rect 10274 -15733 10308 -15699
rect 10532 -15733 10566 -15699
rect 10790 -15733 10824 -15699
rect 11048 -15733 11082 -15699
rect 11912 -15733 11946 -15699
rect 12170 -15733 12204 -15699
rect 12428 -15733 12462 -15699
rect 12686 -15733 12720 -15699
rect 12944 -15733 12978 -15699
rect 13202 -15733 13236 -15699
rect 13460 -15733 13494 -15699
rect 13718 -15733 13752 -15699
rect 14575 -15732 14609 -15698
rect 14833 -15732 14867 -15698
rect 15091 -15732 15125 -15698
rect 15349 -15732 15383 -15698
rect 15607 -15732 15641 -15698
rect 15865 -15732 15899 -15698
rect 16123 -15732 16157 -15698
rect 16381 -15732 16415 -15698
rect 9242 -16043 9276 -16009
rect 9500 -16043 9534 -16009
rect 9758 -16043 9792 -16009
rect 10016 -16043 10050 -16009
rect 10274 -16043 10308 -16009
rect 10532 -16043 10566 -16009
rect 10790 -16043 10824 -16009
rect 11048 -16043 11082 -16009
rect 11912 -16043 11946 -16009
rect 12170 -16043 12204 -16009
rect 12428 -16043 12462 -16009
rect 12686 -16043 12720 -16009
rect 12944 -16043 12978 -16009
rect 13202 -16043 13236 -16009
rect 13460 -16043 13494 -16009
rect 13718 -16043 13752 -16009
rect 14575 -16042 14609 -16008
rect 14833 -16042 14867 -16008
rect 15091 -16042 15125 -16008
rect 15349 -16042 15383 -16008
rect 15607 -16042 15641 -16008
rect 15865 -16042 15899 -16008
rect 16123 -16042 16157 -16008
rect 16381 -16042 16415 -16008
rect 9242 -16151 9276 -16117
rect 9500 -16151 9534 -16117
rect 9758 -16151 9792 -16117
rect 10016 -16151 10050 -16117
rect 10274 -16151 10308 -16117
rect 10532 -16151 10566 -16117
rect 10790 -16151 10824 -16117
rect 11048 -16151 11082 -16117
rect 11912 -16151 11946 -16117
rect 12170 -16151 12204 -16117
rect 12428 -16151 12462 -16117
rect 12686 -16151 12720 -16117
rect 12944 -16151 12978 -16117
rect 13202 -16151 13236 -16117
rect 13460 -16151 13494 -16117
rect 13718 -16151 13752 -16117
rect 14575 -16150 14609 -16116
rect 14833 -16150 14867 -16116
rect 15091 -16150 15125 -16116
rect 15349 -16150 15383 -16116
rect 15607 -16150 15641 -16116
rect 15865 -16150 15899 -16116
rect 16123 -16150 16157 -16116
rect 16381 -16150 16415 -16116
rect 9242 -16461 9276 -16427
rect 9500 -16461 9534 -16427
rect 9758 -16461 9792 -16427
rect 10016 -16461 10050 -16427
rect 10274 -16461 10308 -16427
rect 10532 -16461 10566 -16427
rect 10790 -16461 10824 -16427
rect 11048 -16461 11082 -16427
rect 11912 -16461 11946 -16427
rect 12170 -16461 12204 -16427
rect 12428 -16461 12462 -16427
rect 12686 -16461 12720 -16427
rect 12944 -16461 12978 -16427
rect 13202 -16461 13236 -16427
rect 13460 -16461 13494 -16427
rect 13718 -16461 13752 -16427
rect 14575 -16460 14609 -16426
rect 14833 -16460 14867 -16426
rect 15091 -16460 15125 -16426
rect 15349 -16460 15383 -16426
rect 15607 -16460 15641 -16426
rect 15865 -16460 15899 -16426
rect 16123 -16460 16157 -16426
rect 16381 -16460 16415 -16426
rect 9242 -16569 9276 -16535
rect 9500 -16569 9534 -16535
rect 9758 -16569 9792 -16535
rect 10016 -16569 10050 -16535
rect 10274 -16569 10308 -16535
rect 10532 -16569 10566 -16535
rect 10790 -16569 10824 -16535
rect 11048 -16569 11082 -16535
rect 11912 -16569 11946 -16535
rect 12170 -16569 12204 -16535
rect 12428 -16569 12462 -16535
rect 12686 -16569 12720 -16535
rect 12944 -16569 12978 -16535
rect 13202 -16569 13236 -16535
rect 13460 -16569 13494 -16535
rect 13718 -16569 13752 -16535
rect 14575 -16568 14609 -16534
rect 14833 -16568 14867 -16534
rect 15091 -16568 15125 -16534
rect 15349 -16568 15383 -16534
rect 15607 -16568 15641 -16534
rect 15865 -16568 15899 -16534
rect 16123 -16568 16157 -16534
rect 16381 -16568 16415 -16534
rect 9242 -16879 9276 -16845
rect 9500 -16879 9534 -16845
rect 9758 -16879 9792 -16845
rect 10016 -16879 10050 -16845
rect 10274 -16879 10308 -16845
rect 10532 -16879 10566 -16845
rect 10790 -16879 10824 -16845
rect 11048 -16879 11082 -16845
rect 11912 -16879 11946 -16845
rect 12170 -16879 12204 -16845
rect 12428 -16879 12462 -16845
rect 12686 -16879 12720 -16845
rect 12944 -16879 12978 -16845
rect 13202 -16879 13236 -16845
rect 13460 -16879 13494 -16845
rect 13718 -16879 13752 -16845
rect 14575 -16878 14609 -16844
rect 14833 -16878 14867 -16844
rect 15091 -16878 15125 -16844
rect 15349 -16878 15383 -16844
rect 15607 -16878 15641 -16844
rect 15865 -16878 15899 -16844
rect 16123 -16878 16157 -16844
rect 16381 -16878 16415 -16844
rect 9242 -16987 9276 -16953
rect 9500 -16987 9534 -16953
rect 9758 -16987 9792 -16953
rect 10016 -16987 10050 -16953
rect 10274 -16987 10308 -16953
rect 10532 -16987 10566 -16953
rect 10790 -16987 10824 -16953
rect 11048 -16987 11082 -16953
rect 11912 -16987 11946 -16953
rect 12170 -16987 12204 -16953
rect 12428 -16987 12462 -16953
rect 12686 -16987 12720 -16953
rect 12944 -16987 12978 -16953
rect 13202 -16987 13236 -16953
rect 13460 -16987 13494 -16953
rect 13718 -16987 13752 -16953
rect 14575 -16986 14609 -16952
rect 14833 -16986 14867 -16952
rect 15091 -16986 15125 -16952
rect 15349 -16986 15383 -16952
rect 15607 -16986 15641 -16952
rect 15865 -16986 15899 -16952
rect 16123 -16986 16157 -16952
rect 16381 -16986 16415 -16952
rect 9242 -17297 9276 -17263
rect 9500 -17297 9534 -17263
rect 9758 -17297 9792 -17263
rect 10016 -17297 10050 -17263
rect 10274 -17297 10308 -17263
rect 10532 -17297 10566 -17263
rect 10790 -17297 10824 -17263
rect 11048 -17297 11082 -17263
rect 11912 -17297 11946 -17263
rect 12170 -17297 12204 -17263
rect 12428 -17297 12462 -17263
rect 12686 -17297 12720 -17263
rect 12944 -17297 12978 -17263
rect 13202 -17297 13236 -17263
rect 13460 -17297 13494 -17263
rect 13718 -17297 13752 -17263
rect 14575 -17296 14609 -17262
rect 14833 -17296 14867 -17262
rect 15091 -17296 15125 -17262
rect 15349 -17296 15383 -17262
rect 15607 -17296 15641 -17262
rect 15865 -17296 15899 -17262
rect 16123 -17296 16157 -17262
rect 16381 -17296 16415 -17262
rect 9242 -17405 9276 -17371
rect 9500 -17405 9534 -17371
rect 9758 -17405 9792 -17371
rect 10016 -17405 10050 -17371
rect 10274 -17405 10308 -17371
rect 10532 -17405 10566 -17371
rect 10790 -17405 10824 -17371
rect 11048 -17405 11082 -17371
rect 11912 -17405 11946 -17371
rect 12170 -17405 12204 -17371
rect 12428 -17405 12462 -17371
rect 12686 -17405 12720 -17371
rect 12944 -17405 12978 -17371
rect 13202 -17405 13236 -17371
rect 13460 -17405 13494 -17371
rect 13718 -17405 13752 -17371
rect 14575 -17404 14609 -17370
rect 14833 -17404 14867 -17370
rect 15091 -17404 15125 -17370
rect 15349 -17404 15383 -17370
rect 15607 -17404 15641 -17370
rect 15865 -17404 15899 -17370
rect 16123 -17404 16157 -17370
rect 16381 -17404 16415 -17370
rect 9242 -17715 9276 -17681
rect 9500 -17715 9534 -17681
rect 9758 -17715 9792 -17681
rect 10016 -17715 10050 -17681
rect 10274 -17715 10308 -17681
rect 10532 -17715 10566 -17681
rect 10790 -17715 10824 -17681
rect 11048 -17715 11082 -17681
rect 11912 -17715 11946 -17681
rect 12170 -17715 12204 -17681
rect 12428 -17715 12462 -17681
rect 12686 -17715 12720 -17681
rect 12944 -17715 12978 -17681
rect 13202 -17715 13236 -17681
rect 13460 -17715 13494 -17681
rect 13718 -17715 13752 -17681
rect 14575 -17714 14609 -17680
rect 14833 -17714 14867 -17680
rect 15091 -17714 15125 -17680
rect 15349 -17714 15383 -17680
rect 15607 -17714 15641 -17680
rect 15865 -17714 15899 -17680
rect 16123 -17714 16157 -17680
rect 16381 -17714 16415 -17680
rect 9242 -17823 9276 -17789
rect 9500 -17823 9534 -17789
rect 9758 -17823 9792 -17789
rect 10016 -17823 10050 -17789
rect 10274 -17823 10308 -17789
rect 10532 -17823 10566 -17789
rect 10790 -17823 10824 -17789
rect 11048 -17823 11082 -17789
rect 11912 -17823 11946 -17789
rect 12170 -17823 12204 -17789
rect 12428 -17823 12462 -17789
rect 12686 -17823 12720 -17789
rect 12944 -17823 12978 -17789
rect 13202 -17823 13236 -17789
rect 13460 -17823 13494 -17789
rect 13718 -17823 13752 -17789
rect 14575 -17822 14609 -17788
rect 14833 -17822 14867 -17788
rect 15091 -17822 15125 -17788
rect 15349 -17822 15383 -17788
rect 15607 -17822 15641 -17788
rect 15865 -17822 15899 -17788
rect 16123 -17822 16157 -17788
rect 16381 -17822 16415 -17788
rect 9242 -18133 9276 -18099
rect 9500 -18133 9534 -18099
rect 9758 -18133 9792 -18099
rect 10016 -18133 10050 -18099
rect 10274 -18133 10308 -18099
rect 10532 -18133 10566 -18099
rect 10790 -18133 10824 -18099
rect 11048 -18133 11082 -18099
rect 11912 -18133 11946 -18099
rect 12170 -18133 12204 -18099
rect 12428 -18133 12462 -18099
rect 12686 -18133 12720 -18099
rect 12944 -18133 12978 -18099
rect 13202 -18133 13236 -18099
rect 13460 -18133 13494 -18099
rect 13718 -18133 13752 -18099
rect 14575 -18132 14609 -18098
rect 14833 -18132 14867 -18098
rect 15091 -18132 15125 -18098
rect 15349 -18132 15383 -18098
rect 15607 -18132 15641 -18098
rect 15865 -18132 15899 -18098
rect 16123 -18132 16157 -18098
rect 16381 -18132 16415 -18098
rect 9122 -18475 9156 -18441
rect 9662 -18475 9696 -18441
rect 10142 -18475 10176 -18441
rect 10645 -18473 10679 -18439
rect 11155 -18463 11189 -18429
rect 11792 -18475 11826 -18441
rect 12332 -18475 12366 -18441
rect 12812 -18475 12846 -18441
rect 13315 -18473 13349 -18439
rect 13825 -18463 13859 -18429
rect 14455 -18474 14489 -18440
rect 9122 -18785 9156 -18751
rect 9662 -18785 9696 -18751
rect 10142 -18785 10176 -18751
rect 10645 -18783 10679 -18749
rect 14995 -18474 15029 -18440
rect 15475 -18474 15509 -18440
rect 15978 -18472 16012 -18438
rect 16488 -18462 16522 -18428
rect 11155 -18773 11189 -18739
rect 11792 -18785 11826 -18751
rect 12332 -18785 12366 -18751
rect 12812 -18785 12846 -18751
rect 13315 -18783 13349 -18749
rect 13825 -18773 13859 -18739
rect 14455 -18784 14489 -18750
rect 14995 -18784 15029 -18750
rect 15475 -18784 15509 -18750
rect 15978 -18782 16012 -18748
rect 16488 -18772 16522 -18738
rect 16698 -19575 16732 -19541
rect 9453 -20205 9519 -20167
rect 10060 -20209 10214 -20175
rect 10794 -20207 10860 -20169
rect 11164 -20207 11230 -20169
rect 11586 -20207 11652 -20169
rect 12008 -20207 12074 -20169
rect 12730 -20209 12884 -20175
rect 13495 -20207 13561 -20169
rect 13865 -20207 13931 -20169
rect 14287 -20207 14353 -20169
rect 14709 -20207 14775 -20169
rect 15393 -20208 15547 -20174
rect 10060 -20447 10214 -20413
rect 12730 -20447 12884 -20413
rect 15393 -20446 15547 -20412
rect 17088 -19577 17122 -19543
rect 16698 -20039 16732 -20005
rect 17088 -20041 17122 -20007
rect 16702 -20371 16736 -20337
rect 17092 -20371 17126 -20337
rect 16702 -20565 16736 -20531
rect 17092 -20565 17126 -20531
rect 9242 -21219 9276 -21185
rect 9500 -21219 9534 -21185
rect 9758 -21219 9792 -21185
rect 10016 -21219 10050 -21185
rect 10274 -21219 10308 -21185
rect 10532 -21219 10566 -21185
rect 10790 -21219 10824 -21185
rect 11048 -21219 11082 -21185
rect 11912 -21219 11946 -21185
rect 12170 -21219 12204 -21185
rect 12428 -21219 12462 -21185
rect 12686 -21219 12720 -21185
rect 12944 -21219 12978 -21185
rect 13202 -21219 13236 -21185
rect 13460 -21219 13494 -21185
rect 13718 -21219 13752 -21185
rect 14575 -21218 14609 -21184
rect 14833 -21218 14867 -21184
rect 15091 -21218 15125 -21184
rect 15349 -21218 15383 -21184
rect 15607 -21218 15641 -21184
rect 15865 -21218 15899 -21184
rect 16123 -21218 16157 -21184
rect 16381 -21218 16415 -21184
rect 9242 -21529 9276 -21495
rect 9500 -21529 9534 -21495
rect 9758 -21529 9792 -21495
rect 10016 -21529 10050 -21495
rect 10274 -21529 10308 -21495
rect 10532 -21529 10566 -21495
rect 10790 -21529 10824 -21495
rect 11048 -21529 11082 -21495
rect 11912 -21529 11946 -21495
rect 12170 -21529 12204 -21495
rect 12428 -21529 12462 -21495
rect 12686 -21529 12720 -21495
rect 12944 -21529 12978 -21495
rect 13202 -21529 13236 -21495
rect 13460 -21529 13494 -21495
rect 13718 -21529 13752 -21495
rect 14575 -21528 14609 -21494
rect 14833 -21528 14867 -21494
rect 15091 -21528 15125 -21494
rect 15349 -21528 15383 -21494
rect 15607 -21528 15641 -21494
rect 15865 -21528 15899 -21494
rect 16123 -21528 16157 -21494
rect 16381 -21528 16415 -21494
rect 9242 -21637 9276 -21603
rect 9500 -21637 9534 -21603
rect 9758 -21637 9792 -21603
rect 10016 -21637 10050 -21603
rect 10274 -21637 10308 -21603
rect 10532 -21637 10566 -21603
rect 10790 -21637 10824 -21603
rect 11048 -21637 11082 -21603
rect 11912 -21637 11946 -21603
rect 12170 -21637 12204 -21603
rect 12428 -21637 12462 -21603
rect 12686 -21637 12720 -21603
rect 12944 -21637 12978 -21603
rect 13202 -21637 13236 -21603
rect 13460 -21637 13494 -21603
rect 13718 -21637 13752 -21603
rect 14575 -21636 14609 -21602
rect 14833 -21636 14867 -21602
rect 15091 -21636 15125 -21602
rect 15349 -21636 15383 -21602
rect 15607 -21636 15641 -21602
rect 15865 -21636 15899 -21602
rect 16123 -21636 16157 -21602
rect 16381 -21636 16415 -21602
rect 9242 -21947 9276 -21913
rect 9500 -21947 9534 -21913
rect 9758 -21947 9792 -21913
rect 10016 -21947 10050 -21913
rect 10274 -21947 10308 -21913
rect 10532 -21947 10566 -21913
rect 10790 -21947 10824 -21913
rect 11048 -21947 11082 -21913
rect 11912 -21947 11946 -21913
rect 12170 -21947 12204 -21913
rect 12428 -21947 12462 -21913
rect 12686 -21947 12720 -21913
rect 12944 -21947 12978 -21913
rect 13202 -21947 13236 -21913
rect 13460 -21947 13494 -21913
rect 13718 -21947 13752 -21913
rect 14575 -21946 14609 -21912
rect 14833 -21946 14867 -21912
rect 15091 -21946 15125 -21912
rect 15349 -21946 15383 -21912
rect 15607 -21946 15641 -21912
rect 15865 -21946 15899 -21912
rect 16123 -21946 16157 -21912
rect 16381 -21946 16415 -21912
rect 9242 -22055 9276 -22021
rect 9500 -22055 9534 -22021
rect 9758 -22055 9792 -22021
rect 10016 -22055 10050 -22021
rect 10274 -22055 10308 -22021
rect 10532 -22055 10566 -22021
rect 10790 -22055 10824 -22021
rect 11048 -22055 11082 -22021
rect 11912 -22055 11946 -22021
rect 12170 -22055 12204 -22021
rect 12428 -22055 12462 -22021
rect 12686 -22055 12720 -22021
rect 12944 -22055 12978 -22021
rect 13202 -22055 13236 -22021
rect 13460 -22055 13494 -22021
rect 13718 -22055 13752 -22021
rect 14575 -22054 14609 -22020
rect 14833 -22054 14867 -22020
rect 15091 -22054 15125 -22020
rect 15349 -22054 15383 -22020
rect 15607 -22054 15641 -22020
rect 15865 -22054 15899 -22020
rect 16123 -22054 16157 -22020
rect 16381 -22054 16415 -22020
rect 9242 -22365 9276 -22331
rect 9500 -22365 9534 -22331
rect 9758 -22365 9792 -22331
rect 10016 -22365 10050 -22331
rect 10274 -22365 10308 -22331
rect 10532 -22365 10566 -22331
rect 10790 -22365 10824 -22331
rect 11048 -22365 11082 -22331
rect 11912 -22365 11946 -22331
rect 12170 -22365 12204 -22331
rect 12428 -22365 12462 -22331
rect 12686 -22365 12720 -22331
rect 12944 -22365 12978 -22331
rect 13202 -22365 13236 -22331
rect 13460 -22365 13494 -22331
rect 13718 -22365 13752 -22331
rect 14575 -22364 14609 -22330
rect 14833 -22364 14867 -22330
rect 15091 -22364 15125 -22330
rect 15349 -22364 15383 -22330
rect 15607 -22364 15641 -22330
rect 15865 -22364 15899 -22330
rect 16123 -22364 16157 -22330
rect 16381 -22364 16415 -22330
rect 9242 -22473 9276 -22439
rect 9500 -22473 9534 -22439
rect 9758 -22473 9792 -22439
rect 10016 -22473 10050 -22439
rect 10274 -22473 10308 -22439
rect 10532 -22473 10566 -22439
rect 10790 -22473 10824 -22439
rect 11048 -22473 11082 -22439
rect 11912 -22473 11946 -22439
rect 12170 -22473 12204 -22439
rect 12428 -22473 12462 -22439
rect 12686 -22473 12720 -22439
rect 12944 -22473 12978 -22439
rect 13202 -22473 13236 -22439
rect 13460 -22473 13494 -22439
rect 13718 -22473 13752 -22439
rect 14575 -22472 14609 -22438
rect 14833 -22472 14867 -22438
rect 15091 -22472 15125 -22438
rect 15349 -22472 15383 -22438
rect 15607 -22472 15641 -22438
rect 15865 -22472 15899 -22438
rect 16123 -22472 16157 -22438
rect 16381 -22472 16415 -22438
rect 9242 -22783 9276 -22749
rect 9500 -22783 9534 -22749
rect 9758 -22783 9792 -22749
rect 10016 -22783 10050 -22749
rect 10274 -22783 10308 -22749
rect 10532 -22783 10566 -22749
rect 10790 -22783 10824 -22749
rect 11048 -22783 11082 -22749
rect 11912 -22783 11946 -22749
rect 12170 -22783 12204 -22749
rect 12428 -22783 12462 -22749
rect 12686 -22783 12720 -22749
rect 12944 -22783 12978 -22749
rect 13202 -22783 13236 -22749
rect 13460 -22783 13494 -22749
rect 13718 -22783 13752 -22749
rect 14575 -22782 14609 -22748
rect 14833 -22782 14867 -22748
rect 15091 -22782 15125 -22748
rect 15349 -22782 15383 -22748
rect 15607 -22782 15641 -22748
rect 15865 -22782 15899 -22748
rect 16123 -22782 16157 -22748
rect 16381 -22782 16415 -22748
rect 9242 -22891 9276 -22857
rect 9500 -22891 9534 -22857
rect 9758 -22891 9792 -22857
rect 10016 -22891 10050 -22857
rect 10274 -22891 10308 -22857
rect 10532 -22891 10566 -22857
rect 10790 -22891 10824 -22857
rect 11048 -22891 11082 -22857
rect 11912 -22891 11946 -22857
rect 12170 -22891 12204 -22857
rect 12428 -22891 12462 -22857
rect 12686 -22891 12720 -22857
rect 12944 -22891 12978 -22857
rect 13202 -22891 13236 -22857
rect 13460 -22891 13494 -22857
rect 13718 -22891 13752 -22857
rect 14575 -22890 14609 -22856
rect 14833 -22890 14867 -22856
rect 15091 -22890 15125 -22856
rect 15349 -22890 15383 -22856
rect 15607 -22890 15641 -22856
rect 15865 -22890 15899 -22856
rect 16123 -22890 16157 -22856
rect 16381 -22890 16415 -22856
rect 9242 -23201 9276 -23167
rect 9500 -23201 9534 -23167
rect 9758 -23201 9792 -23167
rect 10016 -23201 10050 -23167
rect 10274 -23201 10308 -23167
rect 10532 -23201 10566 -23167
rect 10790 -23201 10824 -23167
rect 11048 -23201 11082 -23167
rect 11912 -23201 11946 -23167
rect 12170 -23201 12204 -23167
rect 12428 -23201 12462 -23167
rect 12686 -23201 12720 -23167
rect 12944 -23201 12978 -23167
rect 13202 -23201 13236 -23167
rect 13460 -23201 13494 -23167
rect 13718 -23201 13752 -23167
rect 14575 -23200 14609 -23166
rect 14833 -23200 14867 -23166
rect 15091 -23200 15125 -23166
rect 15349 -23200 15383 -23166
rect 15607 -23200 15641 -23166
rect 15865 -23200 15899 -23166
rect 16123 -23200 16157 -23166
rect 16381 -23200 16415 -23166
rect 9242 -23309 9276 -23275
rect 9500 -23309 9534 -23275
rect 9758 -23309 9792 -23275
rect 10016 -23309 10050 -23275
rect 10274 -23309 10308 -23275
rect 10532 -23309 10566 -23275
rect 10790 -23309 10824 -23275
rect 11048 -23309 11082 -23275
rect 11912 -23309 11946 -23275
rect 12170 -23309 12204 -23275
rect 12428 -23309 12462 -23275
rect 12686 -23309 12720 -23275
rect 12944 -23309 12978 -23275
rect 13202 -23309 13236 -23275
rect 13460 -23309 13494 -23275
rect 13718 -23309 13752 -23275
rect 14575 -23308 14609 -23274
rect 14833 -23308 14867 -23274
rect 15091 -23308 15125 -23274
rect 15349 -23308 15383 -23274
rect 15607 -23308 15641 -23274
rect 15865 -23308 15899 -23274
rect 16123 -23308 16157 -23274
rect 16381 -23308 16415 -23274
rect 9242 -23619 9276 -23585
rect 9500 -23619 9534 -23585
rect 9758 -23619 9792 -23585
rect 10016 -23619 10050 -23585
rect 10274 -23619 10308 -23585
rect 10532 -23619 10566 -23585
rect 10790 -23619 10824 -23585
rect 11048 -23619 11082 -23585
rect 11912 -23619 11946 -23585
rect 12170 -23619 12204 -23585
rect 12428 -23619 12462 -23585
rect 12686 -23619 12720 -23585
rect 12944 -23619 12978 -23585
rect 13202 -23619 13236 -23585
rect 13460 -23619 13494 -23585
rect 13718 -23619 13752 -23585
rect 14575 -23618 14609 -23584
rect 14833 -23618 14867 -23584
rect 15091 -23618 15125 -23584
rect 15349 -23618 15383 -23584
rect 15607 -23618 15641 -23584
rect 15865 -23618 15899 -23584
rect 16123 -23618 16157 -23584
rect 16381 -23618 16415 -23584
rect 9242 -23727 9276 -23693
rect 9500 -23727 9534 -23693
rect 9758 -23727 9792 -23693
rect 10016 -23727 10050 -23693
rect 10274 -23727 10308 -23693
rect 10532 -23727 10566 -23693
rect 10790 -23727 10824 -23693
rect 11048 -23727 11082 -23693
rect 11912 -23727 11946 -23693
rect 12170 -23727 12204 -23693
rect 12428 -23727 12462 -23693
rect 12686 -23727 12720 -23693
rect 12944 -23727 12978 -23693
rect 13202 -23727 13236 -23693
rect 13460 -23727 13494 -23693
rect 13718 -23727 13752 -23693
rect 14575 -23726 14609 -23692
rect 14833 -23726 14867 -23692
rect 15091 -23726 15125 -23692
rect 15349 -23726 15383 -23692
rect 15607 -23726 15641 -23692
rect 15865 -23726 15899 -23692
rect 16123 -23726 16157 -23692
rect 16381 -23726 16415 -23692
rect 9242 -24037 9276 -24003
rect 9500 -24037 9534 -24003
rect 9758 -24037 9792 -24003
rect 10016 -24037 10050 -24003
rect 10274 -24037 10308 -24003
rect 10532 -24037 10566 -24003
rect 10790 -24037 10824 -24003
rect 11048 -24037 11082 -24003
rect 11912 -24037 11946 -24003
rect 12170 -24037 12204 -24003
rect 12428 -24037 12462 -24003
rect 12686 -24037 12720 -24003
rect 12944 -24037 12978 -24003
rect 13202 -24037 13236 -24003
rect 13460 -24037 13494 -24003
rect 13718 -24037 13752 -24003
rect 14575 -24036 14609 -24002
rect 14833 -24036 14867 -24002
rect 15091 -24036 15125 -24002
rect 15349 -24036 15383 -24002
rect 15607 -24036 15641 -24002
rect 15865 -24036 15899 -24002
rect 16123 -24036 16157 -24002
rect 16381 -24036 16415 -24002
rect 9122 -24379 9156 -24345
rect 9662 -24379 9696 -24345
rect 10142 -24379 10176 -24345
rect 10645 -24377 10679 -24343
rect 11155 -24367 11189 -24333
rect 11792 -24379 11826 -24345
rect 12332 -24379 12366 -24345
rect 12812 -24379 12846 -24345
rect 13315 -24377 13349 -24343
rect 13825 -24367 13859 -24333
rect 14455 -24378 14489 -24344
rect 9122 -24689 9156 -24655
rect 9662 -24689 9696 -24655
rect 10142 -24689 10176 -24655
rect 10645 -24687 10679 -24653
rect 14995 -24378 15029 -24344
rect 15475 -24378 15509 -24344
rect 15978 -24376 16012 -24342
rect 16488 -24366 16522 -24332
rect 11155 -24677 11189 -24643
rect 11792 -24689 11826 -24655
rect 12332 -24689 12366 -24655
rect 12812 -24689 12846 -24655
rect 13315 -24687 13349 -24653
rect 13825 -24677 13859 -24643
rect 14455 -24688 14489 -24654
rect 14995 -24688 15029 -24654
rect 15475 -24688 15509 -24654
rect 15978 -24686 16012 -24652
rect 16488 -24676 16522 -24642
rect 18052 -7584 19420 -7550
rect 19913 -7584 21278 -7550
rect 18052 -9094 19420 -9060
rect 19913 -9094 21278 -9060
rect 18052 -10604 19420 -10570
rect 19913 -10604 21278 -10570
rect 18052 -12114 19420 -12080
rect 19913 -12114 21278 -12080
rect 18052 -13624 19420 -13590
rect 19913 -13624 21278 -13590
rect 18052 -15134 19420 -15100
rect 19913 -15134 21278 -15100
rect 18052 -16644 19420 -16610
rect 19913 -16644 21278 -16610
rect 18052 -18154 19420 -18120
rect 19913 -18154 21278 -18120
rect 18052 -19664 19420 -19630
rect 19913 -19664 21278 -19630
rect 18052 -21174 19420 -21140
rect 19913 -21174 21278 -21140
rect 18052 -22684 19420 -22650
rect 19913 -22684 21278 -22650
rect 18052 -24194 19420 -24160
rect 19913 -24194 21278 -24160
rect 18052 -25704 19420 -25670
rect 19913 -25704 21278 -25670
<< xpolycontact >>
rect -16256 49248 -16186 49680
rect -16256 44090 -16186 44522
rect -15938 49248 -15868 49680
rect -15938 44090 -15868 44522
rect -15620 49248 -15550 49680
rect -15620 44090 -15550 44522
rect -15302 49248 -15232 49680
rect -15302 44090 -15232 44522
rect -16204 41970 -16134 42402
rect -16204 36812 -16134 37244
rect -15848 41952 -15778 42384
rect -15848 36794 -15778 37226
rect -15530 41952 -15460 42384
rect -15530 36794 -15460 37226
rect -15132 41934 -15062 42366
rect -15132 36776 -15062 37208
rect -16212 35470 -16142 35902
rect -16212 30312 -16142 30744
rect -15874 35490 -15804 35922
rect -15874 30332 -15804 30764
rect -15556 35490 -15486 35922
rect -15556 30332 -15486 30764
rect -15186 35488 -15116 35920
rect -15186 30330 -15116 30762
rect -16190 28718 -16120 29150
rect -16190 23560 -16120 23992
rect -15872 28718 -15802 29150
rect -15872 23560 -15802 23992
rect -15554 28718 -15484 29150
rect -15554 23560 -15484 23992
rect -15236 28718 -15166 29150
rect -15236 23560 -15166 23992
rect 124 10732 556 10802
rect 4406 10732 4838 10802
rect 5354 10732 5786 10802
rect 9636 10732 10068 10802
rect 10584 10732 11016 10802
rect 14866 10732 15298 10802
rect 15814 10732 16246 10802
rect 20096 10732 20528 10802
rect 124 10412 556 10482
rect 4406 10412 4838 10482
rect 5354 10412 5786 10482
rect 9636 10412 10068 10482
rect 10584 10412 11016 10482
rect 14866 10412 15298 10482
rect 15814 10412 16246 10482
rect 20096 10412 20528 10482
rect 124 10092 556 10162
rect 4406 10092 4838 10162
rect 5368 10070 5800 10140
rect 9650 10070 10082 10140
rect 10564 10072 10996 10142
rect 14846 10072 15278 10142
rect 15814 10092 16246 10162
rect 20096 10092 20528 10162
rect 124 9772 556 9842
rect 4406 9772 4838 9842
rect 5368 9752 5800 9822
rect 9650 9752 10082 9822
rect 10564 9754 10996 9824
rect 14846 9754 15278 9824
rect 15814 9772 16246 9842
rect 20096 9772 20528 9842
rect 124 9452 556 9522
rect 4406 9452 4838 9522
rect 5368 9434 5800 9504
rect 9650 9434 10082 9504
rect 10564 9436 10996 9506
rect 14846 9436 15278 9506
rect 15814 9452 16246 9522
rect 20096 9452 20528 9522
rect 124 9132 556 9202
rect 4406 9132 4838 9202
rect 5368 9116 5800 9186
rect 9650 9116 10082 9186
rect 10564 9118 10996 9188
rect 14846 9118 15278 9188
rect 15814 9132 16246 9202
rect 20096 9132 20528 9202
rect 124 8812 556 8882
rect 4406 8812 4838 8882
rect 5368 8798 5800 8868
rect 9650 8798 10082 8868
rect 10564 8800 10996 8870
rect 14846 8800 15278 8870
rect 15814 8812 16246 8882
rect 20096 8812 20528 8882
rect 124 8492 556 8562
rect 4406 8492 4838 8562
rect 5368 8480 5800 8550
rect 9650 8480 10082 8550
rect 10564 8482 10996 8552
rect 14846 8482 15278 8552
rect 15814 8492 16246 8562
rect 20096 8492 20528 8562
rect 124 8172 556 8242
rect 4406 8172 4838 8242
rect 5368 8162 5800 8232
rect 9650 8162 10082 8232
rect 10564 8164 10996 8234
rect 14846 8164 15278 8234
rect 15814 8172 16246 8242
rect 20096 8172 20528 8242
rect 124 7852 556 7922
rect 4406 7852 4838 7922
rect 5368 7844 5800 7914
rect 9650 7844 10082 7914
rect 10564 7846 10996 7916
rect 14846 7846 15278 7916
rect 15814 7852 16246 7922
rect 20096 7852 20528 7922
rect 124 7532 556 7602
rect 4406 7532 4838 7602
rect 5368 7526 5800 7596
rect 9650 7526 10082 7596
rect 10564 7528 10996 7598
rect 14846 7528 15278 7598
rect 15814 7532 16246 7602
rect 20096 7532 20528 7602
rect 124 7212 556 7282
rect 4406 7212 4838 7282
rect 5388 7180 5820 7250
rect 9670 7180 10102 7250
rect 10584 7210 11016 7280
rect 14866 7210 15298 7280
rect 15814 7212 16246 7282
rect 20096 7212 20528 7282
rect 124 6892 556 6962
rect 4406 6892 4838 6962
rect 5388 6860 5820 6930
rect 9670 6860 10102 6930
rect 10584 6892 11016 6962
rect 14866 6892 15298 6962
rect 15814 6892 16246 6962
rect 20096 6892 20528 6962
<< xpolyres >>
rect -16256 44522 -16186 49248
rect -15938 44522 -15868 49248
rect -15620 44522 -15550 49248
rect -15302 44522 -15232 49248
rect -16204 37244 -16134 41970
rect -15848 37226 -15778 41952
rect -15530 37226 -15460 41952
rect -15132 37208 -15062 41934
rect -16212 30744 -16142 35470
rect -15874 30764 -15804 35490
rect -15556 30764 -15486 35490
rect -15186 30762 -15116 35488
rect -16190 23992 -16120 28718
rect -15872 23992 -15802 28718
rect -15554 23992 -15484 28718
rect -15236 23992 -15166 28718
rect 556 10732 4406 10802
rect 5786 10732 9636 10802
rect 11016 10732 14866 10802
rect 16246 10732 20096 10802
rect 556 10412 4406 10482
rect 5786 10412 9636 10482
rect 11016 10412 14866 10482
rect 16246 10412 20096 10482
rect 556 10092 4406 10162
rect 5800 10070 9650 10140
rect 10996 10072 14846 10142
rect 16246 10092 20096 10162
rect 556 9772 4406 9842
rect 5800 9752 9650 9822
rect 10996 9754 14846 9824
rect 16246 9772 20096 9842
rect 556 9452 4406 9522
rect 5800 9434 9650 9504
rect 10996 9436 14846 9506
rect 16246 9452 20096 9522
rect 556 9132 4406 9202
rect 5800 9116 9650 9186
rect 10996 9118 14846 9188
rect 16246 9132 20096 9202
rect 556 8812 4406 8882
rect 5800 8798 9650 8868
rect 10996 8800 14846 8870
rect 16246 8812 20096 8882
rect 556 8492 4406 8562
rect 5800 8480 9650 8550
rect 10996 8482 14846 8552
rect 16246 8492 20096 8562
rect 556 8172 4406 8242
rect 5800 8162 9650 8232
rect 10996 8164 14846 8234
rect 16246 8172 20096 8242
rect 556 7852 4406 7922
rect 5800 7844 9650 7914
rect 10996 7846 14846 7916
rect 16246 7852 20096 7922
rect 556 7532 4406 7602
rect 5800 7526 9650 7596
rect 10996 7528 14846 7598
rect 16246 7532 20096 7602
rect 556 7212 4406 7282
rect 5820 7180 9670 7250
rect 11016 7210 14866 7280
rect 16246 7212 20096 7282
rect 556 6892 4406 6962
rect 5820 6860 9670 6930
rect 11016 6892 14866 6962
rect 16246 6892 20096 6962
<< locali >>
rect -19220 56190 -17382 56450
rect -19220 55462 -18978 56190
rect -17592 55462 -17382 56190
rect -19220 55220 -17382 55462
rect -15220 56190 -13382 56450
rect -15220 55462 -14978 56190
rect -13592 55462 -13382 56190
rect -15220 55220 -13382 55462
rect -11220 56190 -9382 56450
rect -11220 55462 -10978 56190
rect -9592 55462 -9382 56190
rect -11220 55220 -9382 55462
rect -7220 56190 -5382 56450
rect -7220 55462 -6978 56190
rect -5592 55462 -5382 56190
rect -7220 55220 -5382 55462
rect -3220 56190 -1382 56450
rect -3220 55462 -2978 56190
rect -1592 55462 -1382 56190
rect -3220 55220 -1382 55462
rect 780 56190 2618 56450
rect 780 55462 1022 56190
rect 2408 55462 2618 56190
rect 780 55220 2618 55462
rect 4780 56190 6618 56450
rect 4780 55462 5022 56190
rect 6408 55462 6618 56190
rect 4780 55220 6618 55462
rect 8780 56190 10618 56450
rect 8780 55462 9022 56190
rect 10408 55462 10618 56190
rect 8780 55220 10618 55462
rect 12780 56190 14618 56450
rect 12780 55462 13022 56190
rect 14408 55462 14618 56190
rect 12780 55220 14618 55462
rect 16780 56190 18618 56450
rect 16780 55462 17022 56190
rect 18408 55462 18618 56190
rect 16780 55220 18618 55462
rect 20780 56190 22618 56450
rect 20780 55462 21022 56190
rect 22408 55462 22618 56190
rect 20780 55220 22618 55462
rect 24780 56190 26618 56450
rect 24780 55462 25022 56190
rect 26408 55462 26618 56190
rect 24780 55220 26618 55462
rect 28780 56190 30618 56450
rect 28780 55462 29022 56190
rect 30408 55462 30618 56190
rect 28780 55220 30618 55462
rect 32780 56190 34618 56450
rect 32780 55462 33022 56190
rect 34408 55462 34618 56190
rect 32780 55220 34618 55462
rect 36780 56190 38618 56450
rect 36780 55462 37022 56190
rect 38408 55462 38618 56190
rect 36780 55220 38618 55462
rect -20956 54026 -19118 54286
rect -20956 53298 -20714 54026
rect -19328 53298 -19118 54026
rect -20956 53056 -19118 53298
rect 36822 52988 38660 53256
rect 36822 52260 37064 52988
rect 38450 52260 38660 52988
rect 36822 52018 38660 52260
rect -20956 50026 -19118 50286
rect -20956 49298 -20714 50026
rect -19328 49298 -19118 50026
rect -20956 49056 -19118 49298
rect 36822 48988 38660 49256
rect 36822 48260 37064 48988
rect 38450 48260 38660 48988
rect 36822 48018 38660 48260
rect -20956 46026 -19118 46286
rect -20956 45298 -20714 46026
rect -19328 45298 -19118 46026
rect -20956 45056 -19118 45298
rect 36822 44988 38660 45256
rect 36822 44260 37064 44988
rect 38450 44260 38660 44988
rect 36822 44018 38660 44260
rect -20956 42026 -19118 42286
rect -20956 41298 -20714 42026
rect -19328 41298 -19118 42026
rect -20956 41056 -19118 41298
rect 36822 40988 38660 41256
rect 36822 40260 37064 40988
rect 38450 40260 38660 40988
rect 36822 40018 38660 40260
rect -20956 38026 -19118 38286
rect -20956 37298 -20714 38026
rect -19328 37298 -19118 38026
rect -20956 37056 -19118 37298
rect 36822 36988 38660 37256
rect 36822 36260 37064 36988
rect 38450 36260 38660 36988
rect 36822 36018 38660 36260
rect -20956 34026 -19118 34286
rect -20956 33298 -20714 34026
rect -19328 33298 -19118 34026
rect -20956 33056 -19118 33298
rect 36822 32988 38660 33256
rect 36822 32260 37064 32988
rect 38450 32260 38660 32988
rect 36822 32018 38660 32260
rect -20956 30026 -19118 30286
rect -20956 29298 -20714 30026
rect -19328 29298 -19118 30026
rect -20956 29056 -19118 29298
rect 36822 28988 38660 29256
rect 36822 28260 37064 28988
rect 38450 28260 38660 28988
rect 36822 28018 38660 28260
rect -20956 26026 -19118 26286
rect -20956 25298 -20714 26026
rect -19328 25298 -19118 26026
rect -20956 25056 -19118 25298
rect 36822 24988 38660 25256
rect 36822 24260 37064 24988
rect 38450 24260 38660 24988
rect 36822 24018 38660 24260
rect -20956 22026 -19118 22286
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -94226 20649 -93238 20840
rect -94226 20615 -94156 20649
rect -93372 20615 -93238 20649
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -94226 19121 -93238 20615
rect -92574 20649 -91586 20910
rect -92574 20615 -92498 20649
rect -91714 20615 -91586 20649
rect -94226 19087 -94156 19121
rect -93372 19087 -93238 19121
rect -94226 19013 -93238 19087
rect -94226 18979 -94156 19013
rect -93372 18979 -93238 19013
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -94226 17485 -93238 18979
rect -92574 19121 -91586 20615
rect -90968 20649 -89980 20840
rect -90968 20615 -90840 20649
rect -90056 20615 -89980 20649
rect -92574 19087 -92498 19121
rect -91714 19087 -91586 19121
rect -92574 19013 -91586 19087
rect -92574 18979 -92498 19013
rect -91714 18979 -91586 19013
rect -94226 17451 -94156 17485
rect -93372 17451 -93238 17485
rect -94226 17267 -93238 17451
rect -94226 17233 -94154 17267
rect -93370 17233 -93238 17267
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -94226 15739 -93238 17233
rect -92574 17485 -91586 18979
rect -90968 19121 -89980 20615
rect -89268 20649 -88280 20910
rect -89268 20615 -89182 20649
rect -88398 20615 -88280 20649
rect -90968 19087 -90840 19121
rect -90056 19087 -89980 19121
rect -90968 19013 -89980 19087
rect -90968 18979 -90840 19013
rect -90056 18979 -89980 19013
rect -92574 17451 -92498 17485
rect -91714 17451 -91586 17485
rect -92574 17267 -91586 17451
rect -92574 17233 -92496 17267
rect -91712 17233 -91586 17267
rect -94226 15705 -94154 15739
rect -93370 15705 -93238 15739
rect -94226 15631 -93238 15705
rect -94226 15597 -94154 15631
rect -93370 15597 -93238 15631
rect -96266 13740 -95320 15274
rect -94226 14103 -93238 15597
rect -92574 15739 -91586 17233
rect -90968 17485 -89980 18979
rect -89268 19121 -88280 20615
rect -87640 20649 -86652 20886
rect -87640 20615 -87524 20649
rect -86740 20615 -86652 20649
rect -89268 19087 -89182 19121
rect -88398 19087 -88280 19121
rect -89268 19013 -88280 19087
rect -89268 18979 -89182 19013
rect -88398 18979 -88280 19013
rect -90968 17451 -90840 17485
rect -90056 17451 -89980 17485
rect -90968 17267 -89980 17451
rect -90968 17233 -90838 17267
rect -90054 17233 -89980 17267
rect -92574 15705 -92496 15739
rect -91712 15705 -91586 15739
rect -92574 15631 -91586 15705
rect -92574 15597 -92496 15631
rect -91712 15597 -91586 15631
rect -94226 14069 -94154 14103
rect -93370 14069 -93238 14103
rect -94226 13995 -93238 14069
rect -94226 13961 -94154 13995
rect -93370 13961 -93238 13995
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -94226 12467 -93238 13961
rect -92574 14103 -91586 15597
rect -90968 15739 -89980 17233
rect -89268 17485 -88280 18979
rect -87640 19121 -86652 20615
rect -85964 20649 -84976 20910
rect -85964 20615 -85866 20649
rect -85082 20615 -84976 20649
rect -87640 19087 -87524 19121
rect -86740 19087 -86652 19121
rect -87640 19013 -86652 19087
rect -87640 18979 -87524 19013
rect -86740 18979 -86652 19013
rect -89268 17451 -89182 17485
rect -88398 17451 -88280 17485
rect -89268 17267 -88280 17451
rect -89268 17233 -89180 17267
rect -88396 17233 -88280 17267
rect -90968 15705 -90838 15739
rect -90054 15705 -89980 15739
rect -90968 15631 -89980 15705
rect -90968 15597 -90838 15631
rect -90054 15597 -89980 15631
rect -92574 14069 -92496 14103
rect -91712 14069 -91586 14103
rect -92574 13995 -91586 14069
rect -92574 13961 -92496 13995
rect -91712 13961 -91586 13995
rect -94226 12433 -94154 12467
rect -93370 12433 -93238 12467
rect -94226 12359 -93238 12433
rect -94226 12325 -94154 12359
rect -93370 12325 -93238 12359
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -94226 10831 -93238 12325
rect -92574 12467 -91586 13961
rect -90968 14103 -89980 15597
rect -89268 15739 -88280 17233
rect -87640 17485 -86652 18979
rect -85964 19121 -84976 20615
rect -84312 20649 -83324 20864
rect -84312 20615 -84208 20649
rect -83424 20615 -83324 20649
rect -85964 19087 -85866 19121
rect -85082 19087 -84976 19121
rect -85964 19013 -84976 19087
rect -85964 18979 -85866 19013
rect -85082 18979 -84976 19013
rect -87640 17451 -87524 17485
rect -86740 17451 -86652 17485
rect -87640 17267 -86652 17451
rect -87640 17233 -87522 17267
rect -86738 17233 -86652 17267
rect -89268 15705 -89180 15739
rect -88396 15705 -88280 15739
rect -89268 15631 -88280 15705
rect -89268 15597 -89180 15631
rect -88396 15597 -88280 15631
rect -90968 14069 -90838 14103
rect -90054 14069 -89980 14103
rect -90968 13995 -89980 14069
rect -90968 13961 -90838 13995
rect -90054 13961 -89980 13995
rect -92574 12433 -92496 12467
rect -91712 12433 -91586 12467
rect -92574 12359 -91586 12433
rect -92574 12325 -92496 12359
rect -91712 12325 -91586 12359
rect -94226 10797 -94154 10831
rect -93370 10797 -93238 10831
rect -94226 10721 -93238 10797
rect -94226 10687 -94154 10721
rect -93370 10687 -93238 10721
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -94226 9193 -93238 10687
rect -92574 10831 -91586 12325
rect -90968 12467 -89980 13961
rect -89268 14103 -88280 15597
rect -87640 15739 -86652 17233
rect -85964 17485 -84976 18979
rect -84312 19121 -83324 20615
rect -82682 20649 -81694 20886
rect -82682 20615 -82550 20649
rect -81766 20615 -81694 20649
rect -84312 19087 -84208 19121
rect -83424 19087 -83324 19121
rect -84312 19013 -83324 19087
rect -84312 18979 -84208 19013
rect -83424 18979 -83324 19013
rect -85964 17451 -85866 17485
rect -85082 17451 -84976 17485
rect -85964 17267 -84976 17451
rect -85964 17233 -85864 17267
rect -85080 17233 -84976 17267
rect -87640 15705 -87522 15739
rect -86738 15705 -86652 15739
rect -87640 15631 -86652 15705
rect -87640 15597 -87522 15631
rect -86738 15597 -86652 15631
rect -89268 14069 -89180 14103
rect -88396 14069 -88280 14103
rect -89268 13995 -88280 14069
rect -89268 13961 -89180 13995
rect -88396 13961 -88280 13995
rect -90968 12433 -90838 12467
rect -90054 12433 -89980 12467
rect -90968 12359 -89980 12433
rect -90968 12325 -90838 12359
rect -90054 12325 -89980 12359
rect -92574 10797 -92496 10831
rect -91712 10797 -91586 10831
rect -92574 10721 -91586 10797
rect -92574 10687 -92496 10721
rect -91712 10687 -91586 10721
rect -94226 9159 -94154 9193
rect -93370 9159 -93238 9193
rect -94226 9085 -93238 9159
rect -94226 9051 -94154 9085
rect -93370 9051 -93238 9085
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -94226 7557 -93238 9051
rect -92574 9193 -91586 10687
rect -90968 10831 -89980 12325
rect -89268 12467 -88280 13961
rect -87640 14103 -86652 15597
rect -85964 15739 -84976 17233
rect -84312 17485 -83324 18979
rect -82682 19121 -81694 20615
rect -81030 20649 -80042 20864
rect -81030 20615 -80892 20649
rect -80108 20615 -80042 20649
rect -82682 19087 -82550 19121
rect -81766 19087 -81694 19121
rect -82682 19013 -81694 19087
rect -82682 18979 -82550 19013
rect -81766 18979 -81694 19013
rect -84312 17451 -84208 17485
rect -83424 17451 -83324 17485
rect -84312 17267 -83324 17451
rect -84312 17233 -84206 17267
rect -83422 17233 -83324 17267
rect -85964 15705 -85864 15739
rect -85080 15705 -84976 15739
rect -85964 15631 -84976 15705
rect -85964 15597 -85864 15631
rect -85080 15597 -84976 15631
rect -87640 14069 -87522 14103
rect -86738 14069 -86652 14103
rect -87640 13995 -86652 14069
rect -87640 13961 -87522 13995
rect -86738 13961 -86652 13995
rect -89268 12433 -89180 12467
rect -88396 12433 -88280 12467
rect -89268 12359 -88280 12433
rect -89268 12325 -89180 12359
rect -88396 12325 -88280 12359
rect -90968 10797 -90838 10831
rect -90054 10797 -89980 10831
rect -90968 10721 -89980 10797
rect -90968 10687 -90838 10721
rect -90054 10687 -89980 10721
rect -92574 9159 -92496 9193
rect -91712 9159 -91586 9193
rect -92574 9085 -91586 9159
rect -92574 9051 -92496 9085
rect -91712 9051 -91586 9085
rect -94226 7523 -94154 7557
rect -93370 7523 -93238 7557
rect -94226 7449 -93238 7523
rect -94226 7415 -94154 7449
rect -93370 7415 -93238 7449
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -94226 5921 -93238 7415
rect -92574 7557 -91586 9051
rect -90968 9193 -89980 10687
rect -89268 10831 -88280 12325
rect -87640 12467 -86652 13961
rect -85964 14103 -84976 15597
rect -84312 15739 -83324 17233
rect -82682 17485 -81694 18979
rect -81030 19121 -80042 20615
rect -79330 20649 -78342 20886
rect -79330 20615 -79234 20649
rect -78450 20615 -78342 20649
rect -81030 19087 -80892 19121
rect -80108 19087 -80042 19121
rect -81030 19013 -80042 19087
rect -81030 18979 -80892 19013
rect -80108 18979 -80042 19013
rect -82682 17451 -82550 17485
rect -81766 17451 -81694 17485
rect -82682 17267 -81694 17451
rect -82682 17233 -82548 17267
rect -81764 17233 -81694 17267
rect -84312 15705 -84206 15739
rect -83422 15705 -83324 15739
rect -84312 15631 -83324 15705
rect -84312 15597 -84206 15631
rect -83422 15597 -83324 15631
rect -85964 14069 -85864 14103
rect -85080 14069 -84976 14103
rect -85964 13995 -84976 14069
rect -85964 13961 -85864 13995
rect -85080 13961 -84976 13995
rect -87640 12433 -87522 12467
rect -86738 12433 -86652 12467
rect -87640 12359 -86652 12433
rect -87640 12325 -87522 12359
rect -86738 12325 -86652 12359
rect -89268 10797 -89180 10831
rect -88396 10797 -88280 10831
rect -89268 10721 -88280 10797
rect -89268 10687 -89180 10721
rect -88396 10687 -88280 10721
rect -90968 9159 -90838 9193
rect -90054 9159 -89980 9193
rect -90968 9085 -89980 9159
rect -90968 9051 -90838 9085
rect -90054 9051 -89980 9085
rect -92574 7523 -92496 7557
rect -91712 7523 -91586 7557
rect -92574 7449 -91586 7523
rect -92574 7415 -92496 7449
rect -91712 7415 -91586 7449
rect -94226 5887 -94154 5921
rect -93370 5887 -93238 5921
rect -94226 5813 -93238 5887
rect -94226 5779 -94154 5813
rect -93370 5779 -93238 5813
rect -96266 4182 -95320 5274
rect -94226 4285 -93238 5779
rect -92574 5921 -91586 7415
rect -90968 7557 -89980 9051
rect -89268 9193 -88280 10687
rect -87640 10831 -86652 12325
rect -85964 12467 -84976 13961
rect -84312 14103 -83324 15597
rect -82682 15739 -81694 17233
rect -81030 17485 -80042 18979
rect -79330 19121 -78342 20615
rect -77772 20649 -76784 20886
rect -76024 20649 -75036 20910
rect -77772 20615 -77576 20649
rect -76792 20615 -76776 20649
rect -76024 20615 -75918 20649
rect -75134 20615 -75036 20649
rect -79330 19087 -79234 19121
rect -78450 19087 -78342 19121
rect -79330 19013 -78342 19087
rect -79330 18979 -79234 19013
rect -78450 18979 -78342 19013
rect -81030 17451 -80892 17485
rect -80108 17451 -80042 17485
rect -81030 17267 -80042 17451
rect -81030 17233 -80890 17267
rect -80106 17233 -80042 17267
rect -82682 15705 -82548 15739
rect -81764 15705 -81694 15739
rect -82682 15631 -81694 15705
rect -82682 15597 -82548 15631
rect -81764 15597 -81694 15631
rect -84312 14069 -84206 14103
rect -83422 14069 -83324 14103
rect -84312 13995 -83324 14069
rect -84312 13961 -84206 13995
rect -83422 13961 -83324 13995
rect -85964 12433 -85864 12467
rect -85080 12433 -84976 12467
rect -85964 12359 -84976 12433
rect -85964 12325 -85864 12359
rect -85080 12325 -84976 12359
rect -87640 10797 -87522 10831
rect -86738 10797 -86652 10831
rect -87640 10721 -86652 10797
rect -87640 10687 -87522 10721
rect -86738 10687 -86652 10721
rect -89268 9159 -89180 9193
rect -88396 9159 -88280 9193
rect -89268 9085 -88280 9159
rect -89268 9051 -89180 9085
rect -88396 9051 -88280 9085
rect -90968 7523 -90838 7557
rect -90054 7523 -89980 7557
rect -90968 7449 -89980 7523
rect -90968 7415 -90838 7449
rect -90054 7415 -89980 7449
rect -92574 5887 -92496 5921
rect -91712 5887 -91586 5921
rect -92574 5813 -91586 5887
rect -92574 5779 -92496 5813
rect -91712 5779 -91586 5813
rect -94226 4251 -94154 4285
rect -93370 4251 -93238 4285
rect -94226 4220 -93238 4251
rect -92574 4285 -91586 5779
rect -90968 5921 -89980 7415
rect -89268 7557 -88280 9051
rect -87640 9193 -86652 10687
rect -85964 10831 -84976 12325
rect -84312 12467 -83324 13961
rect -82682 14103 -81694 15597
rect -81030 15739 -80042 17233
rect -79330 17485 -78342 18979
rect -77772 19121 -76784 20615
rect -76024 19121 -75036 20615
rect -74372 20649 -73384 20910
rect -74372 20615 -74260 20649
rect -73476 20615 -73384 20649
rect -77772 19087 -77576 19121
rect -76792 19087 -76776 19121
rect -76024 19087 -75918 19121
rect -75134 19087 -75036 19121
rect -77772 19013 -76784 19087
rect -76024 19013 -75036 19087
rect -77772 18979 -77576 19013
rect -76792 18979 -76776 19013
rect -76024 18979 -75918 19013
rect -75134 18979 -75036 19013
rect -79330 17451 -79234 17485
rect -78450 17451 -78342 17485
rect -79330 17267 -78342 17451
rect -79330 17233 -79232 17267
rect -78448 17233 -78342 17267
rect -81030 15705 -80890 15739
rect -80106 15705 -80042 15739
rect -81030 15631 -80042 15705
rect -81030 15597 -80890 15631
rect -80106 15597 -80042 15631
rect -82682 14069 -82548 14103
rect -81764 14069 -81694 14103
rect -82682 13995 -81694 14069
rect -82682 13961 -82548 13995
rect -81764 13961 -81694 13995
rect -84312 12433 -84206 12467
rect -83422 12433 -83324 12467
rect -84312 12359 -83324 12433
rect -84312 12325 -84206 12359
rect -83422 12325 -83324 12359
rect -85964 10797 -85864 10831
rect -85080 10797 -84976 10831
rect -85964 10721 -84976 10797
rect -85964 10687 -85864 10721
rect -85080 10687 -84976 10721
rect -87640 9159 -87522 9193
rect -86738 9159 -86652 9193
rect -87640 9085 -86652 9159
rect -87640 9051 -87522 9085
rect -86738 9051 -86652 9085
rect -89268 7523 -89180 7557
rect -88396 7523 -88280 7557
rect -89268 7449 -88280 7523
rect -89268 7415 -89180 7449
rect -88396 7415 -88280 7449
rect -90968 5887 -90838 5921
rect -90054 5887 -89980 5921
rect -90968 5813 -89980 5887
rect -90968 5779 -90838 5813
rect -90054 5779 -89980 5813
rect -92574 4251 -92496 4285
rect -91712 4251 -91586 4285
rect -92574 4220 -91586 4251
rect -90968 4285 -89980 5779
rect -89268 5921 -88280 7415
rect -87640 7557 -86652 9051
rect -85964 9193 -84976 10687
rect -84312 10831 -83324 12325
rect -82682 12467 -81694 13961
rect -81030 14103 -80042 15597
rect -79330 15739 -78342 17233
rect -77772 17485 -76784 18979
rect -76024 17485 -75036 18979
rect -74372 19121 -73384 20615
rect -72742 20649 -71754 20910
rect -72742 20615 -72602 20649
rect -71818 20615 -71754 20649
rect -74372 19087 -74260 19121
rect -73476 19087 -73384 19121
rect -74372 19013 -73384 19087
rect -74372 18979 -74260 19013
rect -73476 18979 -73384 19013
rect -77772 17451 -77576 17485
rect -76792 17451 -76776 17485
rect -76024 17451 -75918 17485
rect -75134 17451 -75036 17485
rect -77772 17267 -76784 17451
rect -76024 17267 -75036 17451
rect -77772 17233 -77574 17267
rect -76790 17233 -76774 17267
rect -76024 17233 -75916 17267
rect -75132 17233 -75036 17267
rect -79330 15705 -79232 15739
rect -78448 15705 -78342 15739
rect -79330 15631 -78342 15705
rect -79330 15597 -79232 15631
rect -78448 15597 -78342 15631
rect -81030 14069 -80890 14103
rect -80106 14069 -80042 14103
rect -81030 13995 -80042 14069
rect -81030 13961 -80890 13995
rect -80106 13961 -80042 13995
rect -82682 12433 -82548 12467
rect -81764 12433 -81694 12467
rect -82682 12359 -81694 12433
rect -82682 12325 -82548 12359
rect -81764 12325 -81694 12359
rect -84312 10797 -84206 10831
rect -83422 10797 -83324 10831
rect -84312 10721 -83324 10797
rect -84312 10687 -84206 10721
rect -83422 10687 -83324 10721
rect -85964 9159 -85864 9193
rect -85080 9159 -84976 9193
rect -85964 9085 -84976 9159
rect -85964 9051 -85864 9085
rect -85080 9051 -84976 9085
rect -87640 7523 -87522 7557
rect -86738 7523 -86652 7557
rect -87640 7449 -86652 7523
rect -87640 7415 -87522 7449
rect -86738 7415 -86652 7449
rect -89268 5887 -89180 5921
rect -88396 5887 -88280 5921
rect -89268 5813 -88280 5887
rect -89268 5779 -89180 5813
rect -88396 5779 -88280 5813
rect -90968 4251 -90838 4285
rect -90054 4251 -89980 4285
rect -90968 4220 -89980 4251
rect -89268 4285 -88280 5779
rect -87640 5921 -86652 7415
rect -85964 7557 -84976 9051
rect -84312 9193 -83324 10687
rect -82682 10831 -81694 12325
rect -81030 12467 -80042 13961
rect -79330 14103 -78342 15597
rect -77772 15739 -76784 17233
rect -76024 15739 -75036 17233
rect -74372 17485 -73384 18979
rect -72742 19121 -71754 20615
rect -71064 20649 -70076 20910
rect -71064 20615 -70944 20649
rect -70160 20615 -70076 20649
rect -72742 19087 -72602 19121
rect -71818 19087 -71754 19121
rect -72742 19013 -71754 19087
rect -72742 18979 -72602 19013
rect -71818 18979 -71754 19013
rect -74372 17451 -74260 17485
rect -73476 17451 -73384 17485
rect -74372 17267 -73384 17451
rect -74372 17233 -74258 17267
rect -73474 17233 -73384 17267
rect -77772 15705 -77574 15739
rect -76790 15705 -76774 15739
rect -76024 15705 -75916 15739
rect -75132 15705 -75036 15739
rect -77772 15631 -76784 15705
rect -76024 15631 -75036 15705
rect -77772 15597 -77574 15631
rect -76790 15597 -76774 15631
rect -76024 15597 -75916 15631
rect -75132 15597 -75036 15631
rect -79330 14069 -79232 14103
rect -78448 14069 -78342 14103
rect -79330 13995 -78342 14069
rect -79330 13961 -79232 13995
rect -78448 13961 -78342 13995
rect -81030 12433 -80890 12467
rect -80106 12433 -80042 12467
rect -81030 12359 -80042 12433
rect -81030 12325 -80890 12359
rect -80106 12325 -80042 12359
rect -82682 10797 -82548 10831
rect -81764 10797 -81694 10831
rect -82682 10721 -81694 10797
rect -82682 10687 -82548 10721
rect -81764 10687 -81694 10721
rect -84312 9159 -84206 9193
rect -83422 9159 -83324 9193
rect -84312 9085 -83324 9159
rect -84312 9051 -84206 9085
rect -83422 9051 -83324 9085
rect -85964 7523 -85864 7557
rect -85080 7523 -84976 7557
rect -85964 7449 -84976 7523
rect -85964 7415 -85864 7449
rect -85080 7415 -84976 7449
rect -87640 5887 -87522 5921
rect -86738 5887 -86652 5921
rect -87640 5813 -86652 5887
rect -87640 5779 -87522 5813
rect -86738 5779 -86652 5813
rect -89268 4251 -89180 4285
rect -88396 4251 -88280 4285
rect -89268 4220 -88280 4251
rect -87640 4285 -86652 5779
rect -85964 5921 -84976 7415
rect -84312 7557 -83324 9051
rect -82682 9193 -81694 10687
rect -81030 10831 -80042 12325
rect -79330 12467 -78342 13961
rect -77772 14103 -76784 15597
rect -76024 14103 -75036 15597
rect -74372 15739 -73384 17233
rect -72742 17485 -71754 18979
rect -71064 19121 -70076 20615
rect -69366 20649 -68378 20886
rect -69366 20615 -69286 20649
rect -68502 20615 -68378 20649
rect -71064 19087 -70944 19121
rect -70160 19087 -70076 19121
rect -71064 19013 -70076 19087
rect -71064 18979 -70944 19013
rect -70160 18979 -70076 19013
rect -72742 17451 -72602 17485
rect -71818 17451 -71754 17485
rect -72742 17267 -71754 17451
rect -72742 17233 -72600 17267
rect -71816 17233 -71754 17267
rect -74372 15705 -74258 15739
rect -73474 15705 -73384 15739
rect -74372 15631 -73384 15705
rect -74372 15597 -74258 15631
rect -73474 15597 -73384 15631
rect -77772 14069 -77574 14103
rect -76790 14069 -76774 14103
rect -76024 14069 -75916 14103
rect -75132 14069 -75036 14103
rect -77772 13995 -76784 14069
rect -76024 13995 -75036 14069
rect -77772 13961 -77574 13995
rect -76790 13961 -76774 13995
rect -76024 13961 -75916 13995
rect -75132 13961 -75036 13995
rect -79330 12433 -79232 12467
rect -78448 12433 -78342 12467
rect -79330 12359 -78342 12433
rect -79330 12325 -79232 12359
rect -78448 12325 -78342 12359
rect -81030 10797 -80890 10831
rect -80106 10797 -80042 10831
rect -81030 10721 -80042 10797
rect -81030 10687 -80890 10721
rect -80106 10687 -80042 10721
rect -82682 9159 -82548 9193
rect -81764 9159 -81694 9193
rect -82682 9085 -81694 9159
rect -82682 9051 -82548 9085
rect -81764 9051 -81694 9085
rect -84312 7523 -84206 7557
rect -83422 7523 -83324 7557
rect -84312 7449 -83324 7523
rect -84312 7415 -84206 7449
rect -83422 7415 -83324 7449
rect -85964 5887 -85864 5921
rect -85080 5887 -84976 5921
rect -85964 5813 -84976 5887
rect -85964 5779 -85864 5813
rect -85080 5779 -84976 5813
rect -87640 4251 -87522 4285
rect -86738 4251 -86652 4285
rect -87640 4220 -86652 4251
rect -85964 4285 -84976 5779
rect -84312 5921 -83324 7415
rect -82682 7557 -81694 9051
rect -81030 9193 -80042 10687
rect -79330 10831 -78342 12325
rect -77772 12467 -76784 13961
rect -76024 12467 -75036 13961
rect -74372 14103 -73384 15597
rect -72742 15739 -71754 17233
rect -71064 17485 -70076 18979
rect -69366 19121 -68378 20615
rect -67736 20649 -66748 20934
rect -67736 20615 -67628 20649
rect -66844 20615 -66748 20649
rect -69366 19087 -69286 19121
rect -68502 19087 -68378 19121
rect -69366 19013 -68378 19087
rect -69366 18979 -69286 19013
rect -68502 18979 -68378 19013
rect -71064 17451 -70944 17485
rect -70160 17451 -70076 17485
rect -71064 17267 -70076 17451
rect -71064 17233 -70942 17267
rect -70158 17233 -70076 17267
rect -72742 15705 -72600 15739
rect -71816 15705 -71754 15739
rect -72742 15631 -71754 15705
rect -72742 15597 -72600 15631
rect -71816 15597 -71754 15631
rect -74372 14069 -74258 14103
rect -73474 14069 -73384 14103
rect -74372 13995 -73384 14069
rect -74372 13961 -74258 13995
rect -73474 13961 -73384 13995
rect -77772 12433 -77574 12467
rect -76790 12433 -76774 12467
rect -76024 12433 -75916 12467
rect -75132 12433 -75036 12467
rect -77772 12359 -76784 12433
rect -76024 12359 -75036 12433
rect -77772 12325 -77574 12359
rect -76790 12325 -76774 12359
rect -76024 12325 -75916 12359
rect -75132 12325 -75036 12359
rect -79330 10797 -79232 10831
rect -78448 10797 -78342 10831
rect -79330 10721 -78342 10797
rect -79330 10687 -79232 10721
rect -78448 10687 -78342 10721
rect -81030 9159 -80890 9193
rect -80106 9159 -80042 9193
rect -81030 9085 -80042 9159
rect -81030 9051 -80890 9085
rect -80106 9051 -80042 9085
rect -82682 7523 -82548 7557
rect -81764 7523 -81694 7557
rect -82682 7449 -81694 7523
rect -82682 7415 -82548 7449
rect -81764 7415 -81694 7449
rect -84312 5887 -84206 5921
rect -83422 5887 -83324 5921
rect -84312 5813 -83324 5887
rect -84312 5779 -84206 5813
rect -83422 5779 -83324 5813
rect -85964 4251 -85864 4285
rect -85080 4251 -84976 4285
rect -85964 4220 -84976 4251
rect -84312 4285 -83324 5779
rect -82682 5921 -81694 7415
rect -81030 7557 -80042 9051
rect -79330 9193 -78342 10687
rect -77772 10831 -76784 12325
rect -76024 10831 -75036 12325
rect -74372 12467 -73384 13961
rect -72742 14103 -71754 15597
rect -71064 15739 -70076 17233
rect -69366 17485 -68378 18979
rect -67736 19121 -66748 20615
rect -66060 20649 -65072 20910
rect -66060 20615 -65970 20649
rect -65186 20615 -65072 20649
rect -67736 19087 -67628 19121
rect -66844 19087 -66748 19121
rect -67736 19013 -66748 19087
rect -67736 18979 -67628 19013
rect -66844 18979 -66748 19013
rect -69366 17451 -69286 17485
rect -68502 17451 -68378 17485
rect -69366 17267 -68378 17451
rect -69366 17233 -69284 17267
rect -68500 17233 -68378 17267
rect -71064 15705 -70942 15739
rect -70158 15705 -70076 15739
rect -71064 15631 -70076 15705
rect -71064 15597 -70942 15631
rect -70158 15597 -70076 15631
rect -72742 14069 -72600 14103
rect -71816 14069 -71754 14103
rect -72742 13995 -71754 14069
rect -72742 13961 -72600 13995
rect -71816 13961 -71754 13995
rect -74372 12433 -74258 12467
rect -73474 12433 -73384 12467
rect -74372 12359 -73384 12433
rect -74372 12325 -74258 12359
rect -73474 12325 -73384 12359
rect -77772 10797 -77574 10831
rect -76790 10797 -76774 10831
rect -76024 10797 -75916 10831
rect -75132 10797 -75036 10831
rect -77772 10721 -76784 10797
rect -76024 10721 -75036 10797
rect -77772 10687 -77574 10721
rect -76790 10687 -76774 10721
rect -76024 10687 -75916 10721
rect -75132 10687 -75036 10721
rect -79330 9159 -79232 9193
rect -78448 9159 -78342 9193
rect -79330 9085 -78342 9159
rect -79330 9051 -79232 9085
rect -78448 9051 -78342 9085
rect -81030 7523 -80890 7557
rect -80106 7523 -80042 7557
rect -81030 7449 -80042 7523
rect -81030 7415 -80890 7449
rect -80106 7415 -80042 7449
rect -82682 5887 -82548 5921
rect -81764 5887 -81694 5921
rect -82682 5813 -81694 5887
rect -82682 5779 -82548 5813
rect -81764 5779 -81694 5813
rect -84312 4251 -84206 4285
rect -83422 4251 -83324 4285
rect -84312 4220 -83324 4251
rect -82682 4285 -81694 5779
rect -81030 5921 -80042 7415
rect -79330 7557 -78342 9051
rect -77772 9193 -76784 10687
rect -76024 9193 -75036 10687
rect -74372 10831 -73384 12325
rect -72742 12467 -71754 13961
rect -71064 14103 -70076 15597
rect -69366 15739 -68378 17233
rect -67736 17485 -66748 18979
rect -66060 19121 -65072 20615
rect -64408 20649 -63420 20934
rect -64408 20615 -64312 20649
rect -63528 20615 -63420 20649
rect -66060 19087 -65970 19121
rect -65186 19087 -65072 19121
rect -66060 19013 -65072 19087
rect -66060 18979 -65970 19013
rect -65186 18979 -65072 19013
rect -67736 17451 -67628 17485
rect -66844 17451 -66748 17485
rect -67736 17267 -66748 17451
rect -67736 17233 -67626 17267
rect -66842 17233 -66748 17267
rect -69366 15705 -69284 15739
rect -68500 15705 -68378 15739
rect -69366 15631 -68378 15705
rect -69366 15597 -69284 15631
rect -68500 15597 -68378 15631
rect -71064 14069 -70942 14103
rect -70158 14069 -70076 14103
rect -71064 13995 -70076 14069
rect -71064 13961 -70942 13995
rect -70158 13961 -70076 13995
rect -72742 12433 -72600 12467
rect -71816 12433 -71754 12467
rect -72742 12359 -71754 12433
rect -72742 12325 -72600 12359
rect -71816 12325 -71754 12359
rect -74372 10797 -74258 10831
rect -73474 10797 -73384 10831
rect -74372 10721 -73384 10797
rect -74372 10687 -74258 10721
rect -73474 10687 -73384 10721
rect -77772 9159 -77574 9193
rect -76790 9159 -76774 9193
rect -76024 9159 -75916 9193
rect -75132 9159 -75036 9193
rect -77772 9085 -76784 9159
rect -76024 9085 -75036 9159
rect -77772 9051 -77574 9085
rect -76790 9051 -76774 9085
rect -76024 9051 -75916 9085
rect -75132 9051 -75036 9085
rect -79330 7523 -79232 7557
rect -78448 7523 -78342 7557
rect -79330 7449 -78342 7523
rect -79330 7415 -79232 7449
rect -78448 7415 -78342 7449
rect -81030 5887 -80890 5921
rect -80106 5887 -80042 5921
rect -81030 5813 -80042 5887
rect -81030 5779 -80890 5813
rect -80106 5779 -80042 5813
rect -82682 4251 -82548 4285
rect -81764 4251 -81694 4285
rect -82682 4220 -81694 4251
rect -81030 4285 -80042 5779
rect -79330 5921 -78342 7415
rect -77772 7557 -76784 9051
rect -76024 7557 -75036 9051
rect -74372 9193 -73384 10687
rect -72742 10831 -71754 12325
rect -71064 12467 -70076 13961
rect -69366 14103 -68378 15597
rect -67736 15739 -66748 17233
rect -66060 17485 -65072 18979
rect -64408 19121 -63420 20615
rect -62778 20649 -61790 20910
rect -62778 20615 -62654 20649
rect -61870 20615 -61790 20649
rect -64408 19087 -64312 19121
rect -63528 19087 -63420 19121
rect -64408 19013 -63420 19087
rect -64408 18979 -64312 19013
rect -63528 18979 -63420 19013
rect -66060 17451 -65970 17485
rect -65186 17451 -65072 17485
rect -66060 17267 -65072 17451
rect -66060 17233 -65968 17267
rect -65184 17233 -65072 17267
rect -67736 15705 -67626 15739
rect -66842 15705 -66748 15739
rect -67736 15631 -66748 15705
rect -67736 15597 -67626 15631
rect -66842 15597 -66748 15631
rect -69366 14069 -69284 14103
rect -68500 14069 -68378 14103
rect -69366 13995 -68378 14069
rect -69366 13961 -69284 13995
rect -68500 13961 -68378 13995
rect -71064 12433 -70942 12467
rect -70158 12433 -70076 12467
rect -71064 12359 -70076 12433
rect -71064 12325 -70942 12359
rect -70158 12325 -70076 12359
rect -72742 10797 -72600 10831
rect -71816 10797 -71754 10831
rect -72742 10721 -71754 10797
rect -72742 10687 -72600 10721
rect -71816 10687 -71754 10721
rect -74372 9159 -74258 9193
rect -73474 9159 -73384 9193
rect -74372 9085 -73384 9159
rect -74372 9051 -74258 9085
rect -73474 9051 -73384 9085
rect -77772 7523 -77574 7557
rect -76790 7523 -76774 7557
rect -76024 7523 -75916 7557
rect -75132 7523 -75036 7557
rect -77772 7449 -76784 7523
rect -76024 7449 -75036 7523
rect -77772 7415 -77574 7449
rect -76790 7415 -76774 7449
rect -76024 7415 -75916 7449
rect -75132 7415 -75036 7449
rect -79330 5887 -79232 5921
rect -78448 5887 -78342 5921
rect -79330 5813 -78342 5887
rect -79330 5779 -79232 5813
rect -78448 5779 -78342 5813
rect -81030 4251 -80890 4285
rect -80106 4251 -80042 4285
rect -81030 4220 -80042 4251
rect -79330 4285 -78342 5779
rect -77772 5921 -76784 7415
rect -76024 5921 -75036 7415
rect -74372 7557 -73384 9051
rect -72742 9193 -71754 10687
rect -71064 10831 -70076 12325
rect -69366 12467 -68378 13961
rect -67736 14103 -66748 15597
rect -66060 15739 -65072 17233
rect -64408 17485 -63420 18979
rect -62778 19121 -61790 20615
rect -61056 20649 -60068 20910
rect -61056 20615 -60996 20649
rect -60212 20615 -60068 20649
rect -62778 19087 -62654 19121
rect -61870 19087 -61790 19121
rect -62778 19013 -61790 19087
rect -62778 18979 -62654 19013
rect -61870 18979 -61790 19013
rect -64408 17451 -64312 17485
rect -63528 17451 -63420 17485
rect -64408 17267 -63420 17451
rect -64408 17233 -64310 17267
rect -63526 17233 -63420 17267
rect -66060 15705 -65968 15739
rect -65184 15705 -65072 15739
rect -66060 15631 -65072 15705
rect -66060 15597 -65968 15631
rect -65184 15597 -65072 15631
rect -67736 14069 -67626 14103
rect -66842 14069 -66748 14103
rect -67736 13995 -66748 14069
rect -67736 13961 -67626 13995
rect -66842 13961 -66748 13995
rect -69366 12433 -69284 12467
rect -68500 12433 -68378 12467
rect -69366 12359 -68378 12433
rect -69366 12325 -69284 12359
rect -68500 12325 -68378 12359
rect -71064 10797 -70942 10831
rect -70158 10797 -70076 10831
rect -71064 10721 -70076 10797
rect -71064 10687 -70942 10721
rect -70158 10687 -70076 10721
rect -72742 9159 -72600 9193
rect -71816 9159 -71754 9193
rect -72742 9085 -71754 9159
rect -72742 9051 -72600 9085
rect -71816 9051 -71754 9085
rect -74372 7523 -74258 7557
rect -73474 7523 -73384 7557
rect -74372 7449 -73384 7523
rect -74372 7415 -74258 7449
rect -73474 7415 -73384 7449
rect -77772 5887 -77574 5921
rect -76790 5887 -76774 5921
rect -76024 5887 -75916 5921
rect -75132 5887 -75036 5921
rect -77772 5813 -76784 5887
rect -76024 5813 -75036 5887
rect -77772 5779 -77574 5813
rect -76790 5779 -76774 5813
rect -76024 5779 -75916 5813
rect -75132 5779 -75036 5813
rect -79330 4251 -79232 4285
rect -78448 4251 -78342 4285
rect -79330 4220 -78342 4251
rect -77772 4285 -76784 5779
rect -76024 4285 -75036 5779
rect -74372 5921 -73384 7415
rect -72742 7557 -71754 9051
rect -71064 9193 -70076 10687
rect -69366 10831 -68378 12325
rect -67736 12467 -66748 13961
rect -66060 14103 -65072 15597
rect -64408 15739 -63420 17233
rect -62778 17485 -61790 18979
rect -61056 19121 -60068 20615
rect -59450 20649 -58462 20910
rect -59450 20615 -59338 20649
rect -58554 20615 -58462 20649
rect -61056 19087 -60996 19121
rect -60212 19087 -60068 19121
rect -61056 19013 -60068 19087
rect -61056 18979 -60996 19013
rect -60212 18979 -60068 19013
rect -62778 17451 -62654 17485
rect -61870 17451 -61790 17485
rect -62778 17267 -61790 17451
rect -62778 17233 -62652 17267
rect -61868 17233 -61790 17267
rect -64408 15705 -64310 15739
rect -63526 15705 -63420 15739
rect -64408 15631 -63420 15705
rect -64408 15597 -64310 15631
rect -63526 15597 -63420 15631
rect -66060 14069 -65968 14103
rect -65184 14069 -65072 14103
rect -66060 13995 -65072 14069
rect -66060 13961 -65968 13995
rect -65184 13961 -65072 13995
rect -67736 12433 -67626 12467
rect -66842 12433 -66748 12467
rect -67736 12359 -66748 12433
rect -67736 12325 -67626 12359
rect -66842 12325 -66748 12359
rect -69366 10797 -69284 10831
rect -68500 10797 -68378 10831
rect -69366 10721 -68378 10797
rect -69366 10687 -69284 10721
rect -68500 10687 -68378 10721
rect -71064 9159 -70942 9193
rect -70158 9159 -70076 9193
rect -71064 9085 -70076 9159
rect -71064 9051 -70942 9085
rect -70158 9051 -70076 9085
rect -72742 7523 -72600 7557
rect -71816 7523 -71754 7557
rect -72742 7449 -71754 7523
rect -72742 7415 -72600 7449
rect -71816 7415 -71754 7449
rect -74372 5887 -74258 5921
rect -73474 5887 -73384 5921
rect -74372 5813 -73384 5887
rect -74372 5779 -74258 5813
rect -73474 5779 -73384 5813
rect -77772 4251 -77574 4285
rect -76790 4251 -76774 4285
rect -77772 4220 -76774 4251
rect -76024 4251 -75916 4285
rect -75132 4251 -75036 4285
rect -76024 4220 -75036 4251
rect -74372 4285 -73384 5779
rect -72742 5921 -71754 7415
rect -71064 7557 -70076 9051
rect -69366 9193 -68378 10687
rect -67736 10831 -66748 12325
rect -66060 12467 -65072 13961
rect -64408 14103 -63420 15597
rect -62778 15739 -61790 17233
rect -61056 17485 -60068 18979
rect -59450 19121 -58462 20615
rect -57750 20649 -56762 20910
rect -57750 20615 -57680 20649
rect -56896 20615 -56762 20649
rect -59450 19087 -59338 19121
rect -58554 19087 -58462 19121
rect -59450 19013 -58462 19087
rect -59450 18979 -59338 19013
rect -58554 18979 -58462 19013
rect -61056 17451 -60996 17485
rect -60212 17451 -60068 17485
rect -61056 17267 -60068 17451
rect -61056 17233 -60994 17267
rect -60210 17233 -60068 17267
rect -62778 15705 -62652 15739
rect -61868 15705 -61790 15739
rect -62778 15631 -61790 15705
rect -62778 15597 -62652 15631
rect -61868 15597 -61790 15631
rect -64408 14069 -64310 14103
rect -63526 14069 -63420 14103
rect -64408 13995 -63420 14069
rect -64408 13961 -64310 13995
rect -63526 13961 -63420 13995
rect -66060 12433 -65968 12467
rect -65184 12433 -65072 12467
rect -66060 12359 -65072 12433
rect -66060 12325 -65968 12359
rect -65184 12325 -65072 12359
rect -67736 10797 -67626 10831
rect -66842 10797 -66748 10831
rect -67736 10721 -66748 10797
rect -67736 10687 -67626 10721
rect -66842 10687 -66748 10721
rect -69366 9159 -69284 9193
rect -68500 9159 -68378 9193
rect -69366 9085 -68378 9159
rect -69366 9051 -69284 9085
rect -68500 9051 -68378 9085
rect -71064 7523 -70942 7557
rect -70158 7523 -70076 7557
rect -71064 7449 -70076 7523
rect -71064 7415 -70942 7449
rect -70158 7415 -70076 7449
rect -72742 5887 -72600 5921
rect -71816 5887 -71754 5921
rect -72742 5813 -71754 5887
rect -72742 5779 -72600 5813
rect -71816 5779 -71754 5813
rect -74372 4251 -74258 4285
rect -73474 4251 -73384 4285
rect -74372 4220 -73384 4251
rect -72742 4285 -71754 5779
rect -71064 5921 -70076 7415
rect -69366 7557 -68378 9051
rect -67736 9193 -66748 10687
rect -66060 10831 -65072 12325
rect -64408 12467 -63420 13961
rect -62778 14103 -61790 15597
rect -61056 15739 -60068 17233
rect -59450 17485 -58462 18979
rect -57750 19121 -56762 20615
rect -56074 20649 -55086 20910
rect -56074 20615 -56022 20649
rect -55238 20615 -55086 20649
rect -57750 19087 -57680 19121
rect -56896 19087 -56762 19121
rect -57750 19013 -56762 19087
rect -57750 18979 -57680 19013
rect -56896 18979 -56762 19013
rect -59450 17451 -59338 17485
rect -58554 17451 -58462 17485
rect -59450 17267 -58462 17451
rect -59450 17233 -59336 17267
rect -58552 17233 -58462 17267
rect -61056 15705 -60994 15739
rect -60210 15705 -60068 15739
rect -61056 15631 -60068 15705
rect -61056 15597 -60994 15631
rect -60210 15597 -60068 15631
rect -62778 14069 -62652 14103
rect -61868 14069 -61790 14103
rect -62778 13995 -61790 14069
rect -62778 13961 -62652 13995
rect -61868 13961 -61790 13995
rect -64408 12433 -64310 12467
rect -63526 12433 -63420 12467
rect -64408 12359 -63420 12433
rect -64408 12325 -64310 12359
rect -63526 12325 -63420 12359
rect -66060 10797 -65968 10831
rect -65184 10797 -65072 10831
rect -66060 10721 -65072 10797
rect -66060 10687 -65968 10721
rect -65184 10687 -65072 10721
rect -67736 9159 -67626 9193
rect -66842 9159 -66748 9193
rect -67736 9085 -66748 9159
rect -67736 9051 -67626 9085
rect -66842 9051 -66748 9085
rect -69366 7523 -69284 7557
rect -68500 7523 -68378 7557
rect -69366 7449 -68378 7523
rect -69366 7415 -69284 7449
rect -68500 7415 -68378 7449
rect -71064 5887 -70942 5921
rect -70158 5887 -70076 5921
rect -71064 5813 -70076 5887
rect -71064 5779 -70942 5813
rect -70158 5779 -70076 5813
rect -72742 4251 -72600 4285
rect -71816 4251 -71754 4285
rect -72742 4220 -71754 4251
rect -71064 4285 -70076 5779
rect -69366 5921 -68378 7415
rect -67736 7557 -66748 9051
rect -66060 9193 -65072 10687
rect -64408 10831 -63420 12325
rect -62778 12467 -61790 13961
rect -61056 14103 -60068 15597
rect -59450 15739 -58462 17233
rect -57750 17485 -56762 18979
rect -56074 19121 -55086 20615
rect -54444 20649 -53456 20886
rect -54444 20615 -54364 20649
rect -53580 20615 -53456 20649
rect -56074 19087 -56022 19121
rect -55238 19087 -55086 19121
rect -56074 19013 -55086 19087
rect -56074 18979 -56022 19013
rect -55238 18979 -55086 19013
rect -57750 17451 -57680 17485
rect -56896 17451 -56762 17485
rect -57750 17267 -56762 17451
rect -57750 17233 -57678 17267
rect -56894 17233 -56762 17267
rect -59450 15705 -59336 15739
rect -58552 15705 -58462 15739
rect -59450 15631 -58462 15705
rect -59450 15597 -59336 15631
rect -58552 15597 -58462 15631
rect -61056 14069 -60994 14103
rect -60210 14069 -60068 14103
rect -61056 13995 -60068 14069
rect -61056 13961 -60994 13995
rect -60210 13961 -60068 13995
rect -62778 12433 -62652 12467
rect -61868 12433 -61790 12467
rect -62778 12359 -61790 12433
rect -62778 12325 -62652 12359
rect -61868 12325 -61790 12359
rect -64408 10797 -64310 10831
rect -63526 10797 -63420 10831
rect -64408 10721 -63420 10797
rect -64408 10687 -64310 10721
rect -63526 10687 -63420 10721
rect -66060 9159 -65968 9193
rect -65184 9159 -65072 9193
rect -66060 9085 -65072 9159
rect -66060 9051 -65968 9085
rect -65184 9051 -65072 9085
rect -67736 7523 -67626 7557
rect -66842 7523 -66748 7557
rect -67736 7449 -66748 7523
rect -67736 7415 -67626 7449
rect -66842 7415 -66748 7449
rect -69366 5887 -69284 5921
rect -68500 5887 -68378 5921
rect -69366 5813 -68378 5887
rect -69366 5779 -69284 5813
rect -68500 5779 -68378 5813
rect -71064 4251 -70942 4285
rect -70158 4251 -70076 4285
rect -71064 4220 -70076 4251
rect -69366 4285 -68378 5779
rect -67736 5921 -66748 7415
rect -66060 7557 -65072 9051
rect -64408 9193 -63420 10687
rect -62778 10831 -61790 12325
rect -61056 12467 -60068 13961
rect -59450 14103 -58462 15597
rect -57750 15739 -56762 17233
rect -56074 17485 -55086 18979
rect -54444 19121 -53456 20615
rect -52816 20649 -51828 20910
rect -52816 20615 -52706 20649
rect -51922 20615 -51828 20649
rect -54444 19087 -54364 19121
rect -53580 19087 -53456 19121
rect -54444 19013 -53456 19087
rect -54444 18979 -54364 19013
rect -53580 18979 -53456 19013
rect -56074 17451 -56022 17485
rect -55238 17451 -55086 17485
rect -56074 17267 -55086 17451
rect -56074 17233 -56020 17267
rect -55236 17233 -55086 17267
rect -57750 15705 -57678 15739
rect -56894 15705 -56762 15739
rect -57750 15631 -56762 15705
rect -57750 15597 -57678 15631
rect -56894 15597 -56762 15631
rect -59450 14069 -59336 14103
rect -58552 14069 -58462 14103
rect -59450 13995 -58462 14069
rect -59450 13961 -59336 13995
rect -58552 13961 -58462 13995
rect -61056 12433 -60994 12467
rect -60210 12433 -60068 12467
rect -61056 12359 -60068 12433
rect -61056 12325 -60994 12359
rect -60210 12325 -60068 12359
rect -62778 10797 -62652 10831
rect -61868 10797 -61790 10831
rect -62778 10721 -61790 10797
rect -62778 10687 -62652 10721
rect -61868 10687 -61790 10721
rect -64408 9159 -64310 9193
rect -63526 9159 -63420 9193
rect -64408 9085 -63420 9159
rect -64408 9051 -64310 9085
rect -63526 9051 -63420 9085
rect -66060 7523 -65968 7557
rect -65184 7523 -65072 7557
rect -66060 7449 -65072 7523
rect -66060 7415 -65968 7449
rect -65184 7415 -65072 7449
rect -67736 5887 -67626 5921
rect -66842 5887 -66748 5921
rect -67736 5813 -66748 5887
rect -67736 5779 -67626 5813
rect -66842 5779 -66748 5813
rect -69366 4251 -69284 4285
rect -68500 4251 -68378 4285
rect -69366 4220 -68378 4251
rect -67736 4285 -66748 5779
rect -66060 5921 -65072 7415
rect -64408 7557 -63420 9051
rect -62778 9193 -61790 10687
rect -61056 10831 -60068 12325
rect -59450 12467 -58462 13961
rect -57750 14103 -56762 15597
rect -56074 15739 -55086 17233
rect -54444 17485 -53456 18979
rect -52816 19121 -51828 20615
rect -51132 20649 -50144 20864
rect -51132 20615 -51048 20649
rect -50264 20615 -50144 20649
rect -52816 19087 -52706 19121
rect -51922 19087 -51828 19121
rect -52816 19013 -51828 19087
rect -52816 18979 -52706 19013
rect -51922 18979 -51828 19013
rect -54444 17451 -54364 17485
rect -53580 17451 -53456 17485
rect -54444 17267 -53456 17451
rect -54444 17233 -54362 17267
rect -53578 17233 -53456 17267
rect -56074 15705 -56020 15739
rect -55236 15705 -55086 15739
rect -56074 15631 -55086 15705
rect -56074 15597 -56020 15631
rect -55236 15597 -55086 15631
rect -57750 14069 -57678 14103
rect -56894 14069 -56762 14103
rect -57750 13995 -56762 14069
rect -57750 13961 -57678 13995
rect -56894 13961 -56762 13995
rect -59450 12433 -59336 12467
rect -58552 12433 -58462 12467
rect -59450 12359 -58462 12433
rect -59450 12325 -59336 12359
rect -58552 12325 -58462 12359
rect -61056 10797 -60994 10831
rect -60210 10797 -60068 10831
rect -61056 10721 -60068 10797
rect -61056 10687 -60994 10721
rect -60210 10687 -60068 10721
rect -62778 9159 -62652 9193
rect -61868 9159 -61790 9193
rect -62778 9085 -61790 9159
rect -62778 9051 -62652 9085
rect -61868 9051 -61790 9085
rect -64408 7523 -64310 7557
rect -63526 7523 -63420 7557
rect -64408 7449 -63420 7523
rect -64408 7415 -64310 7449
rect -63526 7415 -63420 7449
rect -66060 5887 -65968 5921
rect -65184 5887 -65072 5921
rect -66060 5813 -65072 5887
rect -66060 5779 -65968 5813
rect -65184 5779 -65072 5813
rect -67736 4251 -67626 4285
rect -66842 4251 -66748 4285
rect -67736 4220 -66748 4251
rect -66060 4285 -65072 5779
rect -64408 5921 -63420 7415
rect -62778 7557 -61790 9051
rect -61056 9193 -60068 10687
rect -59450 10831 -58462 12325
rect -57750 12467 -56762 13961
rect -56074 14103 -55086 15597
rect -54444 15739 -53456 17233
rect -52816 17485 -51828 18979
rect -51132 19121 -50144 20615
rect -49458 20649 -48470 20880
rect -49458 20615 -49390 20649
rect -48606 20615 -48470 20649
rect -51132 19087 -51048 19121
rect -50264 19087 -50144 19121
rect -51132 19013 -50144 19087
rect -51132 18979 -51048 19013
rect -50264 18979 -50144 19013
rect -52816 17451 -52706 17485
rect -51922 17451 -51828 17485
rect -52816 17267 -51828 17451
rect -52816 17233 -52704 17267
rect -51920 17233 -51828 17267
rect -54444 15705 -54362 15739
rect -53578 15705 -53456 15739
rect -54444 15631 -53456 15705
rect -54444 15597 -54362 15631
rect -53578 15597 -53456 15631
rect -56074 14069 -56020 14103
rect -55236 14069 -55086 14103
rect -56074 13995 -55086 14069
rect -56074 13961 -56020 13995
rect -55236 13961 -55086 13995
rect -57750 12433 -57678 12467
rect -56894 12433 -56762 12467
rect -57750 12359 -56762 12433
rect -57750 12325 -57678 12359
rect -56894 12325 -56762 12359
rect -59450 10797 -59336 10831
rect -58552 10797 -58462 10831
rect -59450 10721 -58462 10797
rect -59450 10687 -59336 10721
rect -58552 10687 -58462 10721
rect -61056 9159 -60994 9193
rect -60210 9159 -60068 9193
rect -61056 9085 -60068 9159
rect -61056 9051 -60994 9085
rect -60210 9051 -60068 9085
rect -62778 7523 -62652 7557
rect -61868 7523 -61790 7557
rect -62778 7449 -61790 7523
rect -62778 7415 -62652 7449
rect -61868 7415 -61790 7449
rect -64408 5887 -64310 5921
rect -63526 5887 -63420 5921
rect -64408 5813 -63420 5887
rect -64408 5779 -64310 5813
rect -63526 5779 -63420 5813
rect -66060 4251 -65968 4285
rect -65184 4251 -65072 4285
rect -66060 4220 -65072 4251
rect -64408 4285 -63420 5779
rect -62778 5921 -61790 7415
rect -61056 7557 -60068 9051
rect -59450 9193 -58462 10687
rect -57750 10831 -56762 12325
rect -56074 12467 -55086 13961
rect -54444 14103 -53456 15597
rect -52816 15739 -51828 17233
rect -51132 17485 -50144 18979
rect -49458 19121 -48470 20615
rect -47808 20649 -46820 20904
rect -47808 20615 -47732 20649
rect -46948 20615 -46820 20649
rect -49458 19087 -49390 19121
rect -48606 19087 -48470 19121
rect -49458 19013 -48470 19087
rect -49458 18979 -49390 19013
rect -48606 18979 -48470 19013
rect -51132 17451 -51048 17485
rect -50264 17451 -50144 17485
rect -51132 17267 -50144 17451
rect -51132 17233 -51046 17267
rect -50262 17233 -50144 17267
rect -52816 15705 -52704 15739
rect -51920 15705 -51828 15739
rect -52816 15631 -51828 15705
rect -52816 15597 -52704 15631
rect -51920 15597 -51828 15631
rect -54444 14069 -54362 14103
rect -53578 14069 -53456 14103
rect -54444 13995 -53456 14069
rect -54444 13961 -54362 13995
rect -53578 13961 -53456 13995
rect -56074 12433 -56020 12467
rect -55236 12433 -55086 12467
rect -56074 12359 -55086 12433
rect -56074 12325 -56020 12359
rect -55236 12325 -55086 12359
rect -57750 10797 -57678 10831
rect -56894 10797 -56762 10831
rect -57750 10721 -56762 10797
rect -57750 10687 -57678 10721
rect -56894 10687 -56762 10721
rect -59450 9159 -59336 9193
rect -58552 9159 -58462 9193
rect -59450 9085 -58462 9159
rect -59450 9051 -59336 9085
rect -58552 9051 -58462 9085
rect -61056 7523 -60994 7557
rect -60210 7523 -60068 7557
rect -61056 7449 -60068 7523
rect -61056 7415 -60994 7449
rect -60210 7415 -60068 7449
rect -62778 5887 -62652 5921
rect -61868 5887 -61790 5921
rect -62778 5813 -61790 5887
rect -62778 5779 -62652 5813
rect -61868 5779 -61790 5813
rect -64408 4251 -64310 4285
rect -63526 4251 -63420 4285
rect -64408 4220 -63420 4251
rect -62778 4285 -61790 5779
rect -61056 5921 -60068 7415
rect -59450 7557 -58462 9051
rect -57750 9193 -56762 10687
rect -56074 10831 -55086 12325
rect -54444 12467 -53456 13961
rect -52816 14103 -51828 15597
rect -51132 15739 -50144 17233
rect -49458 17485 -48470 18979
rect -47808 19121 -46820 20615
rect -46202 20649 -45214 20880
rect -46202 20615 -46074 20649
rect -45290 20615 -45214 20649
rect -47808 19087 -47732 19121
rect -46948 19087 -46820 19121
rect -47808 19013 -46820 19087
rect -47808 18979 -47732 19013
rect -46948 18979 -46820 19013
rect -49458 17451 -49390 17485
rect -48606 17451 -48470 17485
rect -49458 17267 -48470 17451
rect -49458 17233 -49388 17267
rect -48604 17233 -48470 17267
rect -51132 15705 -51046 15739
rect -50262 15705 -50144 15739
rect -51132 15631 -50144 15705
rect -51132 15597 -51046 15631
rect -50262 15597 -50144 15631
rect -52816 14069 -52704 14103
rect -51920 14069 -51828 14103
rect -52816 13995 -51828 14069
rect -52816 13961 -52704 13995
rect -51920 13961 -51828 13995
rect -54444 12433 -54362 12467
rect -53578 12433 -53456 12467
rect -54444 12359 -53456 12433
rect -54444 12325 -54362 12359
rect -53578 12325 -53456 12359
rect -56074 10797 -56020 10831
rect -55236 10797 -55086 10831
rect -56074 10721 -55086 10797
rect -56074 10687 -56020 10721
rect -55236 10687 -55086 10721
rect -57750 9159 -57678 9193
rect -56894 9159 -56762 9193
rect -57750 9085 -56762 9159
rect -57750 9051 -57678 9085
rect -56894 9051 -56762 9085
rect -59450 7523 -59336 7557
rect -58552 7523 -58462 7557
rect -59450 7449 -58462 7523
rect -59450 7415 -59336 7449
rect -58552 7415 -58462 7449
rect -61056 5887 -60994 5921
rect -60210 5887 -60068 5921
rect -61056 5813 -60068 5887
rect -61056 5779 -60994 5813
rect -60210 5779 -60068 5813
rect -61056 4306 -60068 5779
rect -59450 5921 -58462 7415
rect -57750 7557 -56762 9051
rect -56074 9193 -55086 10687
rect -54444 10831 -53456 12325
rect -52816 12467 -51828 13961
rect -51132 14103 -50144 15597
rect -49458 15739 -48470 17233
rect -47808 17485 -46820 18979
rect -46202 19121 -45214 20615
rect -44504 20649 -43516 20904
rect -44504 20615 -44416 20649
rect -43632 20615 -43516 20649
rect -46202 19087 -46074 19121
rect -45290 19087 -45214 19121
rect -46202 19013 -45214 19087
rect -46202 18979 -46074 19013
rect -45290 18979 -45214 19013
rect -47808 17451 -47732 17485
rect -46948 17451 -46820 17485
rect -47808 17267 -46820 17451
rect -47808 17233 -47730 17267
rect -46946 17233 -46820 17267
rect -49458 15705 -49388 15739
rect -48604 15705 -48470 15739
rect -49458 15631 -48470 15705
rect -49458 15597 -49388 15631
rect -48604 15597 -48470 15631
rect -51132 14069 -51046 14103
rect -50262 14069 -50144 14103
rect -51132 13995 -50144 14069
rect -51132 13961 -51046 13995
rect -50262 13961 -50144 13995
rect -52816 12433 -52704 12467
rect -51920 12433 -51828 12467
rect -52816 12359 -51828 12433
rect -52816 12325 -52704 12359
rect -51920 12325 -51828 12359
rect -54444 10797 -54362 10831
rect -53578 10797 -53456 10831
rect -54444 10721 -53456 10797
rect -54444 10687 -54362 10721
rect -53578 10687 -53456 10721
rect -56074 9159 -56020 9193
rect -55236 9159 -55086 9193
rect -56074 9085 -55086 9159
rect -56074 9051 -56020 9085
rect -55236 9051 -55086 9085
rect -57750 7523 -57678 7557
rect -56894 7523 -56762 7557
rect -57750 7449 -56762 7523
rect -57750 7415 -57678 7449
rect -56894 7415 -56762 7449
rect -59450 5887 -59336 5921
rect -58552 5887 -58462 5921
rect -59450 5813 -58462 5887
rect -59450 5779 -59336 5813
rect -58552 5779 -58462 5813
rect -62778 4251 -62652 4285
rect -61868 4251 -61790 4285
rect -62778 4220 -61790 4251
rect -94232 4182 -61790 4220
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -62542 4086 -61790 4182
rect -61050 4285 -60068 4306
rect -61050 4264 -60994 4285
rect -61050 4230 -61008 4264
rect -60210 4251 -60068 4285
rect -60974 4236 -60068 4251
rect -59450 4285 -58462 5779
rect -57750 5921 -56762 7415
rect -56074 7557 -55086 9051
rect -54444 9193 -53456 10687
rect -52816 10831 -51828 12325
rect -51132 12467 -50144 13961
rect -49458 14103 -48470 15597
rect -47808 15739 -46820 17233
rect -46202 17485 -45214 18979
rect -44504 19121 -43516 20615
rect -42852 20649 -41864 20880
rect -42852 20615 -42758 20649
rect -41974 20615 -41864 20649
rect -44504 19087 -44416 19121
rect -43632 19087 -43516 19121
rect -44504 19013 -43516 19087
rect -44504 18979 -44416 19013
rect -43632 18979 -43516 19013
rect -46202 17451 -46074 17485
rect -45290 17451 -45214 17485
rect -46202 17267 -45214 17451
rect -46202 17233 -46072 17267
rect -45288 17233 -45214 17267
rect -47808 15705 -47730 15739
rect -46946 15705 -46820 15739
rect -47808 15631 -46820 15705
rect -47808 15597 -47730 15631
rect -46946 15597 -46820 15631
rect -49458 14069 -49388 14103
rect -48604 14069 -48470 14103
rect -49458 13995 -48470 14069
rect -49458 13961 -49388 13995
rect -48604 13961 -48470 13995
rect -51132 12433 -51046 12467
rect -50262 12433 -50144 12467
rect -51132 12359 -50144 12433
rect -51132 12325 -51046 12359
rect -50262 12325 -50144 12359
rect -52816 10797 -52704 10831
rect -51920 10797 -51828 10831
rect -52816 10721 -51828 10797
rect -52816 10687 -52704 10721
rect -51920 10687 -51828 10721
rect -54444 9159 -54362 9193
rect -53578 9159 -53456 9193
rect -54444 9085 -53456 9159
rect -54444 9051 -54362 9085
rect -53578 9051 -53456 9085
rect -56074 7523 -56020 7557
rect -55236 7523 -55086 7557
rect -56074 7449 -55086 7523
rect -56074 7415 -56020 7449
rect -55236 7415 -55086 7449
rect -57750 5887 -57678 5921
rect -56894 5887 -56762 5921
rect -57750 5813 -56762 5887
rect -57750 5779 -57678 5813
rect -56894 5779 -56762 5813
rect -59450 4251 -59336 4285
rect -58552 4251 -58462 4285
rect -59450 4236 -58462 4251
rect -57750 4285 -56762 5779
rect -56074 5921 -55086 7415
rect -54444 7557 -53456 9051
rect -52816 9193 -51828 10687
rect -51132 10831 -50144 12325
rect -49458 12467 -48470 13961
rect -47808 14103 -46820 15597
rect -46202 15739 -45214 17233
rect -44504 17485 -43516 18979
rect -42852 19121 -41864 20615
rect -41202 20649 -40214 20904
rect -41202 20615 -41100 20649
rect -40316 20615 -40214 20649
rect -42852 19087 -42758 19121
rect -41974 19087 -41864 19121
rect -42852 19013 -41864 19087
rect -42852 18979 -42758 19013
rect -41974 18979 -41864 19013
rect -44504 17451 -44416 17485
rect -43632 17451 -43516 17485
rect -44504 17267 -43516 17451
rect -44504 17233 -44414 17267
rect -43630 17233 -43516 17267
rect -46202 15705 -46072 15739
rect -45288 15705 -45214 15739
rect -46202 15631 -45214 15705
rect -46202 15597 -46072 15631
rect -45288 15597 -45214 15631
rect -47808 14069 -47730 14103
rect -46946 14069 -46820 14103
rect -47808 13995 -46820 14069
rect -47808 13961 -47730 13995
rect -46946 13961 -46820 13995
rect -49458 12433 -49388 12467
rect -48604 12433 -48470 12467
rect -49458 12359 -48470 12433
rect -49458 12325 -49388 12359
rect -48604 12325 -48470 12359
rect -51132 10797 -51046 10831
rect -50262 10797 -50144 10831
rect -51132 10721 -50144 10797
rect -51132 10687 -51046 10721
rect -50262 10687 -50144 10721
rect -52816 9159 -52704 9193
rect -51920 9159 -51828 9193
rect -52816 9085 -51828 9159
rect -52816 9051 -52704 9085
rect -51920 9051 -51828 9085
rect -54444 7523 -54362 7557
rect -53578 7523 -53456 7557
rect -54444 7449 -53456 7523
rect -54444 7415 -54362 7449
rect -53578 7415 -53456 7449
rect -56074 5887 -56020 5921
rect -55236 5887 -55086 5921
rect -56074 5813 -55086 5887
rect -56074 5779 -56020 5813
rect -55236 5779 -55086 5813
rect -57750 4251 -57678 4285
rect -56894 4251 -56762 4285
rect -57750 4236 -56762 4251
rect -56074 4285 -55086 5779
rect -54444 5921 -53456 7415
rect -52816 7557 -51828 9051
rect -51132 9193 -50144 10687
rect -49458 10831 -48470 12325
rect -47808 12467 -46820 13961
rect -46202 14103 -45214 15597
rect -44504 15739 -43516 17233
rect -42852 17485 -41864 18979
rect -41202 19121 -40214 20615
rect -39550 20649 -38562 20880
rect -39550 20615 -39442 20649
rect -38658 20615 -38562 20649
rect -41202 19087 -41100 19121
rect -40316 19087 -40214 19121
rect -41202 19013 -40214 19087
rect -41202 18979 -41100 19013
rect -40316 18979 -40214 19013
rect -42852 17451 -42758 17485
rect -41974 17451 -41864 17485
rect -42852 17267 -41864 17451
rect -42852 17233 -42756 17267
rect -41972 17233 -41864 17267
rect -44504 15705 -44414 15739
rect -43630 15705 -43516 15739
rect -44504 15631 -43516 15705
rect -44504 15597 -44414 15631
rect -43630 15597 -43516 15631
rect -46202 14069 -46072 14103
rect -45288 14069 -45214 14103
rect -46202 13995 -45214 14069
rect -46202 13961 -46072 13995
rect -45288 13961 -45214 13995
rect -47808 12433 -47730 12467
rect -46946 12433 -46820 12467
rect -47808 12359 -46820 12433
rect -47808 12325 -47730 12359
rect -46946 12325 -46820 12359
rect -49458 10797 -49388 10831
rect -48604 10797 -48470 10831
rect -49458 10721 -48470 10797
rect -49458 10687 -49388 10721
rect -48604 10687 -48470 10721
rect -51132 9159 -51046 9193
rect -50262 9159 -50144 9193
rect -51132 9085 -50144 9159
rect -51132 9051 -51046 9085
rect -50262 9051 -50144 9085
rect -52816 7523 -52704 7557
rect -51920 7523 -51828 7557
rect -52816 7449 -51828 7523
rect -52816 7415 -52704 7449
rect -51920 7415 -51828 7449
rect -54444 5887 -54362 5921
rect -53578 5887 -53456 5921
rect -54444 5813 -53456 5887
rect -54444 5779 -54362 5813
rect -53578 5779 -53456 5813
rect -56074 4251 -56020 4285
rect -55236 4251 -55086 4285
rect -56074 4236 -55086 4251
rect -54444 4285 -53456 5779
rect -52816 5921 -51828 7415
rect -51132 7557 -50144 9051
rect -49458 9193 -48470 10687
rect -47808 10831 -46820 12325
rect -46202 12467 -45214 13961
rect -44504 14103 -43516 15597
rect -42852 15739 -41864 17233
rect -41202 17485 -40214 18979
rect -39550 19121 -38562 20615
rect -37892 20649 -36904 20882
rect -37892 20615 -37784 20649
rect -37000 20615 -36904 20649
rect -39550 19087 -39442 19121
rect -38658 19087 -38562 19121
rect -39550 19013 -38562 19087
rect -39550 18979 -39442 19013
rect -38658 18979 -38562 19013
rect -41202 17451 -41100 17485
rect -40316 17451 -40214 17485
rect -41202 17267 -40214 17451
rect -41202 17233 -41098 17267
rect -40314 17233 -40214 17267
rect -42852 15705 -42756 15739
rect -41972 15705 -41864 15739
rect -42852 15631 -41864 15705
rect -42852 15597 -42756 15631
rect -41972 15597 -41864 15631
rect -44504 14069 -44414 14103
rect -43630 14069 -43516 14103
rect -44504 13995 -43516 14069
rect -44504 13961 -44414 13995
rect -43630 13961 -43516 13995
rect -46202 12433 -46072 12467
rect -45288 12433 -45214 12467
rect -46202 12359 -45214 12433
rect -46202 12325 -46072 12359
rect -45288 12325 -45214 12359
rect -47808 10797 -47730 10831
rect -46946 10797 -46820 10831
rect -47808 10721 -46820 10797
rect -47808 10687 -47730 10721
rect -46946 10687 -46820 10721
rect -49458 9159 -49388 9193
rect -48604 9159 -48470 9193
rect -49458 9085 -48470 9159
rect -49458 9051 -49388 9085
rect -48604 9051 -48470 9085
rect -51132 7523 -51046 7557
rect -50262 7523 -50144 7557
rect -51132 7449 -50144 7523
rect -51132 7415 -51046 7449
rect -50262 7415 -50144 7449
rect -52816 5887 -52704 5921
rect -51920 5887 -51828 5921
rect -52816 5813 -51828 5887
rect -52816 5779 -52704 5813
rect -51920 5779 -51828 5813
rect -54444 4251 -54362 4285
rect -53578 4251 -53456 4285
rect -54444 4236 -53456 4251
rect -52816 4285 -51828 5779
rect -51132 5921 -50144 7415
rect -49458 7557 -48470 9051
rect -47808 9193 -46820 10687
rect -46202 10831 -45214 12325
rect -44504 12467 -43516 13961
rect -42852 14103 -41864 15597
rect -41202 15739 -40214 17233
rect -39550 17485 -38562 18979
rect -37892 19121 -36904 20615
rect -36244 20649 -35256 20882
rect -36244 20615 -36126 20649
rect -35342 20615 -35256 20649
rect -37892 19087 -37784 19121
rect -37000 19087 -36904 19121
rect -37892 19013 -36904 19087
rect -37892 18979 -37784 19013
rect -37000 18979 -36904 19013
rect -39550 17451 -39442 17485
rect -38658 17451 -38562 17485
rect -39550 17267 -38562 17451
rect -39550 17233 -39440 17267
rect -38656 17233 -38562 17267
rect -41202 15705 -41098 15739
rect -40314 15705 -40214 15739
rect -41202 15631 -40214 15705
rect -41202 15597 -41098 15631
rect -40314 15597 -40214 15631
rect -42852 14069 -42756 14103
rect -41972 14069 -41864 14103
rect -42852 13995 -41864 14069
rect -42852 13961 -42756 13995
rect -41972 13961 -41864 13995
rect -44504 12433 -44414 12467
rect -43630 12433 -43516 12467
rect -44504 12359 -43516 12433
rect -44504 12325 -44414 12359
rect -43630 12325 -43516 12359
rect -46202 10797 -46072 10831
rect -45288 10797 -45214 10831
rect -46202 10721 -45214 10797
rect -46202 10687 -46072 10721
rect -45288 10687 -45214 10721
rect -47808 9159 -47730 9193
rect -46946 9159 -46820 9193
rect -47808 9085 -46820 9159
rect -47808 9051 -47730 9085
rect -46946 9051 -46820 9085
rect -49458 7523 -49388 7557
rect -48604 7523 -48470 7557
rect -49458 7449 -48470 7523
rect -49458 7415 -49388 7449
rect -48604 7415 -48470 7449
rect -51132 5887 -51046 5921
rect -50262 5887 -50144 5921
rect -51132 5813 -50144 5887
rect -51132 5779 -51046 5813
rect -50262 5779 -50144 5813
rect -52816 4251 -52704 4285
rect -51920 4251 -51828 4285
rect -52816 4236 -51828 4251
rect -51132 4285 -50144 5779
rect -49458 5921 -48470 7415
rect -47808 7557 -46820 9051
rect -46202 9193 -45214 10687
rect -44504 10831 -43516 12325
rect -42852 12467 -41864 13961
rect -41202 14103 -40214 15597
rect -39550 15739 -38562 17233
rect -37892 17485 -36904 18979
rect -36244 19121 -35256 20615
rect -34550 20649 -33562 20882
rect -34550 20615 -34468 20649
rect -33684 20615 -33562 20649
rect -36244 19087 -36126 19121
rect -35342 19087 -35256 19121
rect -36244 19013 -35256 19087
rect -36244 18979 -36126 19013
rect -35342 18979 -35256 19013
rect -37892 17451 -37784 17485
rect -37000 17451 -36904 17485
rect -37892 17267 -36904 17451
rect -37892 17233 -37782 17267
rect -36998 17233 -36904 17267
rect -39550 15705 -39440 15739
rect -38656 15705 -38562 15739
rect -39550 15631 -38562 15705
rect -39550 15597 -39440 15631
rect -38656 15597 -38562 15631
rect -41202 14069 -41098 14103
rect -40314 14069 -40214 14103
rect -41202 13995 -40214 14069
rect -41202 13961 -41098 13995
rect -40314 13961 -40214 13995
rect -42852 12433 -42756 12467
rect -41972 12433 -41864 12467
rect -42852 12359 -41864 12433
rect -42852 12325 -42756 12359
rect -41972 12325 -41864 12359
rect -44504 10797 -44414 10831
rect -43630 10797 -43516 10831
rect -44504 10721 -43516 10797
rect -44504 10687 -44414 10721
rect -43630 10687 -43516 10721
rect -46202 9159 -46072 9193
rect -45288 9159 -45214 9193
rect -46202 9085 -45214 9159
rect -46202 9051 -46072 9085
rect -45288 9051 -45214 9085
rect -47808 7523 -47730 7557
rect -46946 7523 -46820 7557
rect -47808 7449 -46820 7523
rect -47808 7415 -47730 7449
rect -46946 7415 -46820 7449
rect -49458 5887 -49388 5921
rect -48604 5887 -48470 5921
rect -49458 5813 -48470 5887
rect -49458 5779 -49388 5813
rect -48604 5779 -48470 5813
rect -51132 4251 -51046 4285
rect -50262 4251 -50144 4285
rect -51132 4236 -50144 4251
rect -49458 4285 -48470 5779
rect -47808 5921 -46820 7415
rect -46202 7557 -45214 9051
rect -44504 9193 -43516 10687
rect -42852 10831 -41864 12325
rect -41202 12467 -40214 13961
rect -39550 14103 -38562 15597
rect -37892 15739 -36904 17233
rect -36244 17485 -35256 18979
rect -34550 19121 -33562 20615
rect -32902 20649 -31914 20930
rect -32902 20615 -32810 20649
rect -32026 20615 -31914 20649
rect -34550 19087 -34468 19121
rect -33684 19087 -33562 19121
rect -34550 19013 -33562 19087
rect -34550 18979 -34468 19013
rect -33684 18979 -33562 19013
rect -36244 17451 -36126 17485
rect -35342 17451 -35256 17485
rect -36244 17267 -35256 17451
rect -36244 17233 -36124 17267
rect -35340 17233 -35256 17267
rect -37892 15705 -37782 15739
rect -36998 15705 -36904 15739
rect -37892 15631 -36904 15705
rect -37892 15597 -37782 15631
rect -36998 15597 -36904 15631
rect -39550 14069 -39440 14103
rect -38656 14069 -38562 14103
rect -39550 13995 -38562 14069
rect -39550 13961 -39440 13995
rect -38656 13961 -38562 13995
rect -41202 12433 -41098 12467
rect -40314 12433 -40214 12467
rect -41202 12359 -40214 12433
rect -41202 12325 -41098 12359
rect -40314 12325 -40214 12359
rect -42852 10797 -42756 10831
rect -41972 10797 -41864 10831
rect -42852 10721 -41864 10797
rect -42852 10687 -42756 10721
rect -41972 10687 -41864 10721
rect -44504 9159 -44414 9193
rect -43630 9159 -43516 9193
rect -44504 9085 -43516 9159
rect -44504 9051 -44414 9085
rect -43630 9051 -43516 9085
rect -46202 7523 -46072 7557
rect -45288 7523 -45214 7557
rect -46202 7449 -45214 7523
rect -46202 7415 -46072 7449
rect -45288 7415 -45214 7449
rect -47808 5887 -47730 5921
rect -46946 5887 -46820 5921
rect -47808 5813 -46820 5887
rect -47808 5779 -47730 5813
rect -46946 5779 -46820 5813
rect -49458 4251 -49388 4285
rect -48604 4251 -48470 4285
rect -49458 4236 -48470 4251
rect -47808 4285 -46820 5779
rect -46202 5921 -45214 7415
rect -44504 7557 -43516 9051
rect -42852 9193 -41864 10687
rect -41202 10831 -40214 12325
rect -39550 12467 -38562 13961
rect -37892 14103 -36904 15597
rect -36244 15739 -35256 17233
rect -34550 17485 -33562 18979
rect -32902 19121 -31914 20615
rect -31254 20649 -30266 20906
rect -31254 20615 -31152 20649
rect -30368 20615 -30266 20649
rect -32902 19087 -32810 19121
rect -32026 19087 -31914 19121
rect -32902 19013 -31914 19087
rect -32902 18979 -32810 19013
rect -32026 18979 -31914 19013
rect -34550 17451 -34468 17485
rect -33684 17451 -33562 17485
rect -34550 17267 -33562 17451
rect -34550 17233 -34466 17267
rect -33682 17233 -33562 17267
rect -36244 15705 -36124 15739
rect -35340 15705 -35256 15739
rect -36244 15631 -35256 15705
rect -36244 15597 -36124 15631
rect -35340 15597 -35256 15631
rect -37892 14069 -37782 14103
rect -36998 14069 -36904 14103
rect -37892 13995 -36904 14069
rect -37892 13961 -37782 13995
rect -36998 13961 -36904 13995
rect -39550 12433 -39440 12467
rect -38656 12433 -38562 12467
rect -39550 12359 -38562 12433
rect -39550 12325 -39440 12359
rect -38656 12325 -38562 12359
rect -41202 10797 -41098 10831
rect -40314 10797 -40214 10831
rect -41202 10721 -40214 10797
rect -41202 10687 -41098 10721
rect -40314 10687 -40214 10721
rect -42852 9159 -42756 9193
rect -41972 9159 -41864 9193
rect -42852 9085 -41864 9159
rect -42852 9051 -42756 9085
rect -41972 9051 -41864 9085
rect -44504 7523 -44414 7557
rect -43630 7523 -43516 7557
rect -44504 7449 -43516 7523
rect -44504 7415 -44414 7449
rect -43630 7415 -43516 7449
rect -46202 5887 -46072 5921
rect -45288 5887 -45214 5921
rect -46202 5813 -45214 5887
rect -46202 5779 -46072 5813
rect -45288 5779 -45214 5813
rect -47808 4251 -47730 4285
rect -46946 4251 -46820 4285
rect -47808 4236 -46820 4251
rect -46202 4285 -45214 5779
rect -44504 5921 -43516 7415
rect -42852 7557 -41864 9051
rect -41202 9193 -40214 10687
rect -39550 10831 -38562 12325
rect -37892 12467 -36904 13961
rect -36244 14103 -35256 15597
rect -34550 15739 -33562 17233
rect -32902 17485 -31914 18979
rect -31254 19121 -30266 20615
rect -29606 20649 -28618 20858
rect -29606 20615 -29494 20649
rect -28710 20615 -28618 20649
rect -31254 19087 -31152 19121
rect -30368 19087 -30266 19121
rect -31254 19013 -30266 19087
rect -31254 18979 -31152 19013
rect -30368 18979 -30266 19013
rect -32902 17451 -32810 17485
rect -32026 17451 -31914 17485
rect -32902 17267 -31914 17451
rect -32902 17233 -32808 17267
rect -32024 17233 -31914 17267
rect -34550 15705 -34466 15739
rect -33682 15705 -33562 15739
rect -34550 15631 -33562 15705
rect -34550 15597 -34466 15631
rect -33682 15597 -33562 15631
rect -36244 14069 -36124 14103
rect -35340 14069 -35256 14103
rect -36244 13995 -35256 14069
rect -36244 13961 -36124 13995
rect -35340 13961 -35256 13995
rect -37892 12433 -37782 12467
rect -36998 12433 -36904 12467
rect -37892 12359 -36904 12433
rect -37892 12325 -37782 12359
rect -36998 12325 -36904 12359
rect -39550 10797 -39440 10831
rect -38656 10797 -38562 10831
rect -39550 10721 -38562 10797
rect -39550 10687 -39440 10721
rect -38656 10687 -38562 10721
rect -41202 9159 -41098 9193
rect -40314 9159 -40214 9193
rect -41202 9085 -40214 9159
rect -41202 9051 -41098 9085
rect -40314 9051 -40214 9085
rect -42852 7523 -42756 7557
rect -41972 7523 -41864 7557
rect -42852 7449 -41864 7523
rect -42852 7415 -42756 7449
rect -41972 7415 -41864 7449
rect -44504 5887 -44414 5921
rect -43630 5887 -43516 5921
rect -44504 5813 -43516 5887
rect -44504 5779 -44414 5813
rect -43630 5779 -43516 5813
rect -46202 4251 -46072 4285
rect -45288 4251 -45214 4285
rect -46202 4236 -45214 4251
rect -44504 4285 -43516 5779
rect -42852 5921 -41864 7415
rect -41202 7557 -40214 9051
rect -39550 9193 -38562 10687
rect -37892 10831 -36904 12325
rect -36244 12467 -35256 13961
rect -34550 14103 -33562 15597
rect -32902 15739 -31914 17233
rect -31254 17485 -30266 18979
rect -29606 19121 -28618 20615
rect -27834 19740 -26806 21200
rect -20956 21298 -20714 22026
rect -19328 21298 -19118 22026
rect -20956 21056 -19118 21298
rect 36822 20988 38660 21256
rect 36822 20260 37064 20988
rect 38450 20260 38660 20988
rect 36822 20018 38660 20260
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -29606 19087 -29494 19121
rect -28710 19087 -28618 19121
rect -29606 19013 -28618 19087
rect -29606 18979 -29494 19013
rect -28710 18979 -28618 19013
rect -31254 17451 -31152 17485
rect -30368 17451 -30266 17485
rect -31254 17267 -30266 17451
rect -31254 17233 -31150 17267
rect -30366 17233 -30266 17267
rect -32902 15705 -32808 15739
rect -32024 15705 -31914 15739
rect -32902 15631 -31914 15705
rect -32902 15597 -32808 15631
rect -32024 15597 -31914 15631
rect -34550 14069 -34466 14103
rect -33682 14069 -33562 14103
rect -34550 13995 -33562 14069
rect -34550 13961 -34466 13995
rect -33682 13961 -33562 13995
rect -36244 12433 -36124 12467
rect -35340 12433 -35256 12467
rect -36244 12359 -35256 12433
rect -36244 12325 -36124 12359
rect -35340 12325 -35256 12359
rect -37892 10797 -37782 10831
rect -36998 10797 -36904 10831
rect -37892 10721 -36904 10797
rect -37892 10687 -37782 10721
rect -36998 10687 -36904 10721
rect -39550 9159 -39440 9193
rect -38656 9159 -38562 9193
rect -39550 9085 -38562 9159
rect -39550 9051 -39440 9085
rect -38656 9051 -38562 9085
rect -41202 7523 -41098 7557
rect -40314 7523 -40214 7557
rect -41202 7449 -40214 7523
rect -41202 7415 -41098 7449
rect -40314 7415 -40214 7449
rect -42852 5887 -42756 5921
rect -41972 5887 -41864 5921
rect -42852 5813 -41864 5887
rect -42852 5779 -42756 5813
rect -41972 5779 -41864 5813
rect -44504 4251 -44414 4285
rect -43630 4251 -43516 4285
rect -44504 4236 -43516 4251
rect -42852 4285 -41864 5779
rect -41202 5921 -40214 7415
rect -39550 7557 -38562 9051
rect -37892 9193 -36904 10687
rect -36244 10831 -35256 12325
rect -34550 12467 -33562 13961
rect -32902 14103 -31914 15597
rect -31254 15739 -30266 17233
rect -29606 17485 -28618 18979
rect -27834 17740 -26806 19274
rect -29606 17451 -29494 17485
rect -28710 17451 -28618 17485
rect -29606 17267 -28618 17451
rect -29606 17233 -29492 17267
rect -28708 17233 -28618 17267
rect -31254 15705 -31150 15739
rect -30366 15705 -30266 15739
rect -31254 15631 -30266 15705
rect -31254 15597 -31150 15631
rect -30366 15597 -30266 15631
rect -32902 14069 -32808 14103
rect -32024 14069 -31914 14103
rect -32902 13995 -31914 14069
rect -32902 13961 -32808 13995
rect -32024 13961 -31914 13995
rect -34550 12433 -34466 12467
rect -33682 12433 -33562 12467
rect -34550 12359 -33562 12433
rect -34550 12325 -34466 12359
rect -33682 12325 -33562 12359
rect -36244 10797 -36124 10831
rect -35340 10797 -35256 10831
rect -36244 10721 -35256 10797
rect -36244 10687 -36124 10721
rect -35340 10687 -35256 10721
rect -37892 9159 -37782 9193
rect -36998 9159 -36904 9193
rect -37892 9085 -36904 9159
rect -37892 9051 -37782 9085
rect -36998 9051 -36904 9085
rect -39550 7523 -39440 7557
rect -38656 7523 -38562 7557
rect -39550 7449 -38562 7523
rect -39550 7415 -39440 7449
rect -38656 7415 -38562 7449
rect -41202 5887 -41098 5921
rect -40314 5887 -40214 5921
rect -41202 5813 -40214 5887
rect -41202 5779 -41098 5813
rect -40314 5779 -40214 5813
rect -42852 4251 -42756 4285
rect -41972 4251 -41864 4285
rect -42852 4236 -41864 4251
rect -41202 4285 -40214 5779
rect -39550 5921 -38562 7415
rect -37892 7557 -36904 9051
rect -36244 9193 -35256 10687
rect -34550 10831 -33562 12325
rect -32902 12467 -31914 13961
rect -31254 14103 -30266 15597
rect -29606 15739 -28618 17233
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -29606 15705 -29492 15739
rect -28708 15705 -28618 15739
rect -29606 15631 -28618 15705
rect -29606 15597 -29492 15631
rect -28708 15597 -28618 15631
rect -31254 14069 -31150 14103
rect -30366 14069 -30266 14103
rect -31254 13995 -30266 14069
rect -31254 13961 -31150 13995
rect -30366 13961 -30266 13995
rect -32902 12433 -32808 12467
rect -32024 12433 -31914 12467
rect -32902 12359 -31914 12433
rect -32902 12325 -32808 12359
rect -32024 12325 -31914 12359
rect -34550 10797 -34466 10831
rect -33682 10797 -33562 10831
rect -34550 10721 -33562 10797
rect -34550 10687 -34466 10721
rect -33682 10687 -33562 10721
rect -36244 9159 -36124 9193
rect -35340 9159 -35256 9193
rect -36244 9085 -35256 9159
rect -36244 9051 -36124 9085
rect -35340 9051 -35256 9085
rect -37892 7523 -37782 7557
rect -36998 7523 -36904 7557
rect -37892 7449 -36904 7523
rect -37892 7415 -37782 7449
rect -36998 7415 -36904 7449
rect -39550 5887 -39440 5921
rect -38656 5887 -38562 5921
rect -39550 5813 -38562 5887
rect -39550 5779 -39440 5813
rect -38656 5779 -38562 5813
rect -41202 4251 -41098 4285
rect -40314 4251 -40214 4285
rect -41202 4236 -40214 4251
rect -39550 4285 -38562 5779
rect -37892 5921 -36904 7415
rect -36244 7557 -35256 9051
rect -34550 9193 -33562 10687
rect -32902 10831 -31914 12325
rect -31254 12467 -30266 13961
rect -29606 14103 -28618 15597
rect -27834 15740 -26806 17274
rect -20956 18026 -19118 18286
rect -20956 17298 -20714 18026
rect -19328 17298 -19118 18026
rect -20956 17056 -19118 17298
rect 36822 16988 38660 17256
rect 36822 16260 37064 16988
rect 38450 16260 38660 16988
rect 36822 16018 38660 16260
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -29606 14069 -29492 14103
rect -28708 14069 -28618 14103
rect -29606 13995 -28618 14069
rect -29606 13961 -29492 13995
rect -28708 13961 -28618 13995
rect -31254 12433 -31150 12467
rect -30366 12433 -30266 12467
rect -31254 12359 -30266 12433
rect -31254 12325 -31150 12359
rect -30366 12325 -30266 12359
rect -32902 10797 -32808 10831
rect -32024 10797 -31914 10831
rect -32902 10721 -31914 10797
rect -32902 10687 -32808 10721
rect -32024 10687 -31914 10721
rect -34550 9159 -34466 9193
rect -33682 9159 -33562 9193
rect -34550 9085 -33562 9159
rect -34550 9051 -34466 9085
rect -33682 9051 -33562 9085
rect -36244 7523 -36124 7557
rect -35340 7523 -35256 7557
rect -36244 7449 -35256 7523
rect -36244 7415 -36124 7449
rect -35340 7415 -35256 7449
rect -37892 5887 -37782 5921
rect -36998 5887 -36904 5921
rect -37892 5813 -36904 5887
rect -37892 5779 -37782 5813
rect -36998 5779 -36904 5813
rect -39550 4251 -39440 4285
rect -38656 4251 -38562 4285
rect -39550 4236 -38562 4251
rect -37892 4285 -36904 5779
rect -36244 5921 -35256 7415
rect -34550 7557 -33562 9051
rect -32902 9193 -31914 10687
rect -31254 10831 -30266 12325
rect -29606 12467 -28618 13961
rect -27834 13740 -26806 15274
rect -18294 14908 -16456 15184
rect -18294 14180 -18052 14908
rect -16666 14180 -16456 14908
rect -18294 13938 -16456 14180
rect -14294 15084 -14106 15180
rect -13566 15084 -12456 15180
rect -14294 14908 -12456 15084
rect -14294 14180 -14052 14908
rect -12666 14180 -12456 14908
rect -14294 13938 -12456 14180
rect -10294 14908 -8456 15180
rect -10294 14180 -10052 14908
rect -8666 14180 -8456 14908
rect -10294 13938 -8456 14180
rect -6294 14908 -4456 15180
rect -6294 14180 -6052 14908
rect -4666 14180 -4456 14908
rect -6294 13938 -4456 14180
rect -2294 14908 -456 15180
rect -2294 14180 -2052 14908
rect -666 14180 -456 14908
rect -2294 13938 -456 14180
rect 1706 14908 3544 15180
rect 1706 14180 1948 14908
rect 3334 14180 3544 14908
rect 1706 13938 3544 14180
rect 5706 14908 7544 15180
rect 5706 14180 5948 14908
rect 7334 14180 7544 14908
rect 5706 13938 7544 14180
rect 9706 14908 11544 15180
rect 9706 14180 9948 14908
rect 11334 14180 11544 14908
rect 9706 13938 11544 14180
rect 13706 14908 15544 15180
rect 13706 14180 13948 14908
rect 15334 14180 15544 14908
rect 13706 13938 15544 14180
rect 17706 14908 19544 15180
rect 17706 14180 17948 14908
rect 19334 14180 19544 14908
rect 17706 13938 19544 14180
rect 21706 14908 23544 15180
rect 21706 14180 21948 14908
rect 23334 14180 23544 14908
rect 21706 13938 23544 14180
rect 25706 14908 27544 15180
rect 25706 14180 25948 14908
rect 27334 14180 27544 14908
rect 25706 13938 27544 14180
rect 29706 14908 31544 15180
rect 29706 14180 29948 14908
rect 31334 14180 31544 14908
rect 29706 13938 31544 14180
rect 33706 14908 35544 15180
rect 33706 14180 33948 14908
rect 35334 14180 35544 14908
rect 33706 13938 35544 14180
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -29606 12433 -29492 12467
rect -28708 12433 -28618 12467
rect -29606 12359 -28618 12433
rect -29606 12325 -29492 12359
rect -28708 12325 -28618 12359
rect -31254 10797 -31150 10831
rect -30366 10797 -30266 10831
rect -31254 10721 -30266 10797
rect -31254 10687 -31150 10721
rect -30366 10687 -30266 10721
rect -32902 9159 -32808 9193
rect -32024 9159 -31914 9193
rect -32902 9085 -31914 9159
rect -32902 9051 -32808 9085
rect -32024 9051 -31914 9085
rect -34550 7523 -34466 7557
rect -33682 7523 -33562 7557
rect -34550 7449 -33562 7523
rect -34550 7415 -34466 7449
rect -33682 7415 -33562 7449
rect -36244 5887 -36124 5921
rect -35340 5887 -35256 5921
rect -36244 5813 -35256 5887
rect -36244 5779 -36124 5813
rect -35340 5779 -35256 5813
rect -37892 4251 -37782 4285
rect -36998 4251 -36904 4285
rect -37892 4236 -36904 4251
rect -36244 4285 -35256 5779
rect -34550 5921 -33562 7415
rect -32902 7557 -31914 9051
rect -31254 9193 -30266 10687
rect -29606 10831 -28618 12325
rect -27834 11740 -26806 13274
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect 17792 12068 19104 12262
rect 17792 11574 18000 12068
rect 18960 11574 19104 12068
rect 17792 11354 19104 11574
rect -29606 10797 -29492 10831
rect -28708 10797 -28618 10831
rect -29606 10721 -28618 10797
rect -29606 10687 -29492 10721
rect -28708 10687 -28618 10721
rect -31254 9159 -31150 9193
rect -30366 9159 -30266 9193
rect -31254 9085 -30266 9159
rect -31254 9051 -31150 9085
rect -30366 9051 -30266 9085
rect -32902 7523 -32808 7557
rect -32024 7523 -31914 7557
rect -32902 7449 -31914 7523
rect -32902 7415 -32808 7449
rect -32024 7415 -31914 7449
rect -34550 5887 -34466 5921
rect -33682 5887 -33562 5921
rect -34550 5813 -33562 5887
rect -34550 5779 -34466 5813
rect -33682 5779 -33562 5813
rect -36244 4251 -36124 4285
rect -35340 4251 -35256 4285
rect -36244 4236 -35256 4251
rect -34550 4285 -33562 5779
rect -32902 5921 -31914 7415
rect -31254 7557 -30266 9051
rect -29606 9193 -28618 10687
rect -27834 9740 -26806 11274
rect 116 10802 560 10812
rect 5346 10802 5790 10812
rect 10576 10802 11020 10812
rect 15806 10802 16250 10812
rect 116 10732 124 10802
rect 556 10732 560 10802
rect 5346 10732 5354 10802
rect 5786 10732 5790 10802
rect 10576 10732 10584 10802
rect 11016 10732 11020 10802
rect 15806 10732 15814 10802
rect 16246 10732 16250 10802
rect 116 10720 560 10732
rect 5346 10720 5790 10732
rect 10576 10720 11020 10732
rect 15806 10720 16250 10732
rect 116 10482 560 10492
rect 5346 10482 5790 10492
rect 10576 10482 11020 10492
rect 15806 10482 16250 10492
rect 116 10412 124 10482
rect 556 10412 560 10482
rect 5346 10412 5354 10482
rect 5786 10412 5790 10482
rect 10576 10412 10584 10482
rect 11016 10412 11020 10482
rect 15806 10412 15814 10482
rect 16246 10412 16250 10482
rect 116 10400 560 10412
rect 5346 10400 5790 10412
rect 10576 10400 11020 10412
rect 15806 10400 16250 10412
rect 116 10162 560 10172
rect 15806 10162 16250 10172
rect 116 10092 124 10162
rect 556 10092 560 10162
rect 116 10080 560 10092
rect 15806 10092 15814 10162
rect 16246 10092 16250 10162
rect 15806 10080 16250 10092
rect 116 9842 560 9852
rect 15806 9842 16250 9852
rect 116 9772 124 9842
rect 556 9772 560 9842
rect 116 9760 560 9772
rect 15806 9772 15814 9842
rect 16246 9772 16250 9842
rect 15806 9760 16250 9772
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect 116 9522 560 9532
rect 15806 9522 16250 9532
rect 116 9452 124 9522
rect 556 9452 560 9522
rect 116 9440 560 9452
rect 15806 9452 15814 9522
rect 16246 9452 16250 9522
rect 15806 9440 16250 9452
rect -29606 9159 -29492 9193
rect -28708 9159 -28618 9193
rect -29606 9085 -28618 9159
rect -29606 9051 -29492 9085
rect -28708 9051 -28618 9085
rect -31254 7523 -31150 7557
rect -30366 7523 -30266 7557
rect -31254 7449 -30266 7523
rect -31254 7415 -31150 7449
rect -30366 7415 -30266 7449
rect -32902 5887 -32808 5921
rect -32024 5887 -31914 5921
rect -32902 5813 -31914 5887
rect -32902 5779 -32808 5813
rect -32024 5779 -31914 5813
rect -34550 4251 -34466 4285
rect -33682 4251 -33562 4285
rect -34550 4236 -33562 4251
rect -32902 4285 -31914 5779
rect -31254 5921 -30266 7415
rect -29606 7557 -28618 9051
rect -27834 7740 -26806 9274
rect 116 9202 560 9212
rect 15806 9202 16250 9212
rect 116 9132 124 9202
rect 556 9132 560 9202
rect 116 9120 560 9132
rect 15806 9132 15814 9202
rect 16246 9132 16250 9202
rect 15806 9120 16250 9132
rect 116 8882 560 8892
rect 15806 8882 16250 8892
rect 116 8812 124 8882
rect 556 8812 560 8882
rect 116 8800 560 8812
rect 15806 8812 15814 8882
rect 16246 8812 16250 8882
rect 15806 8800 16250 8812
rect 116 8562 560 8572
rect 15806 8562 16250 8572
rect 116 8492 124 8562
rect 556 8492 560 8562
rect 116 8480 560 8492
rect 15806 8492 15814 8562
rect 16246 8492 16250 8562
rect 15806 8480 16250 8492
rect 116 8242 560 8252
rect 15806 8242 16250 8252
rect 116 8172 124 8242
rect 556 8172 560 8242
rect 116 8160 560 8172
rect 15806 8172 15814 8242
rect 16246 8172 16250 8242
rect 15806 8160 16250 8172
rect 116 7922 560 7932
rect 15806 7922 16250 7932
rect 116 7852 124 7922
rect 556 7852 560 7922
rect 116 7840 560 7852
rect 15806 7852 15814 7922
rect 16246 7852 16250 7922
rect 15806 7840 16250 7852
rect -29606 7523 -29492 7557
rect -28708 7523 -28618 7557
rect -29606 7449 -28618 7523
rect -29606 7415 -29492 7449
rect -28708 7415 -28618 7449
rect -31254 5887 -31150 5921
rect -30366 5887 -30266 5921
rect -31254 5813 -30266 5887
rect -31254 5779 -31150 5813
rect -30366 5779 -30266 5813
rect -32902 4251 -32808 4285
rect -32024 4251 -31914 4285
rect -32902 4236 -31914 4251
rect -31254 4285 -30266 5779
rect -29606 5921 -28618 7415
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect 116 7602 560 7612
rect 15806 7602 16250 7612
rect 116 7532 124 7602
rect 556 7532 560 7602
rect 116 7520 560 7532
rect 15806 7532 15814 7602
rect 16246 7532 16250 7602
rect 15806 7520 16250 7532
rect -29606 5887 -29492 5921
rect -28708 5887 -28618 5921
rect -29606 5813 -28618 5887
rect -29606 5779 -29492 5813
rect -28708 5779 -28618 5813
rect -31254 4251 -31150 4285
rect -30366 4251 -30266 4285
rect -31254 4236 -30266 4251
rect -29606 4285 -28618 5779
rect -27834 5740 -26806 7274
rect 116 7282 560 7292
rect 116 7212 124 7282
rect 556 7212 560 7282
rect 10576 7280 11020 7290
rect 15806 7282 16250 7292
rect 5380 7250 5824 7260
rect 116 7200 560 7212
rect 5380 7180 5388 7250
rect 5820 7180 5824 7250
rect 10576 7210 10584 7280
rect 11016 7210 11020 7280
rect 15806 7212 15814 7282
rect 16246 7212 16250 7282
rect 10576 7198 11020 7210
rect 15806 7200 16250 7212
rect 5380 7168 5824 7180
rect 116 6962 560 6972
rect 10576 6962 11020 6972
rect 15806 6962 16250 6972
rect 116 6892 124 6962
rect 556 6892 560 6962
rect 5380 6930 5824 6940
rect 116 6880 560 6892
rect 5380 6860 5388 6930
rect 5820 6860 5824 6930
rect 10576 6892 10584 6962
rect 11016 6892 11020 6962
rect 15806 6892 15814 6962
rect 16246 6892 16250 6962
rect 10576 6880 11020 6892
rect 15806 6880 16250 6892
rect 5380 6848 5824 6860
rect 5834 6442 7324 6448
rect 3512 6406 7324 6442
rect 3512 6404 5888 6406
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 3520 6034 3558 6404
rect 5866 6366 5910 6368
rect 4534 6328 5910 6366
rect 10298 6452 10416 6478
rect 7618 6406 7694 6426
rect 4534 6034 4572 6328
rect 1280 5776 1374 6016
rect 1700 5776 1794 6016
rect 3350 6005 3760 6034
rect 2708 5963 2724 5997
rect 2808 5963 2824 5997
rect 3350 5971 3380 6005
rect 3464 5971 3638 6005
rect 3722 5971 3760 6005
rect 4358 6005 4768 6034
rect 3350 5960 3760 5971
rect 4358 5971 4380 6005
rect 4464 5971 4638 6005
rect 4722 5971 4768 6005
rect 5270 5975 5286 6009
rect 5370 5975 5386 6009
rect 4358 5960 4768 5971
rect 3958 5876 4026 5908
rect 1280 5678 1794 5776
rect 3142 5832 3570 5834
rect 3142 5768 3572 5832
rect -29606 4251 -29492 4285
rect -28708 4251 -28618 4285
rect -29606 4236 -28618 4251
rect -60974 4230 -28618 4236
rect -61050 4112 -28618 4230
rect -61046 4102 -28618 4112
rect -29606 4096 -28618 4102
rect -61936 3972 -61790 4086
rect -61934 3932 -61840 3972
rect -61638 3971 -61236 3982
rect -61642 3937 -61626 3971
rect -61592 3937 -61434 3971
rect -61400 3937 -61236 3971
rect -61638 3932 -61236 3937
rect -61934 3918 -61848 3932
rect -96396 3740 -62544 3910
rect -61934 3884 -61904 3918
rect -61870 3884 -61848 3918
rect -61934 3864 -61848 3884
rect -61282 3926 -61236 3932
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -61282 3482 -61234 3926
rect -27834 3846 -26806 5274
rect 2620 5660 2654 5676
rect 926 5188 1154 5200
rect 926 5164 1618 5188
rect 1118 5154 1618 5164
rect 2620 5156 2654 5172
rect 2878 5660 2912 5676
rect 2878 5156 2912 5172
rect 1118 5119 1174 5154
rect 1102 5085 1118 5119
rect 1152 5114 1174 5119
rect 1564 5136 1618 5154
rect 1152 5085 1168 5114
rect 1334 5083 1350 5117
rect 1384 5083 1400 5117
rect 1564 5115 1628 5136
rect 1562 5081 1578 5115
rect 1612 5081 1628 5115
rect 1780 5083 1796 5117
rect 1830 5083 1846 5117
rect 1574 5078 1616 5081
rect 1110 4591 1158 4594
rect 1102 4557 1118 4591
rect 1152 4557 1168 4591
rect 1246 4589 1390 4596
rect 1468 4594 1530 4596
rect 1110 4526 1158 4557
rect 1246 4556 1350 4589
rect 930 4478 1200 4480
rect 1246 4478 1282 4556
rect 1334 4555 1350 4556
rect 1384 4555 1400 4589
rect 1468 4587 1618 4594
rect 1694 4589 1832 4592
rect 930 4472 1282 4478
rect 1468 4553 1578 4587
rect 1612 4553 1628 4587
rect 1694 4555 1796 4589
rect 1830 4555 1846 4589
rect 1694 4554 1832 4555
rect 1468 4544 1618 4553
rect 1468 4530 1530 4544
rect 1468 4474 1506 4530
rect 1694 4474 1730 4554
rect 930 4438 1142 4472
rect 1176 4438 1282 4472
rect 1342 4440 1358 4474
rect 1392 4440 1506 4474
rect 1560 4440 1576 4474
rect 1610 4440 1730 4474
rect 1782 4438 1798 4472
rect 1832 4438 1848 4472
rect 930 4434 1200 4438
rect 3144 4358 3186 5768
rect 3528 5756 3572 5768
rect 3530 5734 3572 5756
rect 3960 5756 4026 5876
rect 3276 5668 3310 5684
rect 3266 5180 3276 5238
rect 3530 5668 3574 5734
rect 3530 5644 3534 5668
rect 3310 5180 3318 5238
rect 3266 5048 3318 5180
rect 3568 5644 3574 5668
rect 3792 5668 3826 5684
rect 3534 5164 3568 5180
rect 3784 5180 3792 5234
rect 3826 5180 3836 5234
rect 3784 5060 3836 5180
rect 3960 5060 4022 5756
rect 4528 5732 4966 5832
rect 4276 5668 4310 5684
rect 3598 5048 4022 5060
rect 3266 5040 4022 5048
rect 4270 5180 4276 5202
rect 4530 5668 4574 5732
rect 4530 5646 4534 5668
rect 4310 5180 4316 5202
rect 4270 5070 4316 5180
rect 4568 5646 4574 5668
rect 4792 5668 4826 5684
rect 4534 5164 4568 5180
rect 4786 5180 4792 5214
rect 4826 5180 4832 5214
rect 4786 5070 4832 5180
rect 4270 5040 4832 5070
rect 3266 4976 4832 5040
rect 3266 4974 3838 4976
rect 3944 4974 4832 4976
rect 3514 4972 3588 4974
rect 3784 4972 3836 4974
rect 4270 4972 4832 4974
rect 4274 4964 4832 4972
rect 4928 4694 4966 5732
rect 5182 5672 5216 5688
rect 5182 5168 5216 5184
rect 5440 5672 5474 5688
rect 5440 5168 5474 5184
rect 4902 4658 4968 4694
rect 3144 4320 3994 4358
rect 1396 4168 1486 4172
rect 1142 4162 1178 4166
rect 1396 4164 1426 4168
rect 1126 4128 1142 4162
rect 1176 4128 1192 4162
rect 1342 4130 1358 4164
rect 1392 4130 1426 4164
rect 1466 4130 1486 4168
rect 1560 4164 1626 4166
rect 1560 4130 1576 4164
rect 1610 4130 1626 4164
rect 1694 4164 1782 4172
rect 1694 4130 1704 4164
rect 1738 4162 1782 4164
rect 1738 4130 1798 4162
rect 1142 4092 1178 4128
rect 1396 4126 1486 4130
rect 1578 4092 1612 4130
rect 1694 4128 1798 4130
rect 1832 4128 1848 4162
rect 1694 4126 1782 4128
rect 1694 4120 1750 4126
rect 1142 4052 1612 4092
rect 3950 4182 3990 4320
rect 3862 4134 3996 4182
rect -60278 3740 -26756 3846
rect -61282 3478 -61232 3482
rect -96396 2966 -62544 3274
rect -61898 3443 -61482 3452
rect -61898 3409 -61722 3443
rect -61688 3409 -61530 3443
rect -61496 3409 -61480 3443
rect -61898 3390 -61482 3409
rect -61898 3016 -61860 3390
rect -61280 3332 -61232 3478
rect -61360 3330 -61232 3332
rect -61694 3318 -61232 3330
rect -61694 3284 -61674 3318
rect -61640 3284 -61482 3318
rect -61448 3284 -61232 3318
rect -61694 3278 -61232 3284
rect -61694 3276 -61354 3278
rect -61280 3276 -61232 3278
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect 3950 3436 3990 4134
rect 4924 3904 4968 4658
rect 5866 4026 5910 6328
rect 7618 6306 7630 6406
rect 7682 6306 7694 6406
rect 7618 6286 7694 6306
rect 7794 6402 7880 6426
rect 7794 6318 7810 6402
rect 7862 6318 7880 6402
rect 7794 6294 7880 6318
rect 8522 6424 8622 6444
rect 8522 6326 8534 6424
rect 8612 6326 8622 6424
rect 8522 6294 8622 6326
rect 10298 6320 10312 6452
rect 10400 6320 10416 6452
rect 10298 6300 10416 6320
rect 6168 6094 6682 6190
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 6168 5756 6682 5854
rect 6128 5206 6350 5214
rect 6128 5178 6804 5206
rect 6304 5172 6804 5178
rect 6304 5137 6360 5172
rect 6288 5103 6304 5137
rect 6338 5132 6360 5137
rect 6750 5154 6804 5172
rect 6338 5103 6354 5132
rect 6520 5101 6536 5135
rect 6570 5101 6586 5135
rect 6750 5133 6814 5154
rect 6748 5099 6764 5133
rect 6798 5099 6814 5133
rect 6966 5101 6982 5135
rect 7016 5101 7032 5135
rect 6760 5096 6802 5099
rect 6296 4609 6344 4612
rect 6288 4575 6304 4609
rect 6338 4575 6354 4609
rect 6432 4607 6576 4614
rect 6654 4612 6716 4614
rect 6296 4544 6344 4575
rect 6432 4574 6536 4607
rect 6432 4498 6468 4574
rect 6520 4573 6536 4574
rect 6570 4573 6586 4607
rect 6654 4605 6804 4612
rect 6880 4607 7018 4610
rect 6138 4490 6468 4498
rect 6654 4571 6764 4605
rect 6798 4571 6814 4605
rect 6880 4573 6982 4607
rect 7016 4573 7032 4607
rect 6880 4572 7018 4573
rect 6654 4562 6804 4571
rect 6654 4548 6716 4562
rect 6654 4492 6692 4548
rect 6880 4492 6916 4572
rect 6138 4456 6328 4490
rect 6362 4456 6468 4490
rect 6528 4458 6544 4492
rect 6578 4458 6692 4492
rect 6746 4458 6762 4492
rect 6796 4458 6916 4492
rect 6968 4456 6984 4490
rect 7018 4456 7034 4490
rect 6138 4452 6440 4456
rect 6582 4186 6672 4190
rect 6328 4180 6364 4184
rect 6582 4182 6612 4186
rect 6312 4146 6328 4180
rect 6362 4146 6378 4180
rect 6528 4148 6544 4182
rect 6578 4148 6612 4182
rect 6652 4148 6672 4186
rect 6746 4182 6812 4184
rect 6746 4148 6762 4182
rect 6796 4148 6812 4182
rect 6880 4182 6968 4190
rect 6880 4148 6890 4182
rect 6924 4180 6968 4182
rect 6924 4148 6984 4180
rect 6328 4110 6364 4146
rect 6582 4144 6672 4148
rect 6764 4110 6798 4148
rect 6880 4146 6984 4148
rect 7018 4146 7034 4180
rect 6880 4144 6968 4146
rect 6880 4138 6936 4144
rect 6328 4070 6798 4110
rect 5866 3956 5910 3958
rect 4876 3856 4974 3904
rect 3948 3388 3992 3436
rect 4924 3418 4968 3856
rect -60278 3224 -26756 3274
rect -61898 3008 -61526 3016
rect -61898 2974 -61770 3008
rect -61736 2974 -61578 3008
rect -61544 2974 -61526 3008
rect -61898 2964 -61526 2974
rect -61896 2878 -61292 2894
rect -61896 2826 -61864 2878
rect -61806 2826 -61464 2878
rect -61406 2826 -61292 2878
rect -61896 2812 -61292 2826
rect 3950 2836 3990 3388
rect 4922 3358 4970 3418
rect 4924 2836 4968 3358
rect 3950 2750 3998 2836
rect 4924 2798 4972 2836
rect 3954 2720 3998 2750
rect 2714 2570 2730 2604
rect 2814 2570 2830 2604
rect 3340 2572 3356 2606
rect 3740 2572 3756 2606
rect 2626 2476 2660 2492
rect 2626 2372 2660 2388
rect 2884 2476 2918 2492
rect 2884 2372 2918 2388
rect 3102 2478 3136 2494
rect 3102 2374 3136 2390
rect 3958 2478 3996 2720
rect 4930 2716 4972 2798
rect 4312 2572 4328 2606
rect 4712 2572 4728 2606
rect 3958 2390 3960 2478
rect 3994 2390 3996 2478
rect 3958 2364 3996 2390
rect 4074 2478 4108 2494
rect 4074 2374 4108 2390
rect 4932 2478 4970 2716
rect 5248 2570 5264 2604
rect 5348 2570 5364 2604
rect 4966 2390 4970 2478
rect 4932 2370 4970 2390
rect 5160 2476 5194 2492
rect 5160 2372 5194 2388
rect 5418 2476 5452 2492
rect 5418 2372 5452 2388
rect 3316 1698 4628 1892
rect 3316 1204 3524 1698
rect 4484 1204 4628 1698
rect 7636 1394 7680 6286
rect 7812 1630 7854 6294
rect 8544 5852 8612 6294
rect 8544 5400 8604 5852
rect 9284 5758 9338 5928
rect 9730 5760 9800 5762
rect 9948 5760 10006 5988
rect 10328 5878 10396 6300
rect 12764 6192 12872 6204
rect 12764 6106 12778 6192
rect 12860 6106 12872 6192
rect 12764 6088 12872 6106
rect 14196 6174 14294 6180
rect 14196 6120 14218 6174
rect 14278 6120 14294 6174
rect 14196 6104 14294 6120
rect 14668 6104 14732 6114
rect 11480 5882 11994 5978
rect 8644 5703 8660 5737
rect 8744 5703 8760 5737
rect 9133 5729 9608 5758
rect 9123 5695 9139 5729
rect 9223 5695 9397 5729
rect 9481 5695 9608 5729
rect 9133 5686 9608 5695
rect 9730 5731 10288 5760
rect 9730 5697 9797 5731
rect 9881 5697 10055 5731
rect 10139 5697 10288 5731
rect 9730 5690 10288 5697
rect 9791 5688 10288 5690
rect 8544 4912 8556 5400
rect 8590 4912 8604 5400
rect 8544 4900 8604 4912
rect 8798 5400 8854 5420
rect 9297 5408 9331 5464
rect 8798 4912 8814 5400
rect 8848 4912 8854 5400
rect 8556 4896 8590 4900
rect 8798 4584 8854 4912
rect 9293 5392 9331 5408
rect 9551 5406 9585 5408
rect 9290 4904 9293 4980
rect 9327 5098 9331 5392
rect 9547 5392 9589 5406
rect 9327 4904 9336 4980
rect 9035 4888 9069 4894
rect 9290 4558 9336 4904
rect 9547 4898 9551 5392
rect 9585 4898 9589 5392
rect 9955 5410 9989 5436
rect 9951 5394 9989 5410
rect 9945 5040 9951 5164
rect 9985 5164 9989 5394
rect 10209 5394 10243 5410
rect 9985 5040 9991 5164
rect 9945 5010 9991 5040
rect 9547 4658 9589 4898
rect 9693 4890 9727 4900
rect 9542 4378 9590 4658
rect 9948 4546 9988 5010
rect 10202 4900 10209 4964
rect 10202 4890 10243 4900
rect 10334 5374 10386 5878
rect 10438 5677 10454 5711
rect 10538 5677 10554 5711
rect 11480 5642 11574 5882
rect 11900 5642 11994 5882
rect 11480 5544 11994 5642
rect 10608 5388 10642 5390
rect 10202 4618 10241 4890
rect 10334 4886 10350 5374
rect 10384 4886 10386 5374
rect 10334 4878 10386 4886
rect 10598 5374 10650 5388
rect 10598 4886 10608 5374
rect 10642 4886 10650 5374
rect 10934 5292 11110 5324
rect 10934 5216 10964 5292
rect 11074 5216 11110 5292
rect 10934 5174 11110 5216
rect 11408 5184 11980 5218
rect 10350 4870 10384 4878
rect 10202 4616 10244 4618
rect 9532 4268 9590 4378
rect 9532 3998 9584 4268
rect 8514 3958 9584 3998
rect 8518 3940 9584 3958
rect 9944 4000 9992 4546
rect 10200 4366 10246 4616
rect 10598 4516 10650 4886
rect 10982 4890 11022 5174
rect 11480 5149 11536 5184
rect 11464 5115 11480 5149
rect 11514 5144 11536 5149
rect 11926 5166 11980 5184
rect 11514 5115 11530 5144
rect 11696 5113 11712 5147
rect 11746 5113 11762 5147
rect 11926 5145 11990 5166
rect 11924 5111 11940 5145
rect 11974 5111 11990 5145
rect 12142 5113 12158 5147
rect 12192 5113 12208 5147
rect 11936 5108 11978 5111
rect 10982 4850 11390 4890
rect 10244 4326 10246 4366
rect 10596 4264 10650 4516
rect 11180 4576 11296 4590
rect 11180 4506 11198 4576
rect 11274 4506 11296 4576
rect 11180 4488 11296 4506
rect 9944 3962 10248 4000
rect 8518 3914 8576 3940
rect 9944 3932 10514 3962
rect 9944 3930 9992 3932
rect 8514 3900 8576 3914
rect 10200 3908 10514 3932
rect 8514 3783 8584 3900
rect 9154 3784 9232 3792
rect 10168 3784 10246 3792
rect 8495 3765 8608 3783
rect 9154 3782 9240 3784
rect 9648 3782 9684 3784
rect 10168 3782 10254 3784
rect 8495 3664 8505 3765
rect 8605 3664 8608 3765
rect 8886 3756 9692 3782
rect 9900 3770 10652 3782
rect 10712 3770 10888 3786
rect 9900 3768 10888 3770
rect 9900 3756 10738 3768
rect 8882 3722 8898 3756
rect 8966 3722 9156 3756
rect 9224 3722 9414 3756
rect 9482 3722 9692 3756
rect 9896 3722 9912 3756
rect 9980 3722 10170 3756
rect 10238 3722 10428 3756
rect 10496 3722 10738 3756
rect 8495 3645 8608 3664
rect 8886 3716 9692 3722
rect 9900 3716 10738 3722
rect 10862 3716 10888 3768
rect 8524 2580 8578 3645
rect 8775 3559 8827 3596
rect 8775 3409 8786 3559
rect 8820 3409 8827 3559
rect 8775 3304 8827 3409
rect 8782 3014 8826 3304
rect 8886 3200 8972 3716
rect 9044 3574 9078 3575
rect 9154 3200 9240 3716
rect 8882 3166 8898 3200
rect 8966 3166 8982 3200
rect 9140 3166 9156 3200
rect 9224 3166 9240 3200
rect 8886 3152 8972 3166
rect 9154 3162 9240 3166
rect 9296 3559 9340 3584
rect 9296 3409 9302 3559
rect 9336 3409 9340 3559
rect 8778 3003 8826 3014
rect 8778 2853 8786 3003
rect 8820 2853 8826 3003
rect 8778 2834 8826 2853
rect 9296 3003 9340 3409
rect 9412 3200 9498 3716
rect 9560 3393 9594 3398
rect 9398 3166 9414 3200
rect 9482 3166 9498 3200
rect 9412 3160 9498 3166
rect 9296 2978 9302 3003
rect 9292 2853 9302 2978
rect 9336 2853 9340 3003
rect 9292 2844 9340 2853
rect 8778 2746 8822 2834
rect 9292 2746 9336 2844
rect 9560 2837 9594 2842
rect 8776 2668 9340 2746
rect 8524 2568 8590 2580
rect 8524 2528 8538 2568
rect 8580 2528 8590 2568
rect 8524 2516 8590 2528
rect 9170 2390 9210 2668
rect 9648 2600 9684 3716
rect 9789 3559 9841 3596
rect 9789 3409 9800 3559
rect 9834 3409 9841 3559
rect 9789 3304 9841 3409
rect 9796 3014 9840 3304
rect 9900 3200 9986 3716
rect 10058 3574 10092 3575
rect 10168 3200 10254 3716
rect 9896 3166 9912 3200
rect 9980 3166 9996 3200
rect 10154 3166 10170 3200
rect 10238 3166 10254 3200
rect 9900 3152 9986 3166
rect 10168 3162 10254 3166
rect 10310 3559 10354 3584
rect 10310 3409 10316 3559
rect 10350 3409 10354 3559
rect 9792 3003 9840 3014
rect 9792 2853 9800 3003
rect 9834 2853 9840 3003
rect 9792 2834 9840 2853
rect 10310 3003 10354 3409
rect 10426 3200 10512 3716
rect 10712 3698 10888 3716
rect 10574 3393 10608 3398
rect 10412 3166 10428 3200
rect 10496 3166 10512 3200
rect 10426 3160 10512 3166
rect 10310 2978 10316 3003
rect 10306 2853 10316 2978
rect 10350 2853 10354 3003
rect 10306 2844 10354 2853
rect 9792 2746 9836 2834
rect 10306 2746 10350 2844
rect 10574 2837 10608 2842
rect 9790 2680 10354 2746
rect 9790 2668 10444 2680
rect 10184 2644 10444 2668
rect 10400 2512 10444 2644
rect 10400 2510 10824 2512
rect 10400 2468 10952 2510
rect 10772 2466 10952 2468
rect 11194 2390 11230 4488
rect 9170 2352 11230 2390
rect 11332 3338 11366 4850
rect 11472 4621 11520 4624
rect 11464 4587 11480 4621
rect 11514 4587 11530 4621
rect 11608 4619 11752 4626
rect 11830 4624 11892 4626
rect 11472 4556 11520 4587
rect 11608 4586 11712 4619
rect 11608 4508 11644 4586
rect 11696 4585 11712 4586
rect 11746 4585 11762 4619
rect 11830 4617 11980 4624
rect 12056 4619 12194 4622
rect 11416 4502 11644 4508
rect 11830 4583 11940 4617
rect 11974 4583 11990 4617
rect 12056 4585 12158 4619
rect 12192 4585 12208 4619
rect 12056 4584 12194 4585
rect 11830 4574 11980 4583
rect 11830 4560 11892 4574
rect 11830 4504 11868 4560
rect 12056 4504 12092 4584
rect 11416 4468 11504 4502
rect 11538 4468 11644 4502
rect 11704 4470 11720 4504
rect 11754 4470 11868 4504
rect 11922 4470 11938 4504
rect 11972 4470 12092 4504
rect 12144 4468 12160 4502
rect 12194 4468 12210 4502
rect 11416 4462 11558 4468
rect 11758 4198 11848 4202
rect 11504 4192 11540 4196
rect 11758 4194 11788 4198
rect 11488 4158 11504 4192
rect 11538 4158 11554 4192
rect 11704 4160 11720 4194
rect 11754 4160 11788 4194
rect 11828 4160 11848 4198
rect 11922 4194 11988 4196
rect 11922 4160 11938 4194
rect 11972 4160 11988 4194
rect 12056 4194 12144 4202
rect 12056 4160 12066 4194
rect 12100 4192 12144 4194
rect 12100 4160 12160 4192
rect 11504 4122 11540 4158
rect 11758 4156 11848 4160
rect 11940 4122 11974 4160
rect 12056 4158 12160 4160
rect 12194 4158 12210 4192
rect 12056 4156 12144 4158
rect 12056 4150 12112 4156
rect 11504 4082 11974 4122
rect 11332 3292 12686 3338
rect 11332 2290 11366 3292
rect 9554 2242 11366 2290
rect 9554 1986 9610 2242
rect 10762 2174 12308 2182
rect 10158 2128 12308 2174
rect 10158 1986 10212 2128
rect 10762 2126 12308 2128
rect 9235 1977 9520 1979
rect 9144 1960 9520 1977
rect 9144 1920 9248 1960
rect 9446 1920 9520 1960
rect 9144 1915 9520 1920
rect 9235 1909 9520 1915
rect 9554 1896 9608 1986
rect 9841 1958 10062 1979
rect 9841 1956 9859 1958
rect 9840 1922 9856 1956
rect 9841 1920 9859 1922
rect 9841 1909 10062 1920
rect 9107 1841 9141 1844
rect 9095 1833 9141 1841
rect 9095 1828 9145 1833
rect 9095 1740 9107 1828
rect 9141 1740 9145 1828
rect 9095 1714 9145 1740
rect 9562 1828 9607 1896
rect 9562 1740 9565 1828
rect 9599 1740 9607 1828
rect 9562 1733 9607 1740
rect 9685 1834 9737 1847
rect 10163 1844 10203 1986
rect 9685 1828 9748 1834
rect 9685 1740 9702 1828
rect 9736 1740 9748 1828
rect 9565 1724 9599 1733
rect 9106 1630 9145 1714
rect 9685 1723 9748 1740
rect 10160 1828 10203 1844
rect 10194 1740 10203 1828
rect 10160 1738 10203 1740
rect 10160 1724 10194 1738
rect 9685 1630 9737 1723
rect 7812 1584 9148 1630
rect 9106 1580 9145 1584
rect 9686 1394 9736 1630
rect 7636 1354 9736 1394
rect 10738 1514 12050 1708
rect 3316 984 4628 1204
rect 10738 1020 10946 1514
rect 11906 1020 12050 1514
rect 10738 800 12050 1020
rect 12800 46 12842 6088
rect 13918 5575 13934 5609
rect 14018 5575 14034 5609
rect 14216 5384 14266 6104
rect 14662 6070 16254 6104
rect 14362 5557 14378 5591
rect 14562 5557 14578 5591
rect 13830 5272 13864 5288
rect 13830 4768 13864 4784
rect 14088 5272 14122 5288
rect 14216 5254 14264 5384
rect 14216 5214 14224 5254
rect 14088 4768 14122 4784
rect 14258 5214 14264 5254
rect 14668 5254 14732 6070
rect 15290 5998 16344 6002
rect 15238 5962 16344 5998
rect 14786 5352 14836 5784
rect 14934 5557 14950 5591
rect 15134 5557 15150 5591
rect 14668 5216 14682 5254
rect 14224 4750 14258 4766
rect 14650 4766 14682 4824
rect 14716 5216 14732 5254
rect 14788 5254 14836 5352
rect 14788 5216 14796 5254
rect 14716 4766 14736 4824
rect 14650 4402 14736 4766
rect 14830 5216 14836 5254
rect 15238 5254 15302 5962
rect 16916 5824 17430 5920
rect 15506 5587 15522 5621
rect 15606 5587 15622 5621
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect 15238 5226 15254 5254
rect 14796 4750 14830 4766
rect 15224 4766 15254 4804
rect 15288 5226 15302 5254
rect 15418 5284 15452 5300
rect 15288 4766 15326 4804
rect 15418 4780 15452 4796
rect 15676 5284 15710 5300
rect 17036 5010 17174 5016
rect 17036 4980 17636 5010
rect 17136 4976 17636 4980
rect 17136 4941 17192 4976
rect 17120 4907 17136 4941
rect 17170 4936 17192 4941
rect 17582 4958 17636 4976
rect 17170 4907 17186 4936
rect 17352 4905 17368 4939
rect 17402 4905 17418 4939
rect 17582 4937 17646 4958
rect 17580 4903 17596 4937
rect 17630 4903 17646 4937
rect 17798 4905 17814 4939
rect 17848 4905 17864 4939
rect 17592 4900 17634 4903
rect 15676 4780 15710 4796
rect 15224 4412 15326 4766
rect 17128 4413 17176 4416
rect 14650 4394 14712 4402
rect 14624 4058 14712 4394
rect 15224 4390 15308 4412
rect 14618 3944 14718 4058
rect 15222 4048 15308 4390
rect 17120 4379 17136 4413
rect 17170 4379 17186 4413
rect 17264 4411 17408 4418
rect 17486 4416 17548 4418
rect 17128 4348 17176 4379
rect 17264 4378 17368 4411
rect 17264 4300 17300 4378
rect 17352 4377 17368 4378
rect 17402 4377 17418 4411
rect 17486 4409 17636 4416
rect 17712 4411 17850 4414
rect 16976 4294 17300 4300
rect 17486 4375 17596 4409
rect 17630 4375 17646 4409
rect 17712 4377 17814 4411
rect 17848 4377 17864 4411
rect 17712 4376 17850 4377
rect 17486 4366 17636 4375
rect 17486 4352 17548 4366
rect 17486 4296 17524 4352
rect 17712 4296 17748 4376
rect 16976 4260 17160 4294
rect 17194 4260 17300 4294
rect 17360 4262 17376 4296
rect 17410 4262 17524 4296
rect 17578 4262 17594 4296
rect 17628 4262 17748 4296
rect 17800 4260 17816 4294
rect 17850 4260 17866 4294
rect 15214 3958 15332 4048
rect 17414 3990 17504 3994
rect 17160 3984 17196 3988
rect 17414 3986 17444 3990
rect 14624 3356 14712 3944
rect 14628 3354 14712 3356
rect 15222 3390 15308 3958
rect 17144 3950 17160 3984
rect 17194 3950 17210 3984
rect 17360 3952 17376 3986
rect 17410 3952 17444 3986
rect 17484 3952 17504 3990
rect 17578 3986 17644 3988
rect 17578 3952 17594 3986
rect 17628 3952 17644 3986
rect 17712 3986 17800 3994
rect 17712 3952 17722 3986
rect 17756 3984 17800 3986
rect 17756 3952 17816 3984
rect 17160 3914 17196 3950
rect 17414 3948 17504 3952
rect 17596 3914 17630 3952
rect 17712 3950 17816 3952
rect 17850 3950 17866 3984
rect 17712 3948 17800 3950
rect 17712 3942 17768 3948
rect 17160 3874 17630 3914
rect 26112 3638 26592 3676
rect 26112 3580 26138 3638
rect 25870 3570 26138 3580
rect 13406 3152 13422 3186
rect 13506 3152 13522 3186
rect 13956 3018 13972 3052
rect 14056 3018 14072 3052
rect 14214 3018 14230 3052
rect 14314 3018 14330 3052
rect 14472 3018 14488 3052
rect 14572 3018 14588 3052
rect 14628 2978 14714 3354
rect 15222 3352 15304 3390
rect 15222 3304 15688 3352
rect 15632 3200 15688 3304
rect 25854 3296 26138 3570
rect 14956 3018 14972 3052
rect 15056 3018 15072 3052
rect 15214 3018 15230 3052
rect 15314 3018 15330 3052
rect 15472 3018 15488 3052
rect 15572 3018 15588 3052
rect 14116 2908 14714 2978
rect 15642 2974 15686 3200
rect 16004 3102 16020 3136
rect 16104 3102 16120 3136
rect 15114 2972 15192 2974
rect 15316 2972 15688 2974
rect 13858 2774 13914 2800
rect 13318 2408 13352 2424
rect 13318 1004 13352 1020
rect 13576 2408 13610 2424
rect 13576 1004 13610 1020
rect 13858 2386 13868 2774
rect 13902 2386 13914 2774
rect 13858 1818 13914 2386
rect 14116 2774 14172 2908
rect 14116 2386 14126 2774
rect 14160 2386 14172 2774
rect 14384 2774 14418 2790
rect 13956 2062 13972 2096
rect 14056 2062 14072 2096
rect 13858 1430 13868 1818
rect 13902 1430 13914 1818
rect 13858 862 13914 1430
rect 14116 1818 14172 2386
rect 14376 2386 14384 2772
rect 14632 2774 14688 2908
rect 15114 2904 15688 2972
rect 14868 2780 14902 2790
rect 15120 2784 15170 2904
rect 15634 2898 15686 2904
rect 15384 2788 15418 2790
rect 14418 2386 14432 2772
rect 14632 2718 14642 2774
rect 14214 2062 14230 2096
rect 14314 2062 14330 2096
rect 14116 1430 14126 1818
rect 14160 1430 14172 1818
rect 13956 1106 13972 1140
rect 14056 1106 14072 1140
rect 13858 500 13868 862
rect 13854 474 13868 500
rect 13902 474 13914 862
rect 13854 468 13914 474
rect 14116 862 14172 1430
rect 14376 1818 14432 2386
rect 14634 2386 14642 2718
rect 14676 2768 14688 2774
rect 14856 2774 14912 2780
rect 14676 2386 14690 2768
rect 14472 2062 14488 2096
rect 14572 2062 14588 2096
rect 14376 1430 14384 1818
rect 14418 1430 14432 1818
rect 14214 1106 14230 1140
rect 14314 1106 14330 1140
rect 14116 474 14126 862
rect 14160 474 14172 862
rect 13854 372 13912 468
rect 14116 436 14172 474
rect 14376 862 14432 1430
rect 14634 1818 14690 2386
rect 14634 1430 14642 1818
rect 14676 1430 14690 1818
rect 14472 1106 14488 1140
rect 14572 1106 14588 1140
rect 14376 474 14384 862
rect 14418 506 14432 862
rect 14634 862 14690 1430
rect 14418 474 14434 506
rect 14376 372 14434 474
rect 14634 474 14642 862
rect 14676 474 14690 862
rect 14634 436 14690 474
rect 14856 2386 14868 2774
rect 14902 2386 14912 2774
rect 14856 1818 14912 2386
rect 15118 2774 15174 2784
rect 15118 2386 15126 2774
rect 15160 2386 15174 2774
rect 14956 2062 14972 2096
rect 15056 2062 15072 2096
rect 14856 1430 14868 1818
rect 14902 1430 14912 1818
rect 14856 862 14912 1430
rect 15118 1818 15174 2386
rect 15370 2774 15426 2788
rect 15634 2784 15684 2898
rect 15370 2386 15384 2774
rect 15418 2386 15426 2774
rect 15214 2062 15230 2096
rect 15314 2062 15330 2096
rect 15118 1430 15126 1818
rect 15160 1430 15174 1818
rect 14956 1106 14972 1140
rect 15056 1106 15072 1140
rect 14856 474 14868 862
rect 14902 496 14912 862
rect 15118 862 15174 1430
rect 15370 1818 15426 2386
rect 15628 2774 15684 2784
rect 15628 2386 15642 2774
rect 15676 2386 15684 2774
rect 15472 2062 15488 2096
rect 15572 2062 15588 2096
rect 15370 1430 15384 1818
rect 15418 1430 15426 1818
rect 15214 1106 15230 1140
rect 15314 1106 15330 1140
rect 14902 474 14916 496
rect 14856 448 14916 474
rect 15118 474 15126 862
rect 15160 474 15174 862
rect 15118 452 15174 474
rect 15370 862 15426 1430
rect 15628 1818 15684 2386
rect 15628 1430 15642 1818
rect 15676 1430 15684 1818
rect 15472 1106 15488 1140
rect 15572 1106 15588 1140
rect 15370 474 15384 862
rect 15418 496 15426 862
rect 15628 862 15684 1430
rect 15916 2358 15950 2374
rect 15916 954 15950 970
rect 16174 2358 16208 2374
rect 17370 1832 18682 2026
rect 17370 1338 17578 1832
rect 18538 1338 18682 1832
rect 17370 1118 18682 1338
rect 25854 1342 26050 3296
rect 26112 3246 26138 3296
rect 26538 3580 26592 3638
rect 26538 3572 26954 3580
rect 32438 3576 32484 3578
rect 32246 3574 32498 3576
rect 31600 3572 32242 3574
rect 26538 3550 32242 3572
rect 26538 3304 26988 3550
rect 27236 3304 27988 3550
rect 28236 3304 28988 3550
rect 29236 3304 29988 3550
rect 30236 3304 30988 3550
rect 31236 3326 32242 3550
rect 32484 3326 32504 3574
rect 31236 3304 32504 3326
rect 26538 3300 32504 3304
rect 26538 3296 26616 3300
rect 31600 3296 32504 3300
rect 26538 3246 26592 3296
rect 31986 3294 32504 3296
rect 26112 3216 26592 3246
rect 26206 3204 26522 3216
rect 32206 3058 32504 3294
rect 32200 3050 32504 3058
rect 32200 2904 32496 3050
rect 30282 2903 30482 2904
rect 28544 2899 28744 2900
rect 27392 2895 27592 2896
rect 26780 2887 26980 2888
rect 26780 2854 26930 2887
rect 26162 2356 26256 2358
rect 26160 2352 26368 2356
rect 26160 2182 26176 2352
rect 26352 2182 26368 2352
rect 26780 2300 26816 2854
rect 26914 2853 26930 2854
rect 26964 2853 26980 2887
rect 27392 2862 27542 2895
rect 27090 2832 27124 2848
rect 26886 2794 26920 2810
rect 26886 2466 26920 2482
rect 26974 2794 27008 2810
rect 27090 2504 27124 2520
rect 27178 2834 27212 2848
rect 27178 2504 27212 2520
rect 26974 2466 27008 2482
rect 27146 2461 27180 2462
rect 27118 2427 27134 2461
rect 27168 2427 27184 2461
rect 26740 2282 26816 2300
rect 27146 2370 27182 2427
rect 27392 2370 27428 2862
rect 27526 2861 27542 2862
rect 27576 2861 27592 2895
rect 27970 2891 28170 2892
rect 27970 2858 28120 2891
rect 27702 2840 27736 2856
rect 27498 2802 27532 2818
rect 27498 2474 27532 2490
rect 27586 2802 27620 2818
rect 27702 2512 27736 2528
rect 27790 2842 27824 2856
rect 27790 2512 27824 2528
rect 27586 2474 27620 2490
rect 27758 2469 27792 2470
rect 27730 2435 27746 2469
rect 27780 2435 27796 2469
rect 27146 2318 27428 2370
rect 26740 2280 27076 2282
rect 26160 1840 26368 2182
rect 26678 2264 27030 2280
rect 26678 2190 26690 2264
rect 26780 2248 27030 2264
rect 26780 2246 26812 2248
rect 27014 2246 27030 2248
rect 27064 2246 27080 2280
rect 26780 2190 26796 2246
rect 26678 2176 26796 2190
rect 26886 2196 26920 2212
rect 26982 2196 27016 2212
rect 26966 2104 26982 2150
rect 26886 2056 26920 2072
rect 27078 2196 27112 2212
rect 27016 2104 27032 2150
rect 26982 2056 27016 2072
rect 27078 2056 27112 2072
rect 26918 1988 26934 2022
rect 26968 1988 26984 2022
rect 26928 1968 26984 1988
rect 27146 1968 27182 2318
rect 27392 2290 27428 2318
rect 27758 2350 27794 2435
rect 27970 2350 28006 2858
rect 28104 2857 28120 2858
rect 28154 2857 28170 2891
rect 28544 2866 28694 2899
rect 28280 2836 28314 2852
rect 28168 2814 28210 2816
rect 28076 2798 28110 2814
rect 28076 2470 28110 2486
rect 28164 2798 28210 2814
rect 28198 2508 28210 2798
rect 28280 2508 28314 2524
rect 28368 2838 28402 2852
rect 28368 2508 28402 2524
rect 28164 2470 28198 2486
rect 28336 2465 28370 2466
rect 28308 2431 28324 2465
rect 28358 2431 28374 2465
rect 27758 2316 28006 2350
rect 27392 2288 27688 2290
rect 27392 2256 27642 2288
rect 27626 2254 27642 2256
rect 27676 2254 27692 2288
rect 27498 2204 27532 2220
rect 27486 2080 27498 2132
rect 27594 2204 27628 2220
rect 27532 2080 27548 2132
rect 27582 2080 27594 2132
rect 27690 2204 27724 2220
rect 27628 2080 27640 2132
rect 27486 2074 27548 2080
rect 27498 2064 27532 2074
rect 27594 2064 27628 2080
rect 27690 2064 27724 2080
rect 27530 1996 27546 2030
rect 27580 1996 27596 2030
rect 26928 1934 27182 1968
rect 27540 1976 27596 1996
rect 27758 1976 27794 2316
rect 27970 2286 28006 2316
rect 28336 2358 28372 2431
rect 28544 2358 28580 2866
rect 28678 2865 28694 2866
rect 28728 2865 28744 2899
rect 29122 2899 29322 2900
rect 29122 2866 29272 2899
rect 28854 2844 28888 2860
rect 28742 2822 28784 2824
rect 28650 2806 28684 2822
rect 28650 2478 28684 2494
rect 28738 2806 28784 2822
rect 28772 2508 28784 2806
rect 28854 2516 28888 2532
rect 28942 2846 28976 2860
rect 28942 2516 28976 2532
rect 28738 2478 28772 2494
rect 28910 2473 28944 2474
rect 28882 2439 28898 2473
rect 28932 2439 28948 2473
rect 28336 2322 28580 2358
rect 27970 2284 28266 2286
rect 27970 2252 28220 2284
rect 28204 2250 28220 2252
rect 28254 2250 28270 2284
rect 28076 2200 28110 2216
rect 28172 2200 28206 2216
rect 28156 2100 28172 2138
rect 28076 2060 28110 2076
rect 28268 2200 28302 2216
rect 28206 2100 28220 2138
rect 28172 2060 28206 2076
rect 28268 2060 28302 2076
rect 28108 1992 28124 2026
rect 28158 1992 28174 2026
rect 27540 1942 27794 1976
rect 28118 1972 28174 1992
rect 28336 1972 28372 2322
rect 28544 2294 28580 2322
rect 28910 2364 28946 2439
rect 29122 2364 29158 2866
rect 29256 2865 29272 2866
rect 29306 2865 29322 2899
rect 29700 2899 29900 2900
rect 29700 2866 29850 2899
rect 29432 2844 29466 2860
rect 29228 2806 29262 2822
rect 29228 2478 29262 2494
rect 29316 2806 29350 2822
rect 29432 2516 29466 2532
rect 29520 2846 29554 2860
rect 29520 2516 29554 2532
rect 29316 2478 29350 2494
rect 29488 2473 29522 2474
rect 29460 2439 29476 2473
rect 29510 2439 29526 2473
rect 28910 2328 29158 2364
rect 28544 2292 28840 2294
rect 28544 2260 28794 2292
rect 28778 2258 28794 2260
rect 28828 2258 28844 2292
rect 28650 2208 28684 2224
rect 28746 2208 28780 2224
rect 28730 2106 28746 2172
rect 28650 2068 28684 2084
rect 28842 2208 28876 2224
rect 28780 2116 28798 2172
rect 28780 2106 28794 2116
rect 28746 2068 28780 2084
rect 28842 2068 28876 2084
rect 28682 2000 28698 2034
rect 28732 2000 28748 2034
rect 28118 1938 28372 1972
rect 28692 1980 28748 2000
rect 28910 1980 28946 2328
rect 29122 2294 29158 2328
rect 29488 2368 29524 2439
rect 29700 2368 29736 2866
rect 29834 2865 29850 2866
rect 29884 2865 29900 2899
rect 30282 2870 30432 2903
rect 30010 2844 30044 2860
rect 29806 2806 29840 2822
rect 29806 2478 29840 2494
rect 29894 2806 29928 2822
rect 30010 2516 30044 2532
rect 30098 2846 30132 2860
rect 30098 2516 30132 2532
rect 29894 2478 29928 2494
rect 30066 2473 30100 2474
rect 30038 2439 30054 2473
rect 30088 2439 30104 2473
rect 29488 2332 29736 2368
rect 29122 2292 29418 2294
rect 29122 2260 29372 2292
rect 29356 2258 29372 2260
rect 29406 2258 29422 2292
rect 29228 2208 29262 2224
rect 29324 2208 29358 2224
rect 29310 2108 29324 2162
rect 29228 2068 29262 2084
rect 29420 2208 29454 2224
rect 29358 2126 29376 2162
rect 29358 2108 29374 2126
rect 29324 2068 29358 2084
rect 29420 2068 29454 2084
rect 29260 2000 29276 2034
rect 29310 2000 29326 2034
rect 28692 1946 28946 1980
rect 29270 1980 29326 2000
rect 29488 1980 29524 2332
rect 29700 2294 29736 2332
rect 30066 2374 30102 2439
rect 30282 2374 30318 2870
rect 30416 2869 30432 2870
rect 30466 2869 30482 2903
rect 30858 2899 31058 2900
rect 30858 2866 31008 2899
rect 30592 2848 30626 2864
rect 30388 2810 30422 2826
rect 30388 2482 30422 2498
rect 30476 2810 30510 2826
rect 30592 2520 30626 2536
rect 30680 2850 30714 2864
rect 30680 2520 30714 2536
rect 30476 2482 30510 2498
rect 30648 2477 30682 2478
rect 30620 2443 30636 2477
rect 30670 2443 30686 2477
rect 30066 2338 30318 2374
rect 29700 2292 29996 2294
rect 29700 2260 29950 2292
rect 29934 2258 29950 2260
rect 29984 2258 30000 2292
rect 29806 2208 29840 2224
rect 29902 2208 29936 2224
rect 29886 2106 29902 2162
rect 29806 2068 29840 2084
rect 29998 2208 30032 2224
rect 29936 2120 29954 2162
rect 29936 2106 29950 2120
rect 29902 2068 29936 2084
rect 29998 2068 30032 2084
rect 29838 2000 29854 2034
rect 29888 2000 29904 2034
rect 29270 1946 29524 1980
rect 29848 1980 29904 2000
rect 30066 1980 30102 2338
rect 30282 2298 30318 2338
rect 30648 2374 30684 2443
rect 30858 2374 30894 2866
rect 30992 2865 31008 2866
rect 31042 2865 31058 2899
rect 31428 2895 31628 2896
rect 31428 2862 31578 2895
rect 31168 2844 31202 2860
rect 30964 2806 30998 2822
rect 30964 2478 30998 2494
rect 31052 2806 31086 2822
rect 31168 2516 31202 2532
rect 31256 2846 31290 2860
rect 31256 2516 31290 2532
rect 31052 2478 31086 2494
rect 31224 2473 31258 2474
rect 31196 2439 31212 2473
rect 31246 2439 31262 2473
rect 30648 2338 30896 2374
rect 31224 2364 31260 2439
rect 31428 2364 31464 2862
rect 31562 2861 31578 2862
rect 31612 2861 31628 2895
rect 31738 2840 31772 2856
rect 31534 2802 31568 2818
rect 31534 2474 31568 2490
rect 31622 2802 31656 2818
rect 31738 2512 31772 2528
rect 31826 2842 31860 2856
rect 32200 2684 32212 2904
rect 32196 2660 32212 2684
rect 32460 2660 32496 2904
rect 32196 2650 32496 2660
rect 32196 2646 32476 2650
rect 31826 2512 31860 2528
rect 31622 2474 31656 2490
rect 31794 2469 31828 2470
rect 31766 2435 31782 2469
rect 31816 2435 31832 2469
rect 30282 2296 30578 2298
rect 30282 2264 30532 2296
rect 30516 2262 30532 2264
rect 30566 2262 30582 2296
rect 30388 2212 30422 2228
rect 30484 2212 30518 2228
rect 30468 2114 30484 2168
rect 30388 2072 30422 2088
rect 30580 2212 30614 2228
rect 30518 2126 30534 2168
rect 30518 2114 30532 2126
rect 30484 2072 30518 2088
rect 30580 2072 30614 2088
rect 30420 2004 30436 2038
rect 30470 2004 30486 2038
rect 29848 1946 30102 1980
rect 30430 1984 30486 2004
rect 30648 1984 30684 2338
rect 30858 2294 30894 2338
rect 31224 2328 31464 2364
rect 30858 2292 31154 2294
rect 30858 2260 31108 2292
rect 31092 2258 31108 2260
rect 31142 2258 31158 2292
rect 30964 2208 30998 2224
rect 31060 2208 31094 2224
rect 31044 2106 31060 2158
rect 30964 2068 30998 2084
rect 31156 2208 31190 2224
rect 31094 2106 31108 2158
rect 31060 2068 31094 2084
rect 31156 2068 31190 2084
rect 30996 2000 31012 2034
rect 31046 2000 31062 2034
rect 30430 1950 30684 1984
rect 31006 1980 31062 2000
rect 31224 1980 31260 2328
rect 31428 2290 31464 2328
rect 31428 2288 31724 2290
rect 31428 2256 31678 2288
rect 31662 2254 31678 2256
rect 31712 2254 31728 2288
rect 31534 2204 31568 2220
rect 31306 2074 31396 2090
rect 31306 2012 31320 2074
rect 31382 2030 31396 2074
rect 31630 2204 31664 2220
rect 31616 2108 31630 2160
rect 31534 2064 31568 2080
rect 31726 2204 31760 2220
rect 31664 2108 31680 2160
rect 31630 2064 31664 2080
rect 31726 2064 31760 2080
rect 31382 2012 31582 2030
rect 31306 1998 31582 2012
rect 31006 1946 31260 1980
rect 31322 1996 31582 1998
rect 31616 1996 31634 2030
rect 31322 1978 31634 1996
rect 31576 1976 31634 1978
rect 31794 1976 31830 2435
rect 32096 2344 32164 2346
rect 32096 2340 32208 2344
rect 32096 2170 32120 2340
rect 32204 2214 32220 2340
rect 32204 2170 32222 2214
rect 32096 2132 32222 2170
rect 31576 1942 31830 1976
rect 32026 2106 32222 2132
rect 32364 2206 32976 2274
rect 32364 2106 32424 2206
rect 32026 1918 32424 2106
rect 30402 1840 30828 1844
rect 32026 1840 32220 1918
rect 26160 1670 26168 1840
rect 26344 1670 26628 1840
rect 26804 1670 27228 1840
rect 27404 1670 27828 1840
rect 28004 1670 28428 1840
rect 28604 1670 29028 1840
rect 29204 1670 29628 1840
rect 29804 1670 30228 1840
rect 30404 1670 30828 1840
rect 31004 1670 31428 1840
rect 31604 1670 32028 1840
rect 32204 1670 32220 1840
rect 32364 1746 32424 1918
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 26160 1668 32030 1670
rect 26160 1666 31620 1668
rect 26160 1658 28472 1666
rect 28936 1658 30122 1666
rect 26160 1656 26940 1658
rect 26160 1654 26570 1656
rect 25854 1068 26044 1342
rect 28162 1136 28856 1140
rect 27910 1130 28856 1136
rect 27910 1128 28422 1130
rect 27910 1086 27926 1128
rect 25854 1062 27218 1068
rect 27880 1066 27926 1086
rect 27692 1062 27926 1066
rect 25854 976 27926 1062
rect 16174 954 16208 970
rect 25856 930 27926 976
rect 28126 930 28182 1128
rect 25856 928 28182 930
rect 28382 930 28422 1128
rect 28622 1128 28856 1130
rect 28622 930 28656 1128
rect 28382 928 28656 930
rect 28830 928 28856 1128
rect 29926 1042 30122 1658
rect 28942 1032 30122 1042
rect 28942 1014 30132 1032
rect 28942 1012 29330 1014
rect 28942 1010 29106 1012
rect 25856 916 28856 928
rect 25856 914 28830 916
rect 25856 912 28402 914
rect 25856 910 28148 912
rect 25856 876 28144 910
rect 15418 474 15432 496
rect 15370 456 15432 474
rect 14858 372 14916 448
rect 15374 372 15432 456
rect 15628 474 15642 862
rect 15676 474 15684 862
rect 27896 856 28144 876
rect 27896 844 27926 856
rect 15628 452 15684 474
rect 27912 656 27926 844
rect 28126 844 28144 856
rect 28938 860 28942 944
rect 29030 862 29106 1010
rect 29256 864 29330 1012
rect 29480 864 29546 1014
rect 29696 1012 29946 1014
rect 29696 864 29738 1012
rect 29256 862 29738 864
rect 29888 864 29946 1012
rect 30096 864 30132 1014
rect 29888 862 30132 864
rect 29030 860 30132 862
rect 28126 710 28142 844
rect 28306 840 28364 848
rect 28306 833 28384 840
rect 28306 799 28324 833
rect 28358 799 28384 833
rect 28938 838 30132 860
rect 28306 798 28384 799
rect 28710 831 28760 832
rect 28306 790 28364 798
rect 28710 797 28726 831
rect 28760 797 28776 831
rect 28480 778 28514 794
rect 28280 740 28314 756
rect 28126 656 28280 710
rect 27912 642 28280 656
rect 27912 622 28142 642
rect 13850 264 15432 372
rect 27912 422 27926 622
rect 28126 422 28142 622
rect 27912 382 28142 422
rect 28368 740 28402 756
rect 28314 642 28320 710
rect 28280 412 28314 428
rect 28480 450 28514 466
rect 28568 778 28602 794
rect 28710 790 28760 797
rect 28568 450 28602 466
rect 28682 738 28716 754
rect 28368 412 28402 428
rect 28682 410 28716 426
rect 28770 738 28804 754
rect 28938 502 28986 838
rect 28770 410 28804 426
rect 14728 46 14768 264
rect 12800 2 14768 46
rect 27912 182 27926 382
rect 28126 182 28142 382
rect 28508 373 28524 407
rect 28558 406 28574 407
rect 28558 373 28580 406
rect 28514 364 28580 373
rect 28940 358 28986 502
rect 29938 790 30132 838
rect 29938 640 29956 790
rect 30106 640 30132 790
rect 29938 598 30132 640
rect 29062 442 29150 452
rect 29062 408 29088 442
rect 29122 408 29150 442
rect 29250 442 29338 452
rect 29250 408 29280 442
rect 29314 408 29338 442
rect 29442 442 29530 454
rect 29442 408 29472 442
rect 29506 408 29530 442
rect 29632 442 29720 454
rect 29632 408 29664 442
rect 29698 408 29720 442
rect 29938 448 29962 598
rect 30112 448 30132 598
rect 29938 404 30132 448
rect 28940 342 28944 358
rect 28308 327 28374 328
rect 28712 327 28778 328
rect 28308 293 28324 327
rect 28358 293 28374 327
rect 28708 293 28724 327
rect 28758 293 28778 327
rect 28308 286 28374 293
rect 28480 272 28514 288
rect 27912 144 28142 182
rect 12800 0 14766 2
rect 27912 -48 27924 144
rect 28124 -48 28142 144
rect 27912 -88 28142 -48
rect 27912 -288 27926 -88
rect 28126 -288 28142 -88
rect 28280 234 28314 250
rect 28280 -94 28314 -78
rect 28368 234 28402 250
rect 28480 -56 28514 -40
rect 28568 272 28602 288
rect 28712 286 28778 293
rect 28942 288 28944 342
rect 28568 -56 28602 -40
rect 28680 234 28714 250
rect 28368 -94 28402 -78
rect 28680 -94 28714 -78
rect 28768 234 28802 250
rect 28930 136 28944 288
rect 28934 -72 28944 136
rect 28768 -94 28802 -78
rect 28510 -99 28576 -98
rect 28508 -133 28524 -99
rect 28558 -133 28576 -99
rect 28510 -140 28576 -133
rect 28708 -181 28774 -176
rect 28308 -182 28324 -181
rect 28216 -215 28324 -182
rect 28358 -182 28374 -181
rect 28358 -215 28376 -182
rect 28216 -218 28376 -215
rect 28708 -215 28724 -181
rect 28758 -215 28774 -181
rect 28708 -218 28774 -215
rect 28480 -236 28514 -220
rect 27912 -324 28142 -288
rect 27912 -458 27924 -324
rect 27906 -524 27924 -458
rect 28124 -458 28142 -324
rect 28280 -274 28314 -258
rect 28124 -524 28148 -458
rect 27906 -714 28148 -524
rect 28280 -602 28314 -586
rect 28368 -274 28402 -258
rect 28480 -564 28514 -548
rect 28568 -236 28602 -220
rect 28568 -564 28602 -548
rect 28680 -274 28714 -258
rect 28368 -602 28402 -586
rect 28680 -602 28714 -586
rect 28768 -274 28802 -258
rect 28978 288 28986 358
rect 29040 358 29074 374
rect 28978 -72 28990 288
rect 29028 102 29040 278
rect 29034 -8 29040 102
rect 28944 -282 28978 -266
rect 29136 358 29170 374
rect 29074 -8 29082 184
rect 29126 102 29136 278
rect 29132 -6 29136 102
rect 29040 -282 29074 -266
rect 29232 358 29266 374
rect 29170 -6 29180 186
rect 29222 -66 29232 290
rect 29136 -282 29170 -266
rect 29328 358 29362 374
rect 29266 -66 29278 144
rect 29318 132 29328 296
rect 29316 -78 29328 132
rect 29232 -282 29266 -266
rect 29424 358 29458 374
rect 29362 -78 29372 132
rect 29412 -72 29424 284
rect 29328 -282 29362 -266
rect 29520 358 29554 374
rect 29512 138 29520 286
rect 29458 -72 29468 138
rect 29508 -72 29520 138
rect 29424 -282 29458 -266
rect 29616 358 29650 374
rect 29554 138 29556 286
rect 29554 -72 29564 138
rect 29610 134 29616 280
rect 29604 -76 29616 134
rect 29520 -282 29554 -266
rect 29712 358 29746 374
rect 29650 134 29654 280
rect 29702 144 29712 264
rect 29650 -76 29660 134
rect 29698 -66 29712 144
rect 29616 -282 29650 -266
rect 29808 358 29842 374
rect 29746 -66 29754 144
rect 29712 -282 29746 -266
rect 29938 254 29966 404
rect 30116 254 30132 404
rect 29938 218 30132 254
rect 29938 68 29968 218
rect 30118 68 30132 218
rect 29938 52 30132 68
rect 29936 32 30132 52
rect 29936 -26 29974 32
rect 29808 -282 29842 -266
rect 29938 -118 29974 -26
rect 30124 -118 30132 32
rect 29938 -176 30132 -118
rect 28976 -318 28992 -316
rect 28974 -350 28992 -318
rect 29026 -318 29042 -316
rect 29026 -350 29060 -318
rect 28974 -364 29060 -350
rect 29152 -350 29184 -316
rect 29218 -350 29240 -316
rect 29360 -318 29376 -316
rect 29152 -362 29240 -350
rect 29348 -350 29376 -318
rect 29410 -318 29426 -316
rect 29410 -350 29436 -318
rect 29348 -364 29436 -350
rect 29540 -350 29568 -316
rect 29602 -350 29628 -316
rect 29540 -362 29628 -350
rect 29728 -350 29760 -316
rect 29794 -350 29816 -316
rect 29938 -326 29970 -176
rect 30120 -326 30132 -176
rect 29938 -336 30132 -326
rect 29728 -362 29816 -350
rect 29936 -412 30132 -336
rect 29936 -466 29964 -412
rect 28768 -602 28802 -586
rect 28894 -488 29964 -466
rect 28508 -607 28578 -606
rect 28508 -641 28524 -607
rect 28558 -641 28578 -607
rect 28508 -654 28578 -641
rect 28894 -636 28912 -488
rect 29062 -490 29964 -488
rect 29062 -636 29124 -490
rect 28894 -640 29124 -636
rect 29274 -496 29964 -490
rect 29274 -640 29332 -496
rect 28894 -646 29332 -640
rect 29482 -498 29964 -496
rect 29482 -500 29752 -498
rect 29482 -646 29540 -500
rect 28894 -650 29540 -646
rect 29690 -648 29752 -500
rect 29902 -562 29964 -498
rect 30114 -562 30132 -412
rect 29902 -648 30132 -562
rect 29690 -650 30132 -648
rect 28894 -670 30132 -650
rect 28894 -672 28968 -670
rect 30064 -672 30132 -670
rect 27906 -722 28328 -714
rect 27906 -736 28800 -722
rect 27906 -746 28042 -736
rect 8734 -934 10850 -922
rect 8734 -992 8763 -934
rect 8797 -992 8855 -934
rect 8889 -992 8947 -934
rect 8981 -992 9039 -934
rect 9073 -992 9131 -934
rect 9165 -992 9223 -934
rect 9257 -992 9315 -934
rect 9349 -992 9407 -934
rect 9441 -992 9499 -934
rect 9533 -992 9591 -934
rect 9625 -992 9683 -934
rect 9717 -992 9775 -934
rect 9809 -992 9867 -934
rect 9901 -992 9959 -934
rect 9993 -992 10051 -934
rect 10085 -992 10143 -934
rect 10177 -992 10235 -934
rect 10269 -992 10327 -934
rect 10361 -992 10419 -934
rect 10453 -992 10511 -934
rect 10545 -992 10603 -934
rect 10637 -992 10695 -934
rect 10729 -992 10787 -934
rect 10821 -992 10850 -934
rect 11200 -934 13316 -920
rect 11200 -992 11229 -934
rect 11263 -992 11321 -934
rect 11355 -992 11413 -934
rect 11447 -992 11505 -934
rect 11539 -992 11597 -934
rect 11631 -992 11689 -934
rect 11723 -992 11781 -934
rect 11815 -992 11873 -934
rect 11907 -992 11965 -934
rect 11999 -992 12057 -934
rect 12091 -992 12149 -934
rect 12183 -992 12241 -934
rect 12275 -992 12333 -934
rect 12367 -992 12425 -934
rect 12459 -992 12517 -934
rect 12551 -992 12609 -934
rect 12643 -992 12701 -934
rect 12735 -992 12793 -934
rect 12827 -992 12885 -934
rect 12919 -992 12977 -934
rect 13011 -992 13069 -934
rect 13103 -992 13161 -934
rect 13195 -992 13253 -934
rect 13287 -992 13316 -934
rect 27912 -936 28042 -746
rect 28242 -738 28800 -736
rect 28242 -936 28348 -738
rect 27912 -938 28348 -936
rect 28548 -938 28628 -738
rect 28790 -938 28800 -738
rect 27912 -952 28800 -938
rect 28032 -954 28800 -952
rect 8752 -1042 8803 -1026
rect 8752 -1076 8769 -1042
rect 8752 -1110 8803 -1076
rect 8837 -1058 8903 -992
rect 8837 -1092 8853 -1058
rect 8887 -1092 8903 -1058
rect 8937 -1042 8971 -1026
rect 8752 -1144 8769 -1110
rect 8937 -1110 8971 -1076
rect 8803 -1144 8902 -1126
rect 8752 -1160 8902 -1144
rect 8752 -1270 8822 -1194
rect 8752 -1304 8766 -1270
rect 8800 -1304 8822 -1270
rect 8752 -1324 8822 -1304
rect 8856 -1255 8902 -1160
rect 8856 -1264 8868 -1255
rect 8890 -1298 8902 -1289
rect 8856 -1358 8902 -1298
rect 8752 -1392 8902 -1358
rect 8752 -1400 8803 -1392
rect 8752 -1434 8769 -1400
rect 8937 -1400 8971 -1162
rect 9005 -1186 9070 -1029
rect 9104 -1034 9154 -992
rect 9104 -1068 9120 -1034
rect 9104 -1084 9154 -1068
rect 9188 -1042 9238 -1026
rect 9188 -1076 9204 -1042
rect 9188 -1092 9238 -1076
rect 9281 -1036 9417 -1026
rect 9281 -1070 9297 -1036
rect 9331 -1070 9417 -1036
rect 9532 -1044 9598 -992
rect 9725 -1034 9799 -992
rect 9281 -1092 9417 -1070
rect 9188 -1118 9222 -1092
rect 9143 -1152 9222 -1118
rect 9256 -1128 9349 -1126
rect 9017 -1196 9109 -1186
rect 9017 -1230 9039 -1196
rect 9073 -1209 9109 -1196
rect 9073 -1230 9075 -1209
rect 9017 -1243 9075 -1230
rect 9017 -1396 9109 -1243
rect 8752 -1450 8803 -1434
rect 8837 -1460 8853 -1426
rect 8887 -1460 8903 -1426
rect 9143 -1424 9177 -1152
rect 9256 -1154 9315 -1128
rect 9290 -1162 9315 -1154
rect 9290 -1188 9349 -1162
rect 9256 -1204 9349 -1188
rect 9211 -1264 9281 -1242
rect 9211 -1298 9223 -1264
rect 9257 -1298 9281 -1264
rect 9211 -1316 9281 -1298
rect 9211 -1350 9234 -1316
rect 9268 -1350 9281 -1316
rect 9211 -1366 9281 -1350
rect 9315 -1322 9349 -1204
rect 9383 -1248 9417 -1092
rect 9451 -1060 9485 -1044
rect 9532 -1078 9548 -1044
rect 9582 -1078 9598 -1044
rect 9632 -1060 9666 -1044
rect 9451 -1112 9485 -1094
rect 9725 -1068 9745 -1034
rect 9779 -1068 9799 -1034
rect 9725 -1084 9799 -1068
rect 9833 -1042 9867 -1026
rect 9632 -1112 9666 -1094
rect 9451 -1146 9666 -1112
rect 9833 -1118 9867 -1076
rect 9914 -1035 10088 -1026
rect 9914 -1069 9930 -1035
rect 9964 -1069 10088 -1035
rect 9914 -1094 10088 -1069
rect 10122 -1034 10172 -992
rect 10156 -1068 10172 -1034
rect 10276 -1034 10420 -992
rect 10122 -1084 10172 -1068
rect 10206 -1060 10240 -1044
rect 9755 -1152 9867 -1118
rect 9755 -1180 9789 -1152
rect 9489 -1214 9505 -1180
rect 9539 -1214 9789 -1180
rect 9928 -1162 9939 -1128
rect 9973 -1154 10020 -1128
rect 9928 -1186 9970 -1162
rect 9383 -1268 9721 -1248
rect 9383 -1282 9687 -1268
rect 9315 -1356 9336 -1322
rect 9370 -1356 9386 -1322
rect 9315 -1366 9386 -1356
rect 9420 -1424 9454 -1282
rect 9495 -1332 9591 -1316
rect 9529 -1366 9567 -1332
rect 9625 -1350 9653 -1316
rect 9687 -1318 9721 -1302
rect 9601 -1366 9653 -1350
rect 9755 -1352 9789 -1214
rect 8937 -1450 8971 -1434
rect 8837 -1502 8903 -1460
rect 9043 -1464 9059 -1430
rect 9093 -1464 9109 -1430
rect 9143 -1458 9192 -1424
rect 9226 -1458 9242 -1424
rect 9283 -1458 9299 -1424
rect 9333 -1458 9454 -1424
rect 9629 -1426 9695 -1410
rect 9043 -1502 9109 -1464
rect 9629 -1460 9645 -1426
rect 9679 -1460 9695 -1426
rect 9629 -1502 9695 -1460
rect 9737 -1430 9789 -1352
rect 9827 -1188 9970 -1186
rect 10004 -1188 10020 -1154
rect 10054 -1170 10088 -1094
rect 10276 -1068 10292 -1034
rect 10326 -1068 10370 -1034
rect 10404 -1068 10420 -1034
rect 10454 -1042 10535 -1026
rect 10686 -1034 10720 -992
rect 10206 -1102 10240 -1094
rect 10488 -1076 10535 -1042
rect 10206 -1136 10366 -1102
rect 9827 -1220 9962 -1188
rect 10054 -1204 10248 -1170
rect 10282 -1204 10298 -1170
rect 9827 -1328 9869 -1220
rect 10054 -1222 10088 -1204
rect 9827 -1362 9835 -1328
rect 9827 -1378 9869 -1362
rect 9903 -1264 9973 -1254
rect 9903 -1280 9939 -1264
rect 9903 -1314 9931 -1280
rect 9965 -1314 9973 -1298
rect 9903 -1378 9973 -1314
rect 10007 -1256 10088 -1222
rect 10007 -1412 10041 -1256
rect 10155 -1269 10263 -1238
rect 10332 -1254 10366 -1136
rect 10454 -1110 10535 -1076
rect 10488 -1144 10535 -1110
rect 10454 -1178 10535 -1144
rect 10488 -1212 10535 -1178
rect 10454 -1228 10535 -1212
rect 10332 -1260 10421 -1254
rect 10189 -1278 10263 -1269
rect 10075 -1306 10119 -1290
rect 10109 -1340 10119 -1306
rect 10155 -1312 10171 -1303
rect 10205 -1312 10263 -1278
rect 10075 -1346 10119 -1340
rect 10215 -1332 10263 -1312
rect 10075 -1380 10181 -1346
rect 9851 -1426 10041 -1412
rect 9737 -1464 9757 -1430
rect 9791 -1464 9807 -1430
rect 9851 -1460 9867 -1426
rect 9901 -1460 10041 -1426
rect 9851 -1468 10041 -1460
rect 10075 -1430 10113 -1414
rect 10075 -1464 10079 -1430
rect 10147 -1426 10181 -1380
rect 10249 -1366 10263 -1332
rect 10215 -1392 10263 -1366
rect 10297 -1270 10421 -1260
rect 10297 -1304 10371 -1270
rect 10405 -1304 10421 -1270
rect 10297 -1320 10421 -1304
rect 10469 -1266 10535 -1228
rect 10469 -1301 10488 -1266
rect 10522 -1301 10535 -1266
rect 10297 -1355 10362 -1320
rect 10469 -1354 10535 -1301
rect 10297 -1410 10361 -1355
rect 10147 -1444 10297 -1426
rect 10331 -1444 10361 -1410
rect 10147 -1460 10361 -1444
rect 10401 -1387 10435 -1365
rect 10075 -1502 10113 -1464
rect 10401 -1502 10435 -1421
rect 10469 -1388 10485 -1354
rect 10519 -1388 10535 -1354
rect 10469 -1422 10535 -1388
rect 10469 -1456 10485 -1422
rect 10519 -1456 10535 -1422
rect 10573 -1068 10589 -1034
rect 10623 -1068 10639 -1034
rect 10573 -1102 10639 -1068
rect 10573 -1136 10589 -1102
rect 10623 -1136 10639 -1102
rect 10573 -1254 10639 -1136
rect 11218 -1042 11269 -1026
rect 10686 -1102 10720 -1068
rect 10686 -1170 10720 -1136
rect 10686 -1220 10720 -1204
rect 10770 -1070 10821 -1054
rect 10804 -1104 10821 -1070
rect 10770 -1138 10821 -1104
rect 10804 -1172 10821 -1138
rect 11218 -1076 11235 -1042
rect 11218 -1110 11269 -1076
rect 11303 -1058 11369 -992
rect 11303 -1092 11319 -1058
rect 11353 -1092 11369 -1058
rect 11403 -1042 11437 -1026
rect 11218 -1144 11235 -1110
rect 11403 -1110 11437 -1076
rect 11269 -1144 11368 -1126
rect 11218 -1160 11368 -1144
rect 10770 -1230 10821 -1172
rect 10573 -1270 10745 -1254
rect 10573 -1304 10711 -1270
rect 10573 -1320 10745 -1304
rect 10779 -1265 10821 -1230
rect 10779 -1299 10783 -1265
rect 10817 -1299 10821 -1265
rect 10573 -1400 10623 -1320
rect 10779 -1360 10821 -1299
rect 11218 -1264 11288 -1194
rect 11218 -1298 11230 -1264
rect 11264 -1270 11288 -1264
rect 11218 -1304 11232 -1298
rect 11266 -1304 11288 -1270
rect 11218 -1324 11288 -1304
rect 11322 -1255 11368 -1160
rect 11322 -1264 11334 -1255
rect 11356 -1298 11368 -1289
rect 11322 -1358 11368 -1298
rect 10770 -1376 10821 -1360
rect 10573 -1434 10589 -1400
rect 10573 -1450 10623 -1434
rect 10686 -1406 10720 -1383
rect 10469 -1464 10535 -1456
rect 10686 -1502 10720 -1440
rect 10804 -1410 10821 -1376
rect 10770 -1466 10821 -1410
rect 11218 -1392 11368 -1358
rect 11218 -1400 11269 -1392
rect 11218 -1434 11235 -1400
rect 11403 -1400 11437 -1162
rect 11471 -1186 11536 -1029
rect 11570 -1034 11620 -992
rect 11570 -1068 11586 -1034
rect 11570 -1084 11620 -1068
rect 11654 -1042 11704 -1026
rect 11654 -1076 11670 -1042
rect 11654 -1092 11704 -1076
rect 11747 -1036 11883 -1026
rect 11747 -1070 11763 -1036
rect 11797 -1070 11883 -1036
rect 11998 -1044 12064 -992
rect 12191 -1034 12265 -992
rect 11747 -1092 11883 -1070
rect 11654 -1118 11688 -1092
rect 11609 -1152 11688 -1118
rect 11722 -1128 11815 -1126
rect 11483 -1196 11575 -1186
rect 11483 -1230 11505 -1196
rect 11539 -1209 11575 -1196
rect 11539 -1230 11541 -1209
rect 11483 -1243 11541 -1230
rect 11483 -1396 11575 -1243
rect 11218 -1450 11269 -1434
rect 11303 -1460 11319 -1426
rect 11353 -1460 11369 -1426
rect 11609 -1424 11643 -1152
rect 11722 -1154 11781 -1128
rect 11756 -1162 11781 -1154
rect 11756 -1188 11815 -1162
rect 11722 -1204 11815 -1188
rect 11677 -1264 11747 -1242
rect 11677 -1298 11689 -1264
rect 11723 -1298 11747 -1264
rect 11677 -1316 11747 -1298
rect 11677 -1350 11700 -1316
rect 11734 -1350 11747 -1316
rect 11677 -1366 11747 -1350
rect 11781 -1322 11815 -1204
rect 11849 -1248 11883 -1092
rect 11917 -1060 11951 -1044
rect 11998 -1078 12014 -1044
rect 12048 -1078 12064 -1044
rect 12098 -1060 12132 -1044
rect 11917 -1112 11951 -1094
rect 12191 -1068 12211 -1034
rect 12245 -1068 12265 -1034
rect 12191 -1084 12265 -1068
rect 12299 -1042 12333 -1026
rect 12098 -1112 12132 -1094
rect 11917 -1146 12132 -1112
rect 12299 -1118 12333 -1076
rect 12380 -1035 12554 -1026
rect 12380 -1069 12396 -1035
rect 12430 -1069 12554 -1035
rect 12380 -1094 12554 -1069
rect 12588 -1034 12638 -992
rect 12622 -1068 12638 -1034
rect 12742 -1034 12886 -992
rect 12588 -1084 12638 -1068
rect 12672 -1060 12706 -1044
rect 12221 -1152 12333 -1118
rect 12221 -1180 12255 -1152
rect 11955 -1214 11971 -1180
rect 12005 -1214 12255 -1180
rect 12394 -1162 12405 -1128
rect 12439 -1154 12486 -1128
rect 12394 -1186 12436 -1162
rect 11849 -1268 12187 -1248
rect 11849 -1282 12153 -1268
rect 11781 -1356 11802 -1322
rect 11836 -1356 11852 -1322
rect 11781 -1366 11852 -1356
rect 11886 -1424 11920 -1282
rect 11961 -1332 12057 -1316
rect 11995 -1366 12033 -1332
rect 12091 -1350 12119 -1316
rect 12153 -1318 12187 -1302
rect 12067 -1366 12119 -1350
rect 12221 -1352 12255 -1214
rect 11403 -1450 11437 -1434
rect 11303 -1502 11369 -1460
rect 11509 -1464 11525 -1430
rect 11559 -1464 11575 -1430
rect 11609 -1458 11658 -1424
rect 11692 -1458 11708 -1424
rect 11749 -1458 11765 -1424
rect 11799 -1458 11920 -1424
rect 12095 -1426 12161 -1410
rect 11509 -1502 11575 -1464
rect 12095 -1460 12111 -1426
rect 12145 -1460 12161 -1426
rect 12095 -1502 12161 -1460
rect 12203 -1430 12255 -1352
rect 12293 -1188 12436 -1186
rect 12470 -1188 12486 -1154
rect 12520 -1170 12554 -1094
rect 12742 -1068 12758 -1034
rect 12792 -1068 12836 -1034
rect 12870 -1068 12886 -1034
rect 12920 -1042 13001 -1026
rect 13152 -1034 13186 -992
rect 12672 -1102 12706 -1094
rect 12954 -1076 13001 -1042
rect 12672 -1136 12832 -1102
rect 12293 -1220 12428 -1188
rect 12520 -1204 12714 -1170
rect 12748 -1204 12764 -1170
rect 12293 -1328 12335 -1220
rect 12520 -1222 12554 -1204
rect 12293 -1362 12301 -1328
rect 12293 -1378 12335 -1362
rect 12369 -1264 12439 -1254
rect 12369 -1280 12405 -1264
rect 12369 -1314 12397 -1280
rect 12431 -1314 12439 -1298
rect 12369 -1378 12439 -1314
rect 12473 -1256 12554 -1222
rect 12473 -1412 12507 -1256
rect 12621 -1269 12729 -1238
rect 12798 -1254 12832 -1136
rect 12920 -1110 13001 -1076
rect 12954 -1144 13001 -1110
rect 12920 -1178 13001 -1144
rect 12954 -1212 13001 -1178
rect 12920 -1228 13001 -1212
rect 12798 -1260 12887 -1254
rect 12655 -1278 12729 -1269
rect 12541 -1306 12585 -1290
rect 12575 -1340 12585 -1306
rect 12621 -1312 12637 -1303
rect 12671 -1312 12729 -1278
rect 12541 -1346 12585 -1340
rect 12681 -1332 12729 -1312
rect 12541 -1380 12647 -1346
rect 12317 -1426 12507 -1412
rect 12203 -1464 12223 -1430
rect 12257 -1464 12273 -1430
rect 12317 -1460 12333 -1426
rect 12367 -1460 12507 -1426
rect 12317 -1468 12507 -1460
rect 12541 -1430 12579 -1414
rect 12541 -1464 12545 -1430
rect 12613 -1426 12647 -1380
rect 12715 -1366 12729 -1332
rect 12681 -1392 12729 -1366
rect 12763 -1270 12887 -1260
rect 12763 -1304 12837 -1270
rect 12871 -1304 12887 -1270
rect 12763 -1320 12887 -1304
rect 12763 -1355 12828 -1320
rect 12935 -1354 13001 -1228
rect 12763 -1410 12827 -1355
rect 12613 -1444 12763 -1426
rect 12797 -1444 12827 -1410
rect 12613 -1460 12827 -1444
rect 12867 -1387 12901 -1365
rect 12541 -1502 12579 -1464
rect 12867 -1502 12901 -1421
rect 12935 -1388 12951 -1354
rect 12985 -1388 13001 -1354
rect 12935 -1422 13001 -1388
rect 12935 -1456 12951 -1422
rect 12985 -1456 13001 -1422
rect 13039 -1068 13055 -1034
rect 13089 -1068 13105 -1034
rect 13039 -1102 13105 -1068
rect 13039 -1136 13055 -1102
rect 13089 -1136 13105 -1102
rect 13039 -1254 13105 -1136
rect 13152 -1102 13186 -1068
rect 13152 -1170 13186 -1136
rect 13152 -1220 13186 -1204
rect 13236 -1070 13287 -1054
rect 13270 -1104 13287 -1070
rect 13236 -1138 13287 -1104
rect 13270 -1172 13287 -1138
rect 13236 -1230 13287 -1172
rect 13039 -1270 13211 -1254
rect 13039 -1304 13177 -1270
rect 13039 -1320 13211 -1304
rect 13245 -1264 13287 -1230
rect 13245 -1298 13251 -1264
rect 13285 -1298 13287 -1264
rect 13039 -1400 13089 -1320
rect 13245 -1360 13287 -1298
rect 13236 -1376 13287 -1360
rect 13039 -1434 13055 -1400
rect 13039 -1450 13089 -1434
rect 13152 -1406 13186 -1383
rect 12935 -1464 13001 -1456
rect 13152 -1502 13186 -1440
rect 13270 -1410 13287 -1376
rect 13236 -1466 13287 -1410
rect 8734 -1564 8763 -1502
rect 8797 -1564 8855 -1502
rect 8889 -1564 8947 -1502
rect 8981 -1564 9039 -1502
rect 9073 -1564 9131 -1502
rect 9165 -1564 9223 -1502
rect 9257 -1564 9315 -1502
rect 9349 -1564 9407 -1502
rect 9441 -1564 9499 -1502
rect 9533 -1564 9591 -1502
rect 9625 -1564 9683 -1502
rect 9717 -1564 9775 -1502
rect 9809 -1564 9867 -1502
rect 9901 -1564 9959 -1502
rect 9993 -1564 10051 -1502
rect 10085 -1564 10143 -1502
rect 10177 -1564 10235 -1502
rect 10269 -1564 10327 -1502
rect 10361 -1564 10419 -1502
rect 10453 -1564 10511 -1502
rect 10545 -1564 10603 -1502
rect 10637 -1564 10695 -1502
rect 10729 -1564 10787 -1502
rect 10821 -1564 10850 -1502
rect 8734 -1607 10850 -1564
rect 11200 -1563 11229 -1502
rect 11263 -1563 11321 -1502
rect 11355 -1563 11413 -1502
rect 11447 -1563 11505 -1502
rect 11539 -1563 11597 -1502
rect 11631 -1563 11689 -1502
rect 11723 -1563 11781 -1502
rect 11815 -1563 11873 -1502
rect 11907 -1563 11965 -1502
rect 11999 -1563 12057 -1502
rect 12091 -1563 12149 -1502
rect 12183 -1563 12241 -1502
rect 12275 -1563 12333 -1502
rect 12367 -1563 12425 -1502
rect 12459 -1563 12517 -1502
rect 12551 -1563 12609 -1502
rect 12643 -1563 12701 -1502
rect 12735 -1563 12793 -1502
rect 12827 -1563 12885 -1502
rect 12919 -1563 12977 -1502
rect 13011 -1563 13069 -1502
rect 13103 -1563 13161 -1502
rect 13195 -1563 13253 -1502
rect 13287 -1563 13316 -1502
rect 11200 -1566 13316 -1563
rect 10152 -1736 10428 -1732
rect 10152 -1794 10181 -1736
rect 10215 -1794 10273 -1736
rect 10307 -1794 10365 -1736
rect 10399 -1794 10428 -1736
rect 11200 -1794 11229 -1735
rect 11263 -1794 11321 -1735
rect 11355 -1794 11413 -1735
rect 11447 -1794 11505 -1735
rect 11539 -1794 11597 -1735
rect 11631 -1794 11689 -1735
rect 11723 -1794 11781 -1735
rect 11815 -1794 11873 -1735
rect 11907 -1794 11965 -1735
rect 11999 -1794 12057 -1735
rect 12091 -1794 12149 -1735
rect 12183 -1794 12241 -1735
rect 12275 -1794 12333 -1735
rect 12367 -1794 12425 -1735
rect 12459 -1794 12517 -1735
rect 12551 -1794 12609 -1735
rect 12643 -1794 12701 -1735
rect 12735 -1794 12793 -1735
rect 12827 -1794 12885 -1735
rect 12919 -1794 12977 -1735
rect 13011 -1794 13069 -1735
rect 13103 -1794 13161 -1735
rect 13195 -1794 13253 -1735
rect 13287 -1794 13316 -1735
rect 10177 -1836 10223 -1794
rect 10177 -1870 10189 -1836
rect 10177 -1904 10223 -1870
rect 10177 -1938 10189 -1904
rect 10177 -1972 10223 -1938
rect 10177 -2006 10189 -1972
rect 10177 -2022 10223 -2006
rect 10257 -1836 10323 -1828
rect 10257 -1870 10273 -1836
rect 10307 -1870 10323 -1836
rect 10257 -1904 10323 -1870
rect 10257 -1938 10273 -1904
rect 10307 -1938 10323 -1904
rect 10257 -1972 10323 -1938
rect 10257 -2006 10273 -1972
rect 10307 -2006 10323 -1972
rect 10257 -2024 10323 -2006
rect 10357 -1836 10399 -1794
rect 10391 -1870 10399 -1836
rect 10357 -1904 10399 -1870
rect 10391 -1938 10399 -1904
rect 10357 -1972 10399 -1938
rect 11218 -1844 11269 -1828
rect 11218 -1878 11235 -1844
rect 11218 -1912 11269 -1878
rect 11303 -1860 11369 -1794
rect 11303 -1894 11319 -1860
rect 11353 -1894 11369 -1860
rect 11403 -1844 11437 -1828
rect 11218 -1946 11235 -1912
rect 11403 -1912 11437 -1878
rect 11269 -1946 11368 -1928
rect 11218 -1962 11368 -1946
rect 10391 -2006 10399 -1972
rect 10357 -2022 10399 -2006
rect 10173 -2066 10239 -2056
rect 10173 -2100 10181 -2066
rect 10215 -2072 10239 -2066
rect 10173 -2106 10189 -2100
rect 10223 -2106 10239 -2072
rect 10273 -2096 10323 -2024
rect 10307 -2130 10323 -2096
rect 11218 -2032 11288 -1996
rect 11218 -2066 11230 -2032
rect 11265 -2066 11288 -2032
rect 11218 -2072 11288 -2066
rect 11218 -2106 11232 -2072
rect 11266 -2106 11288 -2072
rect 11218 -2126 11288 -2106
rect 11322 -2057 11368 -1962
rect 11322 -2066 11334 -2057
rect 11356 -2100 11368 -2091
rect 10177 -2156 10223 -2140
rect 10273 -2144 10323 -2130
rect 10177 -2190 10189 -2156
rect 10177 -2228 10223 -2190
rect 10177 -2262 10189 -2228
rect 10177 -2304 10223 -2262
rect 10257 -2156 10323 -2144
rect 10257 -2190 10273 -2156
rect 10307 -2190 10323 -2156
rect 10257 -2228 10323 -2190
rect 10257 -2262 10273 -2228
rect 10307 -2262 10323 -2228
rect 10257 -2270 10323 -2262
rect 10357 -2156 10399 -2140
rect 10391 -2190 10399 -2156
rect 11322 -2160 11368 -2100
rect 10357 -2228 10399 -2190
rect 10391 -2262 10399 -2228
rect 11218 -2194 11368 -2160
rect 11218 -2202 11269 -2194
rect 11218 -2236 11235 -2202
rect 11403 -2202 11437 -1964
rect 11471 -1988 11536 -1831
rect 11570 -1836 11620 -1794
rect 11570 -1870 11586 -1836
rect 11570 -1886 11620 -1870
rect 11654 -1844 11704 -1828
rect 11654 -1878 11670 -1844
rect 11654 -1894 11704 -1878
rect 11747 -1838 11883 -1828
rect 11747 -1872 11763 -1838
rect 11797 -1872 11883 -1838
rect 11998 -1846 12064 -1794
rect 12191 -1836 12265 -1794
rect 11747 -1894 11883 -1872
rect 11654 -1920 11688 -1894
rect 11609 -1954 11688 -1920
rect 11722 -1930 11815 -1928
rect 11483 -2011 11575 -1988
rect 11483 -2028 11541 -2011
rect 11483 -2062 11505 -2028
rect 11539 -2045 11541 -2028
rect 11539 -2062 11575 -2045
rect 11483 -2198 11575 -2062
rect 11218 -2252 11269 -2236
rect 10357 -2304 10399 -2262
rect 11303 -2262 11319 -2228
rect 11353 -2262 11369 -2228
rect 11609 -2226 11643 -1954
rect 11722 -1956 11781 -1930
rect 11756 -1964 11781 -1956
rect 11756 -1990 11815 -1964
rect 11722 -2006 11815 -1990
rect 11677 -2066 11747 -2044
rect 11677 -2100 11689 -2066
rect 11723 -2100 11747 -2066
rect 11677 -2118 11747 -2100
rect 11677 -2152 11700 -2118
rect 11734 -2152 11747 -2118
rect 11677 -2168 11747 -2152
rect 11781 -2124 11815 -2006
rect 11849 -2050 11883 -1894
rect 11917 -1862 11951 -1846
rect 11998 -1880 12014 -1846
rect 12048 -1880 12064 -1846
rect 12098 -1862 12132 -1846
rect 11917 -1914 11951 -1896
rect 12191 -1870 12211 -1836
rect 12245 -1870 12265 -1836
rect 12191 -1886 12265 -1870
rect 12299 -1844 12333 -1828
rect 12098 -1914 12132 -1896
rect 11917 -1948 12132 -1914
rect 12299 -1920 12333 -1878
rect 12380 -1837 12554 -1828
rect 12380 -1871 12396 -1837
rect 12430 -1871 12554 -1837
rect 12380 -1896 12554 -1871
rect 12588 -1836 12638 -1794
rect 12622 -1870 12638 -1836
rect 12742 -1836 12886 -1794
rect 12588 -1886 12638 -1870
rect 12672 -1862 12706 -1846
rect 12221 -1954 12333 -1920
rect 12221 -1982 12255 -1954
rect 11955 -2016 11971 -1982
rect 12005 -2016 12255 -1982
rect 12394 -1964 12405 -1930
rect 12439 -1956 12486 -1930
rect 12394 -1988 12436 -1964
rect 11849 -2070 12187 -2050
rect 11849 -2084 12153 -2070
rect 11781 -2158 11802 -2124
rect 11836 -2158 11852 -2124
rect 11781 -2168 11852 -2158
rect 11886 -2226 11920 -2084
rect 11961 -2134 12057 -2118
rect 11995 -2168 12033 -2134
rect 12091 -2152 12119 -2118
rect 12153 -2120 12187 -2104
rect 12067 -2168 12119 -2152
rect 12221 -2154 12255 -2016
rect 11403 -2252 11437 -2236
rect 11303 -2304 11369 -2262
rect 11509 -2266 11525 -2232
rect 11559 -2266 11575 -2232
rect 11609 -2260 11658 -2226
rect 11692 -2260 11708 -2226
rect 11749 -2260 11765 -2226
rect 11799 -2260 11920 -2226
rect 12095 -2228 12161 -2212
rect 11509 -2304 11575 -2266
rect 12095 -2262 12111 -2228
rect 12145 -2262 12161 -2228
rect 12095 -2304 12161 -2262
rect 12203 -2232 12255 -2154
rect 12293 -1990 12436 -1988
rect 12470 -1990 12486 -1956
rect 12520 -1972 12554 -1896
rect 12742 -1870 12758 -1836
rect 12792 -1870 12836 -1836
rect 12870 -1870 12886 -1836
rect 12920 -1844 13001 -1828
rect 13152 -1836 13186 -1794
rect 12672 -1904 12706 -1896
rect 12954 -1878 13001 -1844
rect 12672 -1938 12832 -1904
rect 12293 -2022 12428 -1990
rect 12520 -2006 12714 -1972
rect 12748 -2006 12764 -1972
rect 12293 -2130 12335 -2022
rect 12520 -2024 12554 -2006
rect 12293 -2164 12301 -2130
rect 12293 -2180 12335 -2164
rect 12369 -2066 12439 -2056
rect 12369 -2082 12405 -2066
rect 12369 -2116 12397 -2082
rect 12431 -2116 12439 -2100
rect 12369 -2180 12439 -2116
rect 12473 -2058 12554 -2024
rect 12473 -2214 12507 -2058
rect 12621 -2071 12729 -2040
rect 12798 -2056 12832 -1938
rect 12920 -1912 13001 -1878
rect 12954 -1946 13001 -1912
rect 12920 -1980 13001 -1946
rect 12954 -2014 13001 -1980
rect 12920 -2030 13001 -2014
rect 12798 -2062 12887 -2056
rect 12655 -2080 12729 -2071
rect 12541 -2108 12585 -2092
rect 12575 -2142 12585 -2108
rect 12621 -2114 12637 -2105
rect 12671 -2114 12729 -2080
rect 12541 -2148 12585 -2142
rect 12681 -2134 12729 -2114
rect 12541 -2182 12647 -2148
rect 12317 -2228 12507 -2214
rect 12203 -2266 12223 -2232
rect 12257 -2266 12273 -2232
rect 12317 -2262 12333 -2228
rect 12367 -2262 12507 -2228
rect 12317 -2270 12507 -2262
rect 12541 -2232 12579 -2216
rect 12541 -2266 12545 -2232
rect 12613 -2228 12647 -2182
rect 12715 -2168 12729 -2134
rect 12681 -2194 12729 -2168
rect 12763 -2072 12887 -2062
rect 12763 -2106 12837 -2072
rect 12871 -2106 12887 -2072
rect 12763 -2122 12887 -2106
rect 12763 -2157 12828 -2122
rect 12935 -2156 13001 -2030
rect 12763 -2212 12827 -2157
rect 12613 -2246 12763 -2228
rect 12797 -2246 12827 -2212
rect 12613 -2262 12827 -2246
rect 12867 -2189 12901 -2167
rect 12541 -2304 12579 -2266
rect 12867 -2304 12901 -2223
rect 12935 -2190 12951 -2156
rect 12985 -2190 13001 -2156
rect 12935 -2224 13001 -2190
rect 12935 -2258 12951 -2224
rect 12985 -2258 13001 -2224
rect 13039 -1870 13055 -1836
rect 13089 -1870 13105 -1836
rect 13039 -1904 13105 -1870
rect 13039 -1938 13055 -1904
rect 13089 -1938 13105 -1904
rect 13039 -2056 13105 -1938
rect 13152 -1904 13186 -1870
rect 13152 -1972 13186 -1938
rect 13152 -2022 13186 -2006
rect 13236 -1872 13287 -1856
rect 13270 -1906 13287 -1872
rect 13236 -1940 13287 -1906
rect 13270 -1974 13287 -1940
rect 13236 -2032 13287 -1974
rect 13039 -2072 13211 -2056
rect 13039 -2106 13177 -2072
rect 13039 -2122 13211 -2106
rect 13245 -2097 13287 -2032
rect 13039 -2202 13089 -2122
rect 13245 -2131 13249 -2097
rect 13283 -2131 13287 -2097
rect 13245 -2162 13287 -2131
rect 13236 -2178 13287 -2162
rect 13039 -2236 13055 -2202
rect 13039 -2252 13089 -2236
rect 13152 -2208 13186 -2185
rect 12935 -2266 13001 -2258
rect 13152 -2304 13186 -2242
rect 13270 -2212 13287 -2178
rect 13236 -2268 13287 -2212
rect 10152 -2364 10181 -2304
rect 10215 -2364 10273 -2304
rect 10307 -2364 10365 -2304
rect 10399 -2364 10428 -2304
rect 10152 -2366 10428 -2364
rect 11200 -2366 11229 -2304
rect 11263 -2366 11321 -2304
rect 11355 -2366 11413 -2304
rect 11447 -2366 11505 -2304
rect 11539 -2366 11597 -2304
rect 11631 -2366 11689 -2304
rect 11723 -2366 11781 -2304
rect 11815 -2366 11873 -2304
rect 11907 -2366 11965 -2304
rect 11999 -2366 12057 -2304
rect 12091 -2366 12149 -2304
rect 12183 -2366 12241 -2304
rect 12275 -2366 12333 -2304
rect 12367 -2366 12425 -2304
rect 12459 -2366 12517 -2304
rect 12551 -2366 12609 -2304
rect 12643 -2366 12701 -2304
rect 12735 -2366 12793 -2304
rect 12827 -2366 12885 -2304
rect 12919 -2366 12977 -2304
rect 13011 -2366 13069 -2304
rect 13103 -2366 13161 -2304
rect 13195 -2366 13253 -2304
rect 13287 -2366 13316 -2304
rect 11200 -2367 13316 -2366
rect -9158 -4204 33162 -4188
rect -9158 -4262 -9129 -4204
rect -9095 -4262 -9037 -4204
rect -9003 -4262 -8945 -4204
rect -8911 -4262 -8853 -4204
rect -8819 -4262 -8761 -4204
rect -8727 -4262 -8669 -4204
rect -8635 -4262 -8577 -4204
rect -8543 -4262 -8485 -4204
rect -8451 -4262 -8393 -4204
rect -8359 -4262 -8301 -4204
rect -8267 -4262 -8209 -4204
rect -8175 -4262 -8117 -4204
rect -8083 -4262 -8025 -4204
rect -7991 -4262 -7933 -4204
rect -7899 -4262 -7841 -4204
rect -7807 -4262 -7749 -4204
rect -7715 -4262 -7657 -4204
rect -7623 -4262 -7565 -4204
rect -7531 -4262 -7473 -4204
rect -7439 -4262 -7381 -4204
rect -7347 -4262 -7289 -4204
rect -7255 -4262 -7197 -4204
rect -7163 -4262 -7105 -4204
rect -7071 -4262 -7013 -4204
rect -6979 -4262 -6921 -4204
rect -6887 -4262 -6829 -4204
rect -6795 -4262 -6737 -4204
rect -6703 -4262 -6645 -4204
rect -6611 -4262 -6553 -4204
rect -6519 -4262 -6461 -4204
rect -6427 -4262 -6369 -4204
rect -6335 -4262 -6277 -4204
rect -6243 -4262 -6185 -4204
rect -6151 -4262 -6093 -4204
rect -6059 -4262 -6001 -4204
rect -5967 -4262 -5909 -4204
rect -5875 -4262 -5817 -4204
rect -5783 -4262 -5725 -4204
rect -5691 -4262 -5633 -4204
rect -5599 -4262 -5541 -4204
rect -5507 -4262 -5449 -4204
rect -5415 -4262 -5357 -4204
rect -5323 -4262 -5265 -4204
rect -5231 -4262 -5173 -4204
rect -5139 -4262 -5081 -4204
rect -5047 -4262 -4989 -4204
rect -4955 -4262 -4897 -4204
rect -4863 -4262 -4805 -4204
rect -4771 -4262 -4713 -4204
rect -4679 -4262 -4621 -4204
rect -4587 -4262 -4529 -4204
rect -4495 -4262 -4437 -4204
rect -4403 -4262 -4345 -4204
rect -4311 -4262 -4253 -4204
rect -4219 -4262 -4161 -4204
rect -4127 -4262 -4069 -4204
rect -4035 -4262 -3977 -4204
rect -3943 -4262 -3885 -4204
rect -3851 -4262 -3793 -4204
rect -3759 -4262 -3701 -4204
rect -3667 -4262 -3609 -4204
rect -3575 -4262 -3517 -4204
rect -3483 -4262 -3425 -4204
rect -3391 -4262 -3333 -4204
rect -3299 -4262 -3241 -4204
rect -3207 -4262 -3149 -4204
rect -3115 -4262 -3057 -4204
rect -3023 -4262 -2965 -4204
rect -2931 -4262 -2873 -4204
rect -2839 -4262 -2781 -4204
rect -2747 -4262 -2689 -4204
rect -2655 -4262 -2597 -4204
rect -2563 -4262 -2505 -4204
rect -2471 -4262 -2413 -4204
rect -2379 -4262 -2321 -4204
rect -2287 -4262 -2229 -4204
rect -2195 -4262 -2137 -4204
rect -2103 -4262 -2045 -4204
rect -2011 -4262 -1953 -4204
rect -1919 -4262 -1861 -4204
rect -1827 -4262 -1769 -4204
rect -1735 -4262 -1677 -4204
rect -1643 -4262 -1585 -4204
rect -1551 -4262 -1493 -4204
rect -1459 -4262 -1401 -4204
rect -1367 -4262 -1309 -4204
rect -1275 -4262 -1217 -4204
rect -1183 -4262 -1125 -4204
rect -1091 -4262 -1033 -4204
rect -999 -4262 -941 -4204
rect -907 -4262 -849 -4204
rect -815 -4262 -757 -4204
rect -723 -4262 -665 -4204
rect -631 -4262 -573 -4204
rect -539 -4262 -481 -4204
rect -447 -4262 -389 -4204
rect -355 -4262 -297 -4204
rect -263 -4262 -205 -4204
rect -171 -4262 -113 -4204
rect -79 -4262 -21 -4204
rect 13 -4262 71 -4204
rect 105 -4262 163 -4204
rect 197 -4262 255 -4204
rect 289 -4262 347 -4204
rect 381 -4262 439 -4204
rect 473 -4262 531 -4204
rect 565 -4262 623 -4204
rect 657 -4262 715 -4204
rect 749 -4262 807 -4204
rect 841 -4262 899 -4204
rect 933 -4262 991 -4204
rect 1025 -4262 1083 -4204
rect 1117 -4262 1175 -4204
rect 1209 -4262 1267 -4204
rect 1301 -4262 1359 -4204
rect 1393 -4262 1451 -4204
rect 1485 -4262 1543 -4204
rect 1577 -4262 1635 -4204
rect 1669 -4262 1727 -4204
rect 1761 -4262 1819 -4204
rect 1853 -4262 1911 -4204
rect 1945 -4262 2003 -4204
rect 2037 -4262 2095 -4204
rect 2129 -4262 2187 -4204
rect 2221 -4262 2279 -4204
rect 2313 -4262 2371 -4204
rect 2405 -4262 2463 -4204
rect 2497 -4262 2555 -4204
rect 2589 -4262 2647 -4204
rect 2681 -4262 2739 -4204
rect 2773 -4262 2831 -4204
rect 2865 -4262 2923 -4204
rect 2957 -4262 3015 -4204
rect 3049 -4262 3107 -4204
rect 3141 -4262 3199 -4204
rect 3233 -4262 3291 -4204
rect 3325 -4262 3383 -4204
rect 3417 -4262 3475 -4204
rect 3509 -4262 3567 -4204
rect 3601 -4262 3659 -4204
rect 3693 -4262 3751 -4204
rect 3785 -4262 3843 -4204
rect 3877 -4262 3935 -4204
rect 3969 -4262 4027 -4204
rect 4061 -4262 4119 -4204
rect 4153 -4262 4211 -4204
rect 4245 -4262 4303 -4204
rect 4337 -4262 4395 -4204
rect 4429 -4262 4487 -4204
rect 4521 -4262 4579 -4204
rect 4613 -4262 4671 -4204
rect 4705 -4262 4763 -4204
rect 4797 -4262 4855 -4204
rect 4889 -4262 4947 -4204
rect 4981 -4262 5039 -4204
rect 5073 -4262 5131 -4204
rect 5165 -4262 5223 -4204
rect 5257 -4262 5315 -4204
rect 5349 -4262 5407 -4204
rect 5441 -4262 5499 -4204
rect 5533 -4262 5591 -4204
rect 5625 -4262 5683 -4204
rect 5717 -4262 5775 -4204
rect 5809 -4262 5867 -4204
rect 5901 -4262 5959 -4204
rect 5993 -4262 6051 -4204
rect 6085 -4262 6143 -4204
rect 6177 -4262 6235 -4204
rect 6269 -4262 6327 -4204
rect 6361 -4262 6419 -4204
rect 6453 -4262 6511 -4204
rect 6545 -4262 6603 -4204
rect 6637 -4262 6695 -4204
rect 6729 -4262 6787 -4204
rect 6821 -4262 6879 -4204
rect 6913 -4262 6971 -4204
rect 7005 -4262 7063 -4204
rect 7097 -4262 7155 -4204
rect 7189 -4262 7247 -4204
rect 7281 -4262 7339 -4204
rect 7373 -4262 7431 -4204
rect 7465 -4262 7523 -4204
rect 7557 -4262 7615 -4204
rect 7649 -4262 7707 -4204
rect 7741 -4262 7799 -4204
rect 7833 -4262 7891 -4204
rect 7925 -4262 7983 -4204
rect 8017 -4262 8075 -4204
rect 8109 -4262 8167 -4204
rect 8201 -4262 8259 -4204
rect 8293 -4262 8351 -4204
rect 8385 -4262 8443 -4204
rect 8477 -4262 8535 -4204
rect 8569 -4262 8627 -4204
rect 8661 -4262 8719 -4204
rect 8753 -4262 8811 -4204
rect 8845 -4262 8903 -4204
rect 8937 -4262 8995 -4204
rect 9029 -4262 9087 -4204
rect 9121 -4262 9179 -4204
rect 9213 -4262 9271 -4204
rect 9305 -4262 9363 -4204
rect 9397 -4262 9455 -4204
rect 9489 -4262 9547 -4204
rect 9581 -4262 9639 -4204
rect 9673 -4262 9731 -4204
rect 9765 -4262 9823 -4204
rect 9857 -4262 9915 -4204
rect 9949 -4262 10007 -4204
rect 10041 -4262 10099 -4204
rect 10133 -4262 10191 -4204
rect 10225 -4262 10283 -4204
rect 10317 -4262 10375 -4204
rect 10409 -4262 10467 -4204
rect 10501 -4262 10559 -4204
rect 10593 -4262 10651 -4204
rect 10685 -4262 10743 -4204
rect 10777 -4262 10835 -4204
rect 10869 -4262 10927 -4204
rect 10961 -4262 11019 -4204
rect 11053 -4262 11111 -4204
rect 11145 -4262 11203 -4204
rect 11237 -4262 11295 -4204
rect 11329 -4262 11387 -4204
rect 11421 -4262 11479 -4204
rect 11513 -4262 11571 -4204
rect 11605 -4262 11663 -4204
rect 11697 -4262 11755 -4204
rect 11789 -4262 11847 -4204
rect 11881 -4262 11939 -4204
rect 11973 -4262 12031 -4204
rect 12065 -4262 12123 -4204
rect 12157 -4262 12215 -4204
rect 12249 -4262 12307 -4204
rect 12341 -4262 12399 -4204
rect 12433 -4262 12491 -4204
rect 12525 -4262 12583 -4204
rect 12617 -4262 12675 -4204
rect 12709 -4262 12767 -4204
rect 12801 -4262 12859 -4204
rect 12893 -4262 12951 -4204
rect 12985 -4262 13043 -4204
rect 13077 -4262 13135 -4204
rect 13169 -4262 13227 -4204
rect 13261 -4262 13319 -4204
rect 13353 -4262 13411 -4204
rect 13445 -4262 13503 -4204
rect 13537 -4262 13595 -4204
rect 13629 -4262 13687 -4204
rect 13721 -4262 13779 -4204
rect 13813 -4262 13871 -4204
rect 13905 -4262 13963 -4204
rect 13997 -4262 14055 -4204
rect 14089 -4262 14147 -4204
rect 14181 -4262 14239 -4204
rect 14273 -4262 14331 -4204
rect 14365 -4262 14423 -4204
rect 14457 -4262 14515 -4204
rect 14549 -4262 14607 -4204
rect 14641 -4262 14699 -4204
rect 14733 -4262 14791 -4204
rect 14825 -4262 14883 -4204
rect 14917 -4262 14975 -4204
rect 15009 -4262 15067 -4204
rect 15101 -4262 15159 -4204
rect 15193 -4262 15251 -4204
rect 15285 -4262 15343 -4204
rect 15377 -4262 15435 -4204
rect 15469 -4262 15527 -4204
rect 15561 -4262 15619 -4204
rect 15653 -4262 15711 -4204
rect 15745 -4262 15803 -4204
rect 15837 -4262 15895 -4204
rect 15929 -4262 15987 -4204
rect 16021 -4262 16079 -4204
rect 16113 -4262 16171 -4204
rect 16205 -4262 16263 -4204
rect 16297 -4262 16355 -4204
rect 16389 -4262 16447 -4204
rect 16481 -4262 16539 -4204
rect 16573 -4262 16631 -4204
rect 16665 -4262 16723 -4204
rect 16757 -4262 16815 -4204
rect 16849 -4262 16907 -4204
rect 16941 -4262 16999 -4204
rect 17033 -4262 17091 -4204
rect 17125 -4262 17183 -4204
rect 17217 -4262 17275 -4204
rect 17309 -4262 17367 -4204
rect 17401 -4262 17459 -4204
rect 17493 -4262 17551 -4204
rect 17585 -4262 17643 -4204
rect 17677 -4262 17735 -4204
rect 17769 -4262 17827 -4204
rect 17861 -4262 17919 -4204
rect 17953 -4262 18011 -4204
rect 18045 -4262 18103 -4204
rect 18137 -4262 18195 -4204
rect 18229 -4262 18287 -4204
rect 18321 -4262 18379 -4204
rect 18413 -4262 18471 -4204
rect 18505 -4262 18563 -4204
rect 18597 -4262 18655 -4204
rect 18689 -4262 18747 -4204
rect 18781 -4262 18839 -4204
rect 18873 -4262 18931 -4204
rect 18965 -4262 19023 -4204
rect 19057 -4262 19115 -4204
rect 19149 -4262 19207 -4204
rect 19241 -4262 19299 -4204
rect 19333 -4262 19391 -4204
rect 19425 -4262 19483 -4204
rect 19517 -4262 19575 -4204
rect 19609 -4262 19667 -4204
rect 19701 -4262 19759 -4204
rect 19793 -4262 19851 -4204
rect 19885 -4262 19943 -4204
rect 19977 -4262 20035 -4204
rect 20069 -4262 20127 -4204
rect 20161 -4262 20219 -4204
rect 20253 -4262 20311 -4204
rect 20345 -4262 20403 -4204
rect 20437 -4262 20495 -4204
rect 20529 -4262 20587 -4204
rect 20621 -4262 20679 -4204
rect 20713 -4262 20771 -4204
rect 20805 -4262 20863 -4204
rect 20897 -4262 20955 -4204
rect 20989 -4262 21047 -4204
rect 21081 -4262 21139 -4204
rect 21173 -4262 21231 -4204
rect 21265 -4262 21323 -4204
rect 21357 -4262 21415 -4204
rect 21449 -4262 21507 -4204
rect 21541 -4262 21599 -4204
rect 21633 -4262 21691 -4204
rect 21725 -4262 21783 -4204
rect 21817 -4262 21875 -4204
rect 21909 -4262 21967 -4204
rect 22001 -4262 22059 -4204
rect 22093 -4262 22151 -4204
rect 22185 -4262 22243 -4204
rect 22277 -4262 22335 -4204
rect 22369 -4262 22427 -4204
rect 22461 -4262 22519 -4204
rect 22553 -4262 22611 -4204
rect 22645 -4262 22703 -4204
rect 22737 -4262 22795 -4204
rect 22829 -4262 22887 -4204
rect 22921 -4262 22979 -4204
rect 23013 -4262 23071 -4204
rect 23105 -4262 23163 -4204
rect 23197 -4262 23255 -4204
rect 23289 -4262 23347 -4204
rect 23381 -4262 23439 -4204
rect 23473 -4262 23531 -4204
rect 23565 -4262 23623 -4204
rect 23657 -4262 23715 -4204
rect 23749 -4262 23807 -4204
rect 23841 -4262 23899 -4204
rect 23933 -4262 23991 -4204
rect 24025 -4262 24083 -4204
rect 24117 -4262 24175 -4204
rect 24209 -4262 24267 -4204
rect 24301 -4262 24359 -4204
rect 24393 -4262 24451 -4204
rect 24485 -4262 24543 -4204
rect 24577 -4262 24635 -4204
rect 24669 -4262 24727 -4204
rect 24761 -4262 24819 -4204
rect 24853 -4262 24911 -4204
rect 24945 -4262 25003 -4204
rect 25037 -4262 25095 -4204
rect 25129 -4262 25187 -4204
rect 25221 -4262 25279 -4204
rect 25313 -4262 25371 -4204
rect 25405 -4262 25463 -4204
rect 25497 -4262 25555 -4204
rect 25589 -4262 25647 -4204
rect 25681 -4262 25739 -4204
rect 25773 -4262 25831 -4204
rect 25865 -4262 25923 -4204
rect 25957 -4262 26015 -4204
rect 26049 -4262 26107 -4204
rect 26141 -4262 26199 -4204
rect 26233 -4262 26291 -4204
rect 26325 -4262 26383 -4204
rect 26417 -4262 26475 -4204
rect 26509 -4262 26567 -4204
rect 26601 -4262 26659 -4204
rect 26693 -4262 26751 -4204
rect 26785 -4262 26843 -4204
rect 26877 -4262 26935 -4204
rect 26969 -4262 27027 -4204
rect 27061 -4262 27119 -4204
rect 27153 -4262 27211 -4204
rect 27245 -4262 27303 -4204
rect 27337 -4262 27395 -4204
rect 27429 -4262 27487 -4204
rect 27521 -4262 27579 -4204
rect 27613 -4262 27671 -4204
rect 27705 -4262 27763 -4204
rect 27797 -4262 27855 -4204
rect 27889 -4262 27947 -4204
rect 27981 -4262 28039 -4204
rect 28073 -4262 28131 -4204
rect 28165 -4262 28223 -4204
rect 28257 -4262 28315 -4204
rect 28349 -4262 28407 -4204
rect 28441 -4262 28499 -4204
rect 28533 -4262 28591 -4204
rect 28625 -4262 28683 -4204
rect 28717 -4262 28775 -4204
rect 28809 -4262 28867 -4204
rect 28901 -4262 28959 -4204
rect 28993 -4262 29051 -4204
rect 29085 -4262 29143 -4204
rect 29177 -4262 29235 -4204
rect 29269 -4262 29327 -4204
rect 29361 -4262 29419 -4204
rect 29453 -4262 29511 -4204
rect 29545 -4262 29603 -4204
rect 29637 -4262 29695 -4204
rect 29729 -4262 29787 -4204
rect 29821 -4262 29879 -4204
rect 29913 -4262 29971 -4204
rect 30005 -4262 30063 -4204
rect 30097 -4262 30155 -4204
rect 30189 -4262 30247 -4204
rect 30281 -4262 30339 -4204
rect 30373 -4262 30431 -4204
rect 30465 -4262 30523 -4204
rect 30557 -4262 30615 -4204
rect 30649 -4262 30707 -4204
rect 30741 -4262 30799 -4204
rect 30833 -4262 30891 -4204
rect 30925 -4262 30983 -4204
rect 31017 -4262 31075 -4204
rect 31109 -4262 31167 -4204
rect 31201 -4262 31259 -4204
rect 31293 -4262 31351 -4204
rect 31385 -4262 31443 -4204
rect 31477 -4262 31535 -4204
rect 31569 -4262 31627 -4204
rect 31661 -4262 31719 -4204
rect 31753 -4262 31811 -4204
rect 31845 -4262 31903 -4204
rect 31937 -4262 31995 -4204
rect 32029 -4262 32087 -4204
rect 32121 -4262 32179 -4204
rect 32213 -4262 32271 -4204
rect 32305 -4262 32363 -4204
rect 32397 -4262 32455 -4204
rect 32489 -4262 32547 -4204
rect 32581 -4262 32639 -4204
rect 32673 -4262 32731 -4204
rect 32765 -4262 32823 -4204
rect 32857 -4262 32915 -4204
rect 32949 -4262 33007 -4204
rect 33041 -4262 33099 -4204
rect 33133 -4262 33162 -4204
rect -9140 -4312 -9089 -4296
rect -9140 -4346 -9123 -4312
rect -9140 -4380 -9089 -4346
rect -9055 -4328 -8989 -4262
rect -9055 -4362 -9039 -4328
rect -9005 -4362 -8989 -4328
rect -8955 -4312 -8921 -4296
rect -9140 -4414 -9123 -4380
rect -8955 -4380 -8921 -4346
rect -9089 -4414 -8990 -4396
rect -9140 -4430 -8990 -4414
rect -9158 -4540 -9070 -4464
rect -9158 -4574 -9126 -4540
rect -9092 -4574 -9070 -4540
rect -9158 -4594 -9070 -4574
rect -9036 -4525 -8990 -4430
rect -9036 -4534 -9024 -4525
rect -9002 -4568 -8990 -4559
rect -9036 -4628 -8990 -4568
rect -9140 -4662 -8990 -4628
rect -9140 -4670 -9089 -4662
rect -9140 -4704 -9123 -4670
rect -8955 -4670 -8921 -4432
rect -8887 -4456 -8822 -4299
rect -8788 -4304 -8738 -4262
rect -8788 -4338 -8772 -4304
rect -8788 -4354 -8738 -4338
rect -8704 -4312 -8654 -4296
rect -8704 -4346 -8688 -4312
rect -8704 -4362 -8654 -4346
rect -8611 -4306 -8475 -4296
rect -8611 -4340 -8595 -4306
rect -8561 -4340 -8475 -4306
rect -8360 -4314 -8294 -4262
rect -8167 -4304 -8093 -4262
rect -8611 -4362 -8475 -4340
rect -8704 -4388 -8670 -4362
rect -8749 -4422 -8670 -4388
rect -8636 -4398 -8543 -4396
rect -8875 -4479 -8783 -4456
rect -8875 -4513 -8817 -4479
rect -8875 -4614 -8783 -4513
rect -8875 -4648 -8851 -4614
rect -8813 -4648 -8783 -4614
rect -8875 -4666 -8783 -4648
rect -9140 -4720 -9089 -4704
rect -9055 -4730 -9039 -4696
rect -9005 -4730 -8989 -4696
rect -8749 -4694 -8715 -4422
rect -8636 -4424 -8577 -4398
rect -8602 -4432 -8577 -4424
rect -8602 -4458 -8543 -4432
rect -8636 -4474 -8543 -4458
rect -8681 -4534 -8611 -4512
rect -8681 -4568 -8669 -4534
rect -8635 -4568 -8611 -4534
rect -8681 -4586 -8611 -4568
rect -8681 -4620 -8658 -4586
rect -8624 -4620 -8611 -4586
rect -8681 -4636 -8611 -4620
rect -8577 -4592 -8543 -4474
rect -8509 -4518 -8475 -4362
rect -8441 -4330 -8407 -4314
rect -8360 -4348 -8344 -4314
rect -8310 -4348 -8294 -4314
rect -8260 -4330 -8226 -4314
rect -8441 -4382 -8407 -4364
rect -8167 -4338 -8147 -4304
rect -8113 -4338 -8093 -4304
rect -8167 -4354 -8093 -4338
rect -8059 -4312 -8025 -4296
rect -8260 -4382 -8226 -4364
rect -8441 -4416 -8226 -4382
rect -8059 -4388 -8025 -4346
rect -7978 -4305 -7804 -4296
rect -7978 -4339 -7962 -4305
rect -7928 -4339 -7804 -4305
rect -7978 -4364 -7804 -4339
rect -7770 -4304 -7720 -4262
rect -7736 -4338 -7720 -4304
rect -7616 -4304 -7472 -4262
rect -7770 -4354 -7720 -4338
rect -7686 -4330 -7652 -4314
rect -8137 -4422 -8025 -4388
rect -8137 -4450 -8103 -4422
rect -8403 -4484 -8387 -4450
rect -8353 -4484 -8103 -4450
rect -7964 -4432 -7953 -4398
rect -7919 -4424 -7872 -4398
rect -7964 -4456 -7922 -4432
rect -8509 -4538 -8171 -4518
rect -8509 -4552 -8205 -4538
rect -8577 -4626 -8556 -4592
rect -8522 -4626 -8506 -4592
rect -8577 -4636 -8506 -4626
rect -8472 -4694 -8438 -4552
rect -8397 -4602 -8301 -4586
rect -8363 -4636 -8325 -4602
rect -8267 -4620 -8239 -4586
rect -8205 -4588 -8171 -4572
rect -8291 -4636 -8239 -4620
rect -8137 -4622 -8103 -4484
rect -8955 -4720 -8921 -4704
rect -9055 -4772 -8989 -4730
rect -8849 -4734 -8833 -4700
rect -8799 -4734 -8783 -4700
rect -8749 -4728 -8700 -4694
rect -8666 -4728 -8650 -4694
rect -8609 -4728 -8593 -4694
rect -8559 -4728 -8438 -4694
rect -8263 -4696 -8197 -4680
rect -8849 -4772 -8783 -4734
rect -8263 -4730 -8247 -4696
rect -8213 -4730 -8197 -4696
rect -8263 -4772 -8197 -4730
rect -8155 -4700 -8103 -4622
rect -8065 -4458 -7922 -4456
rect -7888 -4458 -7872 -4424
rect -7838 -4440 -7804 -4364
rect -7616 -4338 -7600 -4304
rect -7566 -4338 -7522 -4304
rect -7488 -4338 -7472 -4304
rect -7438 -4312 -7357 -4296
rect -7206 -4304 -7172 -4262
rect -7686 -4372 -7652 -4364
rect -7404 -4346 -7357 -4312
rect -7686 -4406 -7526 -4372
rect -8065 -4490 -7930 -4458
rect -7838 -4474 -7644 -4440
rect -7610 -4474 -7594 -4440
rect -8065 -4598 -8023 -4490
rect -7838 -4492 -7804 -4474
rect -8065 -4632 -8057 -4598
rect -8065 -4648 -8023 -4632
rect -7989 -4534 -7919 -4524
rect -7989 -4550 -7953 -4534
rect -7989 -4584 -7961 -4550
rect -7927 -4584 -7919 -4568
rect -7989 -4648 -7919 -4584
rect -7885 -4526 -7804 -4492
rect -7885 -4682 -7851 -4526
rect -7737 -4539 -7629 -4508
rect -7560 -4524 -7526 -4406
rect -7438 -4380 -7357 -4346
rect -7404 -4414 -7357 -4380
rect -7438 -4448 -7357 -4414
rect -7404 -4482 -7357 -4448
rect -7438 -4498 -7357 -4482
rect -7560 -4530 -7471 -4524
rect -7703 -4548 -7629 -4539
rect -7817 -4576 -7773 -4560
rect -7783 -4610 -7773 -4576
rect -7737 -4582 -7721 -4573
rect -7687 -4582 -7629 -4548
rect -7817 -4616 -7773 -4610
rect -7677 -4602 -7629 -4582
rect -7817 -4650 -7711 -4616
rect -8041 -4696 -7851 -4682
rect -8155 -4734 -8135 -4700
rect -8101 -4734 -8085 -4700
rect -8041 -4730 -8025 -4696
rect -7991 -4730 -7851 -4696
rect -8041 -4738 -7851 -4730
rect -7817 -4700 -7779 -4684
rect -7817 -4734 -7813 -4700
rect -7745 -4696 -7711 -4650
rect -7643 -4636 -7629 -4602
rect -7677 -4662 -7629 -4636
rect -7595 -4540 -7471 -4530
rect -7595 -4574 -7521 -4540
rect -7487 -4574 -7471 -4540
rect -7595 -4590 -7471 -4574
rect -7595 -4625 -7530 -4590
rect -7423 -4624 -7357 -4498
rect -7595 -4680 -7531 -4625
rect -7745 -4714 -7595 -4696
rect -7561 -4714 -7531 -4680
rect -7745 -4730 -7531 -4714
rect -7491 -4657 -7457 -4635
rect -7817 -4772 -7779 -4734
rect -7491 -4772 -7457 -4691
rect -7423 -4658 -7407 -4624
rect -7373 -4658 -7357 -4624
rect -7423 -4692 -7357 -4658
rect -7423 -4726 -7407 -4692
rect -7373 -4726 -7357 -4692
rect -7319 -4338 -7303 -4304
rect -7269 -4338 -7253 -4304
rect -7319 -4372 -7253 -4338
rect -7319 -4406 -7303 -4372
rect -7269 -4406 -7253 -4372
rect -7319 -4524 -7253 -4406
rect -7024 -4312 -6973 -4296
rect -7206 -4372 -7172 -4338
rect -7206 -4440 -7172 -4406
rect -7206 -4490 -7172 -4474
rect -7122 -4340 -7071 -4324
rect -7088 -4374 -7071 -4340
rect -7122 -4408 -7071 -4374
rect -7088 -4442 -7071 -4408
rect -7024 -4346 -7007 -4312
rect -7024 -4380 -6973 -4346
rect -6939 -4328 -6873 -4262
rect -6939 -4362 -6923 -4328
rect -6889 -4362 -6873 -4328
rect -6839 -4312 -6805 -4296
rect -7024 -4414 -7007 -4380
rect -6839 -4380 -6805 -4346
rect -6973 -4414 -6874 -4396
rect -7024 -4430 -6874 -4414
rect -7122 -4464 -7071 -4442
rect -7122 -4500 -6954 -4464
rect -7113 -4515 -6954 -4500
rect -7319 -4540 -7147 -4524
rect -7319 -4574 -7181 -4540
rect -7319 -4590 -7147 -4574
rect -7113 -4549 -7082 -4515
rect -7044 -4540 -6954 -4515
rect -7044 -4549 -7010 -4540
rect -7113 -4574 -7010 -4549
rect -6976 -4574 -6954 -4540
rect -7319 -4670 -7269 -4590
rect -7113 -4594 -6954 -4574
rect -6920 -4525 -6874 -4430
rect -6920 -4534 -6908 -4525
rect -6886 -4568 -6874 -4559
rect -7113 -4630 -7071 -4594
rect -6920 -4628 -6874 -4568
rect -7122 -4646 -7071 -4630
rect -7319 -4704 -7303 -4670
rect -7319 -4720 -7269 -4704
rect -7206 -4676 -7172 -4653
rect -7423 -4734 -7357 -4726
rect -7206 -4772 -7172 -4710
rect -7088 -4680 -7071 -4646
rect -7122 -4736 -7071 -4680
rect -7024 -4662 -6874 -4628
rect -7024 -4670 -6973 -4662
rect -7024 -4704 -7007 -4670
rect -6839 -4670 -6805 -4432
rect -6771 -4456 -6706 -4299
rect -6672 -4304 -6622 -4262
rect -6672 -4338 -6656 -4304
rect -6672 -4354 -6622 -4338
rect -6588 -4312 -6538 -4296
rect -6588 -4346 -6572 -4312
rect -6588 -4362 -6538 -4346
rect -6495 -4306 -6359 -4296
rect -6495 -4340 -6479 -4306
rect -6445 -4340 -6359 -4306
rect -6244 -4314 -6178 -4262
rect -6051 -4304 -5977 -4262
rect -6495 -4362 -6359 -4340
rect -6588 -4388 -6554 -4362
rect -6633 -4422 -6554 -4388
rect -6520 -4398 -6427 -4396
rect -6759 -4479 -6667 -4456
rect -6759 -4513 -6701 -4479
rect -6759 -4614 -6667 -4513
rect -6759 -4648 -6735 -4614
rect -6697 -4648 -6667 -4614
rect -6759 -4666 -6667 -4648
rect -7024 -4720 -6973 -4704
rect -6939 -4730 -6923 -4696
rect -6889 -4730 -6873 -4696
rect -6633 -4694 -6599 -4422
rect -6520 -4424 -6461 -4398
rect -6486 -4432 -6461 -4424
rect -6486 -4458 -6427 -4432
rect -6520 -4474 -6427 -4458
rect -6565 -4534 -6495 -4512
rect -6565 -4568 -6553 -4534
rect -6519 -4568 -6495 -4534
rect -6565 -4586 -6495 -4568
rect -6565 -4620 -6542 -4586
rect -6508 -4620 -6495 -4586
rect -6565 -4636 -6495 -4620
rect -6461 -4592 -6427 -4474
rect -6393 -4518 -6359 -4362
rect -6325 -4330 -6291 -4314
rect -6244 -4348 -6228 -4314
rect -6194 -4348 -6178 -4314
rect -6144 -4330 -6110 -4314
rect -6325 -4382 -6291 -4364
rect -6051 -4338 -6031 -4304
rect -5997 -4338 -5977 -4304
rect -6051 -4354 -5977 -4338
rect -5943 -4312 -5909 -4296
rect -6144 -4382 -6110 -4364
rect -6325 -4416 -6110 -4382
rect -5943 -4388 -5909 -4346
rect -5862 -4305 -5688 -4296
rect -5862 -4339 -5846 -4305
rect -5812 -4339 -5688 -4305
rect -5862 -4364 -5688 -4339
rect -5654 -4304 -5604 -4262
rect -5620 -4338 -5604 -4304
rect -5500 -4304 -5356 -4262
rect -5654 -4354 -5604 -4338
rect -5570 -4330 -5536 -4314
rect -6021 -4422 -5909 -4388
rect -6021 -4450 -5987 -4422
rect -6287 -4484 -6271 -4450
rect -6237 -4484 -5987 -4450
rect -5848 -4432 -5837 -4398
rect -5803 -4424 -5756 -4398
rect -5848 -4456 -5806 -4432
rect -6393 -4538 -6055 -4518
rect -6393 -4552 -6089 -4538
rect -6461 -4626 -6440 -4592
rect -6406 -4626 -6390 -4592
rect -6461 -4636 -6390 -4626
rect -6356 -4694 -6322 -4552
rect -6281 -4602 -6185 -4586
rect -6247 -4636 -6209 -4602
rect -6151 -4620 -6123 -4586
rect -6089 -4588 -6055 -4572
rect -6175 -4636 -6123 -4620
rect -6021 -4622 -5987 -4484
rect -6839 -4720 -6805 -4704
rect -6939 -4772 -6873 -4730
rect -6733 -4734 -6717 -4700
rect -6683 -4734 -6667 -4700
rect -6633 -4728 -6584 -4694
rect -6550 -4728 -6534 -4694
rect -6493 -4728 -6477 -4694
rect -6443 -4728 -6322 -4694
rect -6147 -4696 -6081 -4680
rect -6733 -4772 -6667 -4734
rect -6147 -4730 -6131 -4696
rect -6097 -4730 -6081 -4696
rect -6147 -4772 -6081 -4730
rect -6039 -4700 -5987 -4622
rect -5949 -4458 -5806 -4456
rect -5772 -4458 -5756 -4424
rect -5722 -4440 -5688 -4364
rect -5500 -4338 -5484 -4304
rect -5450 -4338 -5406 -4304
rect -5372 -4338 -5356 -4304
rect -5322 -4312 -5241 -4296
rect -5090 -4304 -5056 -4262
rect -5570 -4372 -5536 -4364
rect -5288 -4346 -5241 -4312
rect -5570 -4406 -5410 -4372
rect -5949 -4490 -5814 -4458
rect -5722 -4474 -5528 -4440
rect -5494 -4474 -5478 -4440
rect -5949 -4598 -5907 -4490
rect -5722 -4492 -5688 -4474
rect -5949 -4632 -5941 -4598
rect -5949 -4648 -5907 -4632
rect -5873 -4534 -5803 -4524
rect -5873 -4550 -5837 -4534
rect -5873 -4584 -5845 -4550
rect -5811 -4584 -5803 -4568
rect -5873 -4648 -5803 -4584
rect -5769 -4526 -5688 -4492
rect -5769 -4682 -5735 -4526
rect -5621 -4539 -5513 -4508
rect -5444 -4524 -5410 -4406
rect -5322 -4380 -5241 -4346
rect -5288 -4414 -5241 -4380
rect -5322 -4448 -5241 -4414
rect -5288 -4482 -5241 -4448
rect -5322 -4498 -5241 -4482
rect -5444 -4530 -5355 -4524
rect -5587 -4548 -5513 -4539
rect -5701 -4576 -5657 -4560
rect -5667 -4610 -5657 -4576
rect -5621 -4582 -5605 -4573
rect -5571 -4582 -5513 -4548
rect -5701 -4616 -5657 -4610
rect -5561 -4602 -5513 -4582
rect -5701 -4650 -5595 -4616
rect -5925 -4696 -5735 -4682
rect -6039 -4734 -6019 -4700
rect -5985 -4734 -5969 -4700
rect -5925 -4730 -5909 -4696
rect -5875 -4730 -5735 -4696
rect -5925 -4738 -5735 -4730
rect -5701 -4700 -5663 -4684
rect -5701 -4734 -5697 -4700
rect -5629 -4696 -5595 -4650
rect -5527 -4636 -5513 -4602
rect -5561 -4662 -5513 -4636
rect -5479 -4540 -5355 -4530
rect -5479 -4574 -5405 -4540
rect -5371 -4574 -5355 -4540
rect -5479 -4590 -5355 -4574
rect -5479 -4625 -5414 -4590
rect -5307 -4624 -5241 -4498
rect -5479 -4680 -5415 -4625
rect -5629 -4714 -5479 -4696
rect -5445 -4714 -5415 -4680
rect -5629 -4730 -5415 -4714
rect -5375 -4657 -5341 -4635
rect -5701 -4772 -5663 -4734
rect -5375 -4772 -5341 -4691
rect -5307 -4658 -5291 -4624
rect -5257 -4658 -5241 -4624
rect -5307 -4692 -5241 -4658
rect -5307 -4726 -5291 -4692
rect -5257 -4726 -5241 -4692
rect -5203 -4338 -5187 -4304
rect -5153 -4338 -5137 -4304
rect -5203 -4372 -5137 -4338
rect -5203 -4406 -5187 -4372
rect -5153 -4406 -5137 -4372
rect -5203 -4524 -5137 -4406
rect -4908 -4312 -4857 -4296
rect -5090 -4372 -5056 -4338
rect -5090 -4440 -5056 -4406
rect -5090 -4490 -5056 -4474
rect -5006 -4340 -4955 -4324
rect -4972 -4374 -4955 -4340
rect -5006 -4408 -4955 -4374
rect -4972 -4442 -4955 -4408
rect -4908 -4346 -4891 -4312
rect -4908 -4380 -4857 -4346
rect -4823 -4328 -4757 -4262
rect -4823 -4362 -4807 -4328
rect -4773 -4362 -4757 -4328
rect -4723 -4312 -4689 -4296
rect -4908 -4414 -4891 -4380
rect -4723 -4380 -4689 -4346
rect -4857 -4414 -4758 -4396
rect -4908 -4430 -4758 -4414
rect -5006 -4464 -4955 -4442
rect -5006 -4500 -4838 -4464
rect -4997 -4515 -4838 -4500
rect -5203 -4540 -5031 -4524
rect -5203 -4574 -5065 -4540
rect -5203 -4590 -5031 -4574
rect -4997 -4549 -4966 -4515
rect -4928 -4540 -4838 -4515
rect -4928 -4549 -4894 -4540
rect -4997 -4574 -4894 -4549
rect -4860 -4574 -4838 -4540
rect -5203 -4670 -5153 -4590
rect -4997 -4594 -4838 -4574
rect -4804 -4525 -4758 -4430
rect -4804 -4534 -4792 -4525
rect -4770 -4568 -4758 -4559
rect -4997 -4630 -4955 -4594
rect -4804 -4628 -4758 -4568
rect -5006 -4646 -4955 -4630
rect -5203 -4704 -5187 -4670
rect -5203 -4720 -5153 -4704
rect -5090 -4676 -5056 -4653
rect -5307 -4734 -5241 -4726
rect -5090 -4772 -5056 -4710
rect -4972 -4680 -4955 -4646
rect -5006 -4736 -4955 -4680
rect -4908 -4662 -4758 -4628
rect -4908 -4670 -4857 -4662
rect -4908 -4704 -4891 -4670
rect -4723 -4670 -4689 -4432
rect -4655 -4456 -4590 -4299
rect -4556 -4304 -4506 -4262
rect -4556 -4338 -4540 -4304
rect -4556 -4354 -4506 -4338
rect -4472 -4312 -4422 -4296
rect -4472 -4346 -4456 -4312
rect -4472 -4362 -4422 -4346
rect -4379 -4306 -4243 -4296
rect -4379 -4340 -4363 -4306
rect -4329 -4340 -4243 -4306
rect -4128 -4314 -4062 -4262
rect -3935 -4304 -3861 -4262
rect -4379 -4362 -4243 -4340
rect -4472 -4388 -4438 -4362
rect -4517 -4422 -4438 -4388
rect -4404 -4398 -4311 -4396
rect -4643 -4479 -4551 -4456
rect -4643 -4513 -4585 -4479
rect -4643 -4614 -4551 -4513
rect -4643 -4648 -4619 -4614
rect -4581 -4648 -4551 -4614
rect -4643 -4666 -4551 -4648
rect -4908 -4720 -4857 -4704
rect -4823 -4730 -4807 -4696
rect -4773 -4730 -4757 -4696
rect -4517 -4694 -4483 -4422
rect -4404 -4424 -4345 -4398
rect -4370 -4432 -4345 -4424
rect -4370 -4458 -4311 -4432
rect -4404 -4474 -4311 -4458
rect -4449 -4534 -4379 -4512
rect -4449 -4568 -4437 -4534
rect -4403 -4568 -4379 -4534
rect -4449 -4586 -4379 -4568
rect -4449 -4620 -4426 -4586
rect -4392 -4620 -4379 -4586
rect -4449 -4636 -4379 -4620
rect -4345 -4592 -4311 -4474
rect -4277 -4518 -4243 -4362
rect -4209 -4330 -4175 -4314
rect -4128 -4348 -4112 -4314
rect -4078 -4348 -4062 -4314
rect -4028 -4330 -3994 -4314
rect -4209 -4382 -4175 -4364
rect -3935 -4338 -3915 -4304
rect -3881 -4338 -3861 -4304
rect -3935 -4354 -3861 -4338
rect -3827 -4312 -3793 -4296
rect -4028 -4382 -3994 -4364
rect -4209 -4416 -3994 -4382
rect -3827 -4388 -3793 -4346
rect -3746 -4305 -3572 -4296
rect -3746 -4339 -3730 -4305
rect -3696 -4339 -3572 -4305
rect -3746 -4364 -3572 -4339
rect -3538 -4304 -3488 -4262
rect -3504 -4338 -3488 -4304
rect -3384 -4304 -3240 -4262
rect -3538 -4354 -3488 -4338
rect -3454 -4330 -3420 -4314
rect -3905 -4422 -3793 -4388
rect -3905 -4450 -3871 -4422
rect -4171 -4484 -4155 -4450
rect -4121 -4484 -3871 -4450
rect -3732 -4432 -3721 -4398
rect -3687 -4424 -3640 -4398
rect -3732 -4456 -3690 -4432
rect -4277 -4538 -3939 -4518
rect -4277 -4552 -3973 -4538
rect -4345 -4626 -4324 -4592
rect -4290 -4626 -4274 -4592
rect -4345 -4636 -4274 -4626
rect -4240 -4694 -4206 -4552
rect -4165 -4602 -4069 -4586
rect -4131 -4636 -4093 -4602
rect -4035 -4620 -4007 -4586
rect -3973 -4588 -3939 -4572
rect -4059 -4636 -4007 -4620
rect -3905 -4622 -3871 -4484
rect -4723 -4720 -4689 -4704
rect -4823 -4772 -4757 -4730
rect -4617 -4734 -4601 -4700
rect -4567 -4734 -4551 -4700
rect -4517 -4728 -4468 -4694
rect -4434 -4728 -4418 -4694
rect -4377 -4728 -4361 -4694
rect -4327 -4728 -4206 -4694
rect -4031 -4696 -3965 -4680
rect -4617 -4772 -4551 -4734
rect -4031 -4730 -4015 -4696
rect -3981 -4730 -3965 -4696
rect -4031 -4772 -3965 -4730
rect -3923 -4700 -3871 -4622
rect -3833 -4458 -3690 -4456
rect -3656 -4458 -3640 -4424
rect -3606 -4440 -3572 -4364
rect -3384 -4338 -3368 -4304
rect -3334 -4338 -3290 -4304
rect -3256 -4338 -3240 -4304
rect -3206 -4312 -3125 -4296
rect -2974 -4304 -2940 -4262
rect -3454 -4372 -3420 -4364
rect -3172 -4346 -3125 -4312
rect -3454 -4406 -3294 -4372
rect -3833 -4490 -3698 -4458
rect -3606 -4474 -3412 -4440
rect -3378 -4474 -3362 -4440
rect -3833 -4598 -3791 -4490
rect -3606 -4492 -3572 -4474
rect -3833 -4632 -3825 -4598
rect -3833 -4648 -3791 -4632
rect -3757 -4534 -3687 -4524
rect -3757 -4550 -3721 -4534
rect -3757 -4584 -3729 -4550
rect -3695 -4584 -3687 -4568
rect -3757 -4648 -3687 -4584
rect -3653 -4526 -3572 -4492
rect -3653 -4682 -3619 -4526
rect -3505 -4539 -3397 -4508
rect -3328 -4524 -3294 -4406
rect -3206 -4380 -3125 -4346
rect -3172 -4414 -3125 -4380
rect -3206 -4448 -3125 -4414
rect -3172 -4482 -3125 -4448
rect -3206 -4498 -3125 -4482
rect -3328 -4530 -3239 -4524
rect -3471 -4548 -3397 -4539
rect -3585 -4576 -3541 -4560
rect -3551 -4610 -3541 -4576
rect -3505 -4582 -3489 -4573
rect -3455 -4582 -3397 -4548
rect -3585 -4616 -3541 -4610
rect -3445 -4602 -3397 -4582
rect -3585 -4650 -3479 -4616
rect -3809 -4696 -3619 -4682
rect -3923 -4734 -3903 -4700
rect -3869 -4734 -3853 -4700
rect -3809 -4730 -3793 -4696
rect -3759 -4730 -3619 -4696
rect -3809 -4738 -3619 -4730
rect -3585 -4700 -3547 -4684
rect -3585 -4734 -3581 -4700
rect -3513 -4696 -3479 -4650
rect -3411 -4636 -3397 -4602
rect -3445 -4662 -3397 -4636
rect -3363 -4540 -3239 -4530
rect -3363 -4574 -3289 -4540
rect -3255 -4574 -3239 -4540
rect -3363 -4590 -3239 -4574
rect -3363 -4625 -3298 -4590
rect -3191 -4624 -3125 -4498
rect -3363 -4680 -3299 -4625
rect -3513 -4714 -3363 -4696
rect -3329 -4714 -3299 -4680
rect -3513 -4730 -3299 -4714
rect -3259 -4657 -3225 -4635
rect -3585 -4772 -3547 -4734
rect -3259 -4772 -3225 -4691
rect -3191 -4658 -3175 -4624
rect -3141 -4658 -3125 -4624
rect -3191 -4692 -3125 -4658
rect -3191 -4726 -3175 -4692
rect -3141 -4726 -3125 -4692
rect -3087 -4338 -3071 -4304
rect -3037 -4338 -3021 -4304
rect -3087 -4372 -3021 -4338
rect -3087 -4406 -3071 -4372
rect -3037 -4406 -3021 -4372
rect -3087 -4524 -3021 -4406
rect -2792 -4312 -2741 -4296
rect -2974 -4372 -2940 -4338
rect -2974 -4440 -2940 -4406
rect -2974 -4490 -2940 -4474
rect -2890 -4340 -2839 -4324
rect -2856 -4374 -2839 -4340
rect -2890 -4408 -2839 -4374
rect -2856 -4442 -2839 -4408
rect -2792 -4346 -2775 -4312
rect -2792 -4380 -2741 -4346
rect -2707 -4328 -2641 -4262
rect -2707 -4362 -2691 -4328
rect -2657 -4362 -2641 -4328
rect -2607 -4312 -2573 -4296
rect -2792 -4414 -2775 -4380
rect -2607 -4380 -2573 -4346
rect -2741 -4414 -2642 -4396
rect -2792 -4430 -2642 -4414
rect -2890 -4464 -2839 -4442
rect -2890 -4500 -2722 -4464
rect -2881 -4515 -2722 -4500
rect -3087 -4540 -2915 -4524
rect -3087 -4574 -2949 -4540
rect -3087 -4590 -2915 -4574
rect -2881 -4549 -2850 -4515
rect -2812 -4540 -2722 -4515
rect -2812 -4549 -2778 -4540
rect -2881 -4574 -2778 -4549
rect -2744 -4574 -2722 -4540
rect -3087 -4670 -3037 -4590
rect -2881 -4594 -2722 -4574
rect -2688 -4525 -2642 -4430
rect -2688 -4534 -2676 -4525
rect -2654 -4568 -2642 -4559
rect -2881 -4630 -2839 -4594
rect -2688 -4628 -2642 -4568
rect -2890 -4646 -2839 -4630
rect -3087 -4704 -3071 -4670
rect -3087 -4720 -3037 -4704
rect -2974 -4676 -2940 -4653
rect -3191 -4734 -3125 -4726
rect -2974 -4772 -2940 -4710
rect -2856 -4680 -2839 -4646
rect -2890 -4736 -2839 -4680
rect -2792 -4662 -2642 -4628
rect -2792 -4670 -2741 -4662
rect -2792 -4704 -2775 -4670
rect -2607 -4670 -2573 -4432
rect -2539 -4456 -2474 -4299
rect -2440 -4304 -2390 -4262
rect -2440 -4338 -2424 -4304
rect -2440 -4354 -2390 -4338
rect -2356 -4312 -2306 -4296
rect -2356 -4346 -2340 -4312
rect -2356 -4362 -2306 -4346
rect -2263 -4306 -2127 -4296
rect -2263 -4340 -2247 -4306
rect -2213 -4340 -2127 -4306
rect -2012 -4314 -1946 -4262
rect -1819 -4304 -1745 -4262
rect -2263 -4362 -2127 -4340
rect -2356 -4388 -2322 -4362
rect -2401 -4422 -2322 -4388
rect -2288 -4398 -2195 -4396
rect -2527 -4479 -2435 -4456
rect -2527 -4513 -2469 -4479
rect -2527 -4614 -2435 -4513
rect -2527 -4648 -2503 -4614
rect -2465 -4648 -2435 -4614
rect -2527 -4666 -2435 -4648
rect -2792 -4720 -2741 -4704
rect -2707 -4730 -2691 -4696
rect -2657 -4730 -2641 -4696
rect -2401 -4694 -2367 -4422
rect -2288 -4424 -2229 -4398
rect -2254 -4432 -2229 -4424
rect -2254 -4458 -2195 -4432
rect -2288 -4474 -2195 -4458
rect -2333 -4534 -2263 -4512
rect -2333 -4568 -2321 -4534
rect -2287 -4568 -2263 -4534
rect -2333 -4586 -2263 -4568
rect -2333 -4620 -2310 -4586
rect -2276 -4620 -2263 -4586
rect -2333 -4636 -2263 -4620
rect -2229 -4592 -2195 -4474
rect -2161 -4518 -2127 -4362
rect -2093 -4330 -2059 -4314
rect -2012 -4348 -1996 -4314
rect -1962 -4348 -1946 -4314
rect -1912 -4330 -1878 -4314
rect -2093 -4382 -2059 -4364
rect -1819 -4338 -1799 -4304
rect -1765 -4338 -1745 -4304
rect -1819 -4354 -1745 -4338
rect -1711 -4312 -1677 -4296
rect -1912 -4382 -1878 -4364
rect -2093 -4416 -1878 -4382
rect -1711 -4388 -1677 -4346
rect -1630 -4305 -1456 -4296
rect -1630 -4339 -1614 -4305
rect -1580 -4339 -1456 -4305
rect -1630 -4364 -1456 -4339
rect -1422 -4304 -1372 -4262
rect -1388 -4338 -1372 -4304
rect -1268 -4304 -1124 -4262
rect -1422 -4354 -1372 -4338
rect -1338 -4330 -1304 -4314
rect -1789 -4422 -1677 -4388
rect -1789 -4450 -1755 -4422
rect -2055 -4484 -2039 -4450
rect -2005 -4484 -1755 -4450
rect -1616 -4432 -1605 -4398
rect -1571 -4424 -1524 -4398
rect -1616 -4456 -1574 -4432
rect -2161 -4538 -1823 -4518
rect -2161 -4552 -1857 -4538
rect -2229 -4626 -2208 -4592
rect -2174 -4626 -2158 -4592
rect -2229 -4636 -2158 -4626
rect -2124 -4694 -2090 -4552
rect -2049 -4602 -1953 -4586
rect -2015 -4636 -1977 -4602
rect -1919 -4620 -1891 -4586
rect -1857 -4588 -1823 -4572
rect -1943 -4636 -1891 -4620
rect -1789 -4622 -1755 -4484
rect -2607 -4720 -2573 -4704
rect -2707 -4772 -2641 -4730
rect -2501 -4734 -2485 -4700
rect -2451 -4734 -2435 -4700
rect -2401 -4728 -2352 -4694
rect -2318 -4728 -2302 -4694
rect -2261 -4728 -2245 -4694
rect -2211 -4728 -2090 -4694
rect -1915 -4696 -1849 -4680
rect -2501 -4772 -2435 -4734
rect -1915 -4730 -1899 -4696
rect -1865 -4730 -1849 -4696
rect -1915 -4772 -1849 -4730
rect -1807 -4700 -1755 -4622
rect -1717 -4458 -1574 -4456
rect -1540 -4458 -1524 -4424
rect -1490 -4440 -1456 -4364
rect -1268 -4338 -1252 -4304
rect -1218 -4338 -1174 -4304
rect -1140 -4338 -1124 -4304
rect -1090 -4312 -1009 -4296
rect -858 -4304 -824 -4262
rect -1338 -4372 -1304 -4364
rect -1056 -4346 -1009 -4312
rect -1338 -4406 -1178 -4372
rect -1717 -4490 -1582 -4458
rect -1490 -4474 -1296 -4440
rect -1262 -4474 -1246 -4440
rect -1717 -4598 -1675 -4490
rect -1490 -4492 -1456 -4474
rect -1717 -4632 -1709 -4598
rect -1717 -4648 -1675 -4632
rect -1641 -4534 -1571 -4524
rect -1641 -4550 -1605 -4534
rect -1641 -4584 -1613 -4550
rect -1579 -4584 -1571 -4568
rect -1641 -4648 -1571 -4584
rect -1537 -4526 -1456 -4492
rect -1537 -4682 -1503 -4526
rect -1389 -4539 -1281 -4508
rect -1212 -4524 -1178 -4406
rect -1090 -4380 -1009 -4346
rect -1056 -4414 -1009 -4380
rect -1090 -4448 -1009 -4414
rect -1056 -4482 -1009 -4448
rect -1090 -4498 -1009 -4482
rect -1212 -4530 -1123 -4524
rect -1355 -4548 -1281 -4539
rect -1469 -4576 -1425 -4560
rect -1435 -4610 -1425 -4576
rect -1389 -4582 -1373 -4573
rect -1339 -4582 -1281 -4548
rect -1469 -4616 -1425 -4610
rect -1329 -4602 -1281 -4582
rect -1469 -4650 -1363 -4616
rect -1693 -4696 -1503 -4682
rect -1807 -4734 -1787 -4700
rect -1753 -4734 -1737 -4700
rect -1693 -4730 -1677 -4696
rect -1643 -4730 -1503 -4696
rect -1693 -4738 -1503 -4730
rect -1469 -4700 -1431 -4684
rect -1469 -4734 -1465 -4700
rect -1397 -4696 -1363 -4650
rect -1295 -4636 -1281 -4602
rect -1329 -4662 -1281 -4636
rect -1247 -4540 -1123 -4530
rect -1247 -4574 -1173 -4540
rect -1139 -4574 -1123 -4540
rect -1247 -4590 -1123 -4574
rect -1247 -4625 -1182 -4590
rect -1075 -4624 -1009 -4498
rect -1247 -4680 -1183 -4625
rect -1397 -4714 -1247 -4696
rect -1213 -4714 -1183 -4680
rect -1397 -4730 -1183 -4714
rect -1143 -4657 -1109 -4635
rect -1469 -4772 -1431 -4734
rect -1143 -4772 -1109 -4691
rect -1075 -4658 -1059 -4624
rect -1025 -4658 -1009 -4624
rect -1075 -4692 -1009 -4658
rect -1075 -4726 -1059 -4692
rect -1025 -4726 -1009 -4692
rect -971 -4338 -955 -4304
rect -921 -4338 -905 -4304
rect -971 -4372 -905 -4338
rect -971 -4406 -955 -4372
rect -921 -4406 -905 -4372
rect -971 -4524 -905 -4406
rect -676 -4312 -625 -4296
rect -858 -4372 -824 -4338
rect -858 -4440 -824 -4406
rect -858 -4490 -824 -4474
rect -774 -4340 -723 -4324
rect -740 -4374 -723 -4340
rect -774 -4408 -723 -4374
rect -740 -4442 -723 -4408
rect -676 -4346 -659 -4312
rect -676 -4380 -625 -4346
rect -591 -4328 -525 -4262
rect -591 -4362 -575 -4328
rect -541 -4362 -525 -4328
rect -491 -4312 -457 -4296
rect -676 -4414 -659 -4380
rect -491 -4380 -457 -4346
rect -625 -4414 -526 -4396
rect -676 -4430 -526 -4414
rect -774 -4464 -723 -4442
rect -774 -4500 -606 -4464
rect -765 -4515 -606 -4500
rect -971 -4540 -799 -4524
rect -971 -4574 -833 -4540
rect -971 -4590 -799 -4574
rect -765 -4549 -734 -4515
rect -696 -4540 -606 -4515
rect -696 -4549 -662 -4540
rect -765 -4574 -662 -4549
rect -628 -4574 -606 -4540
rect -971 -4670 -921 -4590
rect -765 -4594 -606 -4574
rect -572 -4525 -526 -4430
rect -572 -4534 -560 -4525
rect -538 -4568 -526 -4559
rect -765 -4630 -723 -4594
rect -572 -4628 -526 -4568
rect -774 -4646 -723 -4630
rect -971 -4704 -955 -4670
rect -971 -4720 -921 -4704
rect -858 -4676 -824 -4653
rect -1075 -4734 -1009 -4726
rect -858 -4772 -824 -4710
rect -740 -4680 -723 -4646
rect -774 -4736 -723 -4680
rect -676 -4662 -526 -4628
rect -676 -4670 -625 -4662
rect -676 -4704 -659 -4670
rect -491 -4670 -457 -4432
rect -423 -4456 -358 -4299
rect -324 -4304 -274 -4262
rect -324 -4338 -308 -4304
rect -324 -4354 -274 -4338
rect -240 -4312 -190 -4296
rect -240 -4346 -224 -4312
rect -240 -4362 -190 -4346
rect -147 -4306 -11 -4296
rect -147 -4340 -131 -4306
rect -97 -4340 -11 -4306
rect 104 -4314 170 -4262
rect 297 -4304 371 -4262
rect -147 -4362 -11 -4340
rect -240 -4388 -206 -4362
rect -285 -4422 -206 -4388
rect -172 -4398 -79 -4396
rect -411 -4479 -319 -4456
rect -411 -4513 -353 -4479
rect -411 -4614 -319 -4513
rect -411 -4648 -387 -4614
rect -349 -4648 -319 -4614
rect -411 -4666 -319 -4648
rect -676 -4720 -625 -4704
rect -591 -4730 -575 -4696
rect -541 -4730 -525 -4696
rect -285 -4694 -251 -4422
rect -172 -4424 -113 -4398
rect -138 -4432 -113 -4424
rect -138 -4458 -79 -4432
rect -172 -4474 -79 -4458
rect -217 -4534 -147 -4512
rect -217 -4568 -205 -4534
rect -171 -4568 -147 -4534
rect -217 -4586 -147 -4568
rect -217 -4620 -194 -4586
rect -160 -4620 -147 -4586
rect -217 -4636 -147 -4620
rect -113 -4592 -79 -4474
rect -45 -4518 -11 -4362
rect 23 -4330 57 -4314
rect 104 -4348 120 -4314
rect 154 -4348 170 -4314
rect 204 -4330 238 -4314
rect 23 -4382 57 -4364
rect 297 -4338 317 -4304
rect 351 -4338 371 -4304
rect 297 -4354 371 -4338
rect 405 -4312 439 -4296
rect 204 -4382 238 -4364
rect 23 -4416 238 -4382
rect 405 -4388 439 -4346
rect 486 -4305 660 -4296
rect 486 -4339 502 -4305
rect 536 -4339 660 -4305
rect 486 -4364 660 -4339
rect 694 -4304 744 -4262
rect 728 -4338 744 -4304
rect 848 -4304 992 -4262
rect 694 -4354 744 -4338
rect 778 -4330 812 -4314
rect 327 -4422 439 -4388
rect 327 -4450 361 -4422
rect 61 -4484 77 -4450
rect 111 -4484 361 -4450
rect 500 -4432 511 -4398
rect 545 -4424 592 -4398
rect 500 -4456 542 -4432
rect -45 -4538 293 -4518
rect -45 -4552 259 -4538
rect -113 -4626 -92 -4592
rect -58 -4626 -42 -4592
rect -113 -4636 -42 -4626
rect -8 -4694 26 -4552
rect 67 -4602 163 -4586
rect 101 -4636 139 -4602
rect 197 -4620 225 -4586
rect 259 -4588 293 -4572
rect 173 -4636 225 -4620
rect 327 -4622 361 -4484
rect -491 -4720 -457 -4704
rect -591 -4772 -525 -4730
rect -385 -4734 -369 -4700
rect -335 -4734 -319 -4700
rect -285 -4728 -236 -4694
rect -202 -4728 -186 -4694
rect -145 -4728 -129 -4694
rect -95 -4728 26 -4694
rect 201 -4696 267 -4680
rect -385 -4772 -319 -4734
rect 201 -4730 217 -4696
rect 251 -4730 267 -4696
rect 201 -4772 267 -4730
rect 309 -4700 361 -4622
rect 399 -4458 542 -4456
rect 576 -4458 592 -4424
rect 626 -4440 660 -4364
rect 848 -4338 864 -4304
rect 898 -4338 942 -4304
rect 976 -4338 992 -4304
rect 1026 -4312 1107 -4296
rect 1258 -4304 1292 -4262
rect 778 -4372 812 -4364
rect 1060 -4346 1107 -4312
rect 778 -4406 938 -4372
rect 399 -4490 534 -4458
rect 626 -4474 820 -4440
rect 854 -4474 870 -4440
rect 399 -4598 441 -4490
rect 626 -4492 660 -4474
rect 399 -4632 407 -4598
rect 399 -4648 441 -4632
rect 475 -4534 545 -4524
rect 475 -4550 511 -4534
rect 475 -4584 503 -4550
rect 537 -4584 545 -4568
rect 475 -4648 545 -4584
rect 579 -4526 660 -4492
rect 579 -4682 613 -4526
rect 727 -4539 835 -4508
rect 904 -4524 938 -4406
rect 1026 -4380 1107 -4346
rect 1060 -4414 1107 -4380
rect 1026 -4448 1107 -4414
rect 1060 -4482 1107 -4448
rect 1026 -4498 1107 -4482
rect 904 -4530 993 -4524
rect 761 -4548 835 -4539
rect 647 -4576 691 -4560
rect 681 -4610 691 -4576
rect 727 -4582 743 -4573
rect 777 -4582 835 -4548
rect 647 -4616 691 -4610
rect 787 -4602 835 -4582
rect 647 -4650 753 -4616
rect 423 -4696 613 -4682
rect 309 -4734 329 -4700
rect 363 -4734 379 -4700
rect 423 -4730 439 -4696
rect 473 -4730 613 -4696
rect 423 -4738 613 -4730
rect 647 -4700 685 -4684
rect 647 -4734 651 -4700
rect 719 -4696 753 -4650
rect 821 -4636 835 -4602
rect 787 -4662 835 -4636
rect 869 -4540 993 -4530
rect 869 -4574 943 -4540
rect 977 -4574 993 -4540
rect 869 -4590 993 -4574
rect 869 -4625 934 -4590
rect 1041 -4624 1107 -4498
rect 869 -4680 933 -4625
rect 719 -4714 869 -4696
rect 903 -4714 933 -4680
rect 719 -4730 933 -4714
rect 973 -4657 1007 -4635
rect 647 -4772 685 -4734
rect 973 -4772 1007 -4691
rect 1041 -4658 1057 -4624
rect 1091 -4658 1107 -4624
rect 1041 -4692 1107 -4658
rect 1041 -4726 1057 -4692
rect 1091 -4726 1107 -4692
rect 1145 -4338 1161 -4304
rect 1195 -4338 1211 -4304
rect 1145 -4372 1211 -4338
rect 1145 -4406 1161 -4372
rect 1195 -4406 1211 -4372
rect 1145 -4524 1211 -4406
rect 1440 -4312 1491 -4296
rect 1258 -4372 1292 -4338
rect 1258 -4440 1292 -4406
rect 1258 -4490 1292 -4474
rect 1342 -4340 1393 -4324
rect 1376 -4374 1393 -4340
rect 1342 -4408 1393 -4374
rect 1376 -4442 1393 -4408
rect 1440 -4346 1457 -4312
rect 1440 -4380 1491 -4346
rect 1525 -4328 1591 -4262
rect 1525 -4362 1541 -4328
rect 1575 -4362 1591 -4328
rect 1625 -4312 1659 -4296
rect 1440 -4414 1457 -4380
rect 1625 -4380 1659 -4346
rect 1491 -4414 1590 -4396
rect 1440 -4430 1590 -4414
rect 1342 -4464 1393 -4442
rect 1342 -4500 1510 -4464
rect 1351 -4515 1510 -4500
rect 1145 -4540 1317 -4524
rect 1145 -4574 1283 -4540
rect 1145 -4590 1317 -4574
rect 1351 -4549 1382 -4515
rect 1420 -4540 1510 -4515
rect 1420 -4549 1454 -4540
rect 1351 -4574 1454 -4549
rect 1488 -4574 1510 -4540
rect 1145 -4670 1195 -4590
rect 1351 -4594 1510 -4574
rect 1544 -4525 1590 -4430
rect 1544 -4534 1556 -4525
rect 1578 -4568 1590 -4559
rect 1351 -4630 1393 -4594
rect 1544 -4628 1590 -4568
rect 1342 -4646 1393 -4630
rect 1145 -4704 1161 -4670
rect 1145 -4720 1195 -4704
rect 1258 -4676 1292 -4653
rect 1041 -4734 1107 -4726
rect 1258 -4772 1292 -4710
rect 1376 -4680 1393 -4646
rect 1342 -4736 1393 -4680
rect 1440 -4662 1590 -4628
rect 1440 -4670 1491 -4662
rect 1440 -4704 1457 -4670
rect 1625 -4670 1659 -4432
rect 1693 -4456 1758 -4299
rect 1792 -4304 1842 -4262
rect 1792 -4338 1808 -4304
rect 1792 -4354 1842 -4338
rect 1876 -4312 1926 -4296
rect 1876 -4346 1892 -4312
rect 1876 -4362 1926 -4346
rect 1969 -4306 2105 -4296
rect 1969 -4340 1985 -4306
rect 2019 -4340 2105 -4306
rect 2220 -4314 2286 -4262
rect 2413 -4304 2487 -4262
rect 1969 -4362 2105 -4340
rect 1876 -4388 1910 -4362
rect 1831 -4422 1910 -4388
rect 1944 -4398 2037 -4396
rect 1705 -4479 1797 -4456
rect 1705 -4513 1763 -4479
rect 1705 -4614 1797 -4513
rect 1705 -4648 1729 -4614
rect 1767 -4648 1797 -4614
rect 1705 -4666 1797 -4648
rect 1440 -4720 1491 -4704
rect 1525 -4730 1541 -4696
rect 1575 -4730 1591 -4696
rect 1831 -4694 1865 -4422
rect 1944 -4424 2003 -4398
rect 1978 -4432 2003 -4424
rect 1978 -4458 2037 -4432
rect 1944 -4474 2037 -4458
rect 1899 -4534 1969 -4512
rect 1899 -4568 1911 -4534
rect 1945 -4568 1969 -4534
rect 1899 -4586 1969 -4568
rect 1899 -4620 1922 -4586
rect 1956 -4620 1969 -4586
rect 1899 -4636 1969 -4620
rect 2003 -4592 2037 -4474
rect 2071 -4518 2105 -4362
rect 2139 -4330 2173 -4314
rect 2220 -4348 2236 -4314
rect 2270 -4348 2286 -4314
rect 2320 -4330 2354 -4314
rect 2139 -4382 2173 -4364
rect 2413 -4338 2433 -4304
rect 2467 -4338 2487 -4304
rect 2413 -4354 2487 -4338
rect 2521 -4312 2555 -4296
rect 2320 -4382 2354 -4364
rect 2139 -4416 2354 -4382
rect 2521 -4388 2555 -4346
rect 2602 -4305 2776 -4296
rect 2602 -4339 2618 -4305
rect 2652 -4339 2776 -4305
rect 2602 -4364 2776 -4339
rect 2810 -4304 2860 -4262
rect 2844 -4338 2860 -4304
rect 2964 -4304 3108 -4262
rect 2810 -4354 2860 -4338
rect 2894 -4330 2928 -4314
rect 2443 -4422 2555 -4388
rect 2443 -4450 2477 -4422
rect 2177 -4484 2193 -4450
rect 2227 -4484 2477 -4450
rect 2616 -4432 2627 -4398
rect 2661 -4424 2708 -4398
rect 2616 -4456 2658 -4432
rect 2071 -4538 2409 -4518
rect 2071 -4552 2375 -4538
rect 2003 -4626 2024 -4592
rect 2058 -4626 2074 -4592
rect 2003 -4636 2074 -4626
rect 2108 -4694 2142 -4552
rect 2183 -4602 2279 -4586
rect 2217 -4636 2255 -4602
rect 2313 -4620 2341 -4586
rect 2375 -4588 2409 -4572
rect 2289 -4636 2341 -4620
rect 2443 -4622 2477 -4484
rect 1625 -4720 1659 -4704
rect 1525 -4772 1591 -4730
rect 1731 -4734 1747 -4700
rect 1781 -4734 1797 -4700
rect 1831 -4728 1880 -4694
rect 1914 -4728 1930 -4694
rect 1971 -4728 1987 -4694
rect 2021 -4728 2142 -4694
rect 2317 -4696 2383 -4680
rect 1731 -4772 1797 -4734
rect 2317 -4730 2333 -4696
rect 2367 -4730 2383 -4696
rect 2317 -4772 2383 -4730
rect 2425 -4700 2477 -4622
rect 2515 -4458 2658 -4456
rect 2692 -4458 2708 -4424
rect 2742 -4440 2776 -4364
rect 2964 -4338 2980 -4304
rect 3014 -4338 3058 -4304
rect 3092 -4338 3108 -4304
rect 3142 -4312 3223 -4296
rect 3374 -4304 3408 -4262
rect 2894 -4372 2928 -4364
rect 3176 -4346 3223 -4312
rect 2894 -4406 3054 -4372
rect 2515 -4490 2650 -4458
rect 2742 -4474 2936 -4440
rect 2970 -4474 2986 -4440
rect 2515 -4598 2557 -4490
rect 2742 -4492 2776 -4474
rect 2515 -4632 2523 -4598
rect 2515 -4648 2557 -4632
rect 2591 -4534 2661 -4524
rect 2591 -4550 2627 -4534
rect 2591 -4584 2619 -4550
rect 2653 -4584 2661 -4568
rect 2591 -4648 2661 -4584
rect 2695 -4526 2776 -4492
rect 2695 -4682 2729 -4526
rect 2843 -4539 2951 -4508
rect 3020 -4524 3054 -4406
rect 3142 -4380 3223 -4346
rect 3176 -4414 3223 -4380
rect 3142 -4448 3223 -4414
rect 3176 -4482 3223 -4448
rect 3142 -4498 3223 -4482
rect 3020 -4530 3109 -4524
rect 2877 -4548 2951 -4539
rect 2763 -4576 2807 -4560
rect 2797 -4610 2807 -4576
rect 2843 -4582 2859 -4573
rect 2893 -4582 2951 -4548
rect 2763 -4616 2807 -4610
rect 2903 -4602 2951 -4582
rect 2763 -4650 2869 -4616
rect 2539 -4696 2729 -4682
rect 2425 -4734 2445 -4700
rect 2479 -4734 2495 -4700
rect 2539 -4730 2555 -4696
rect 2589 -4730 2729 -4696
rect 2539 -4738 2729 -4730
rect 2763 -4700 2801 -4684
rect 2763 -4734 2767 -4700
rect 2835 -4696 2869 -4650
rect 2937 -4636 2951 -4602
rect 2903 -4662 2951 -4636
rect 2985 -4540 3109 -4530
rect 2985 -4574 3059 -4540
rect 3093 -4574 3109 -4540
rect 2985 -4590 3109 -4574
rect 2985 -4625 3050 -4590
rect 3157 -4624 3223 -4498
rect 2985 -4680 3049 -4625
rect 2835 -4714 2985 -4696
rect 3019 -4714 3049 -4680
rect 2835 -4730 3049 -4714
rect 3089 -4657 3123 -4635
rect 2763 -4772 2801 -4734
rect 3089 -4772 3123 -4691
rect 3157 -4658 3173 -4624
rect 3207 -4658 3223 -4624
rect 3157 -4692 3223 -4658
rect 3157 -4726 3173 -4692
rect 3207 -4726 3223 -4692
rect 3261 -4338 3277 -4304
rect 3311 -4338 3327 -4304
rect 3261 -4372 3327 -4338
rect 3261 -4406 3277 -4372
rect 3311 -4406 3327 -4372
rect 3261 -4524 3327 -4406
rect 3556 -4312 3607 -4296
rect 3374 -4372 3408 -4338
rect 3374 -4440 3408 -4406
rect 3374 -4490 3408 -4474
rect 3458 -4340 3509 -4324
rect 3492 -4374 3509 -4340
rect 3458 -4408 3509 -4374
rect 3492 -4442 3509 -4408
rect 3556 -4346 3573 -4312
rect 3556 -4380 3607 -4346
rect 3641 -4328 3707 -4262
rect 3641 -4362 3657 -4328
rect 3691 -4362 3707 -4328
rect 3741 -4312 3775 -4296
rect 3556 -4414 3573 -4380
rect 3741 -4380 3775 -4346
rect 3607 -4414 3706 -4396
rect 3556 -4430 3706 -4414
rect 3458 -4464 3509 -4442
rect 3458 -4500 3626 -4464
rect 3467 -4515 3626 -4500
rect 3261 -4540 3433 -4524
rect 3261 -4574 3399 -4540
rect 3261 -4590 3433 -4574
rect 3467 -4549 3498 -4515
rect 3536 -4540 3626 -4515
rect 3536 -4549 3570 -4540
rect 3467 -4574 3570 -4549
rect 3604 -4574 3626 -4540
rect 3261 -4670 3311 -4590
rect 3467 -4594 3626 -4574
rect 3660 -4525 3706 -4430
rect 3660 -4534 3672 -4525
rect 3694 -4568 3706 -4559
rect 3467 -4630 3509 -4594
rect 3660 -4628 3706 -4568
rect 3458 -4646 3509 -4630
rect 3261 -4704 3277 -4670
rect 3261 -4720 3311 -4704
rect 3374 -4676 3408 -4653
rect 3157 -4734 3223 -4726
rect 3374 -4772 3408 -4710
rect 3492 -4680 3509 -4646
rect 3458 -4736 3509 -4680
rect 3556 -4662 3706 -4628
rect 3556 -4670 3607 -4662
rect 3556 -4704 3573 -4670
rect 3741 -4670 3775 -4432
rect 3809 -4456 3874 -4299
rect 3908 -4304 3958 -4262
rect 3908 -4338 3924 -4304
rect 3908 -4354 3958 -4338
rect 3992 -4312 4042 -4296
rect 3992 -4346 4008 -4312
rect 3992 -4362 4042 -4346
rect 4085 -4306 4221 -4296
rect 4085 -4340 4101 -4306
rect 4135 -4340 4221 -4306
rect 4336 -4314 4402 -4262
rect 4529 -4304 4603 -4262
rect 4085 -4362 4221 -4340
rect 3992 -4388 4026 -4362
rect 3947 -4422 4026 -4388
rect 4060 -4398 4153 -4396
rect 3821 -4479 3913 -4456
rect 3821 -4513 3879 -4479
rect 3821 -4614 3913 -4513
rect 3821 -4648 3845 -4614
rect 3883 -4648 3913 -4614
rect 3821 -4666 3913 -4648
rect 3556 -4720 3607 -4704
rect 3641 -4730 3657 -4696
rect 3691 -4730 3707 -4696
rect 3947 -4694 3981 -4422
rect 4060 -4424 4119 -4398
rect 4094 -4432 4119 -4424
rect 4094 -4458 4153 -4432
rect 4060 -4474 4153 -4458
rect 4015 -4534 4085 -4512
rect 4015 -4568 4027 -4534
rect 4061 -4568 4085 -4534
rect 4015 -4586 4085 -4568
rect 4015 -4620 4038 -4586
rect 4072 -4620 4085 -4586
rect 4015 -4636 4085 -4620
rect 4119 -4592 4153 -4474
rect 4187 -4518 4221 -4362
rect 4255 -4330 4289 -4314
rect 4336 -4348 4352 -4314
rect 4386 -4348 4402 -4314
rect 4436 -4330 4470 -4314
rect 4255 -4382 4289 -4364
rect 4529 -4338 4549 -4304
rect 4583 -4338 4603 -4304
rect 4529 -4354 4603 -4338
rect 4637 -4312 4671 -4296
rect 4436 -4382 4470 -4364
rect 4255 -4416 4470 -4382
rect 4637 -4388 4671 -4346
rect 4718 -4305 4892 -4296
rect 4718 -4339 4734 -4305
rect 4768 -4339 4892 -4305
rect 4718 -4364 4892 -4339
rect 4926 -4304 4976 -4262
rect 4960 -4338 4976 -4304
rect 5080 -4304 5224 -4262
rect 4926 -4354 4976 -4338
rect 5010 -4330 5044 -4314
rect 4559 -4422 4671 -4388
rect 4559 -4450 4593 -4422
rect 4293 -4484 4309 -4450
rect 4343 -4484 4593 -4450
rect 4732 -4432 4743 -4398
rect 4777 -4424 4824 -4398
rect 4732 -4456 4774 -4432
rect 4187 -4538 4525 -4518
rect 4187 -4552 4491 -4538
rect 4119 -4626 4140 -4592
rect 4174 -4626 4190 -4592
rect 4119 -4636 4190 -4626
rect 4224 -4694 4258 -4552
rect 4299 -4602 4395 -4586
rect 4333 -4636 4371 -4602
rect 4429 -4620 4457 -4586
rect 4491 -4588 4525 -4572
rect 4405 -4636 4457 -4620
rect 4559 -4622 4593 -4484
rect 3741 -4720 3775 -4704
rect 3641 -4772 3707 -4730
rect 3847 -4734 3863 -4700
rect 3897 -4734 3913 -4700
rect 3947 -4728 3996 -4694
rect 4030 -4728 4046 -4694
rect 4087 -4728 4103 -4694
rect 4137 -4728 4258 -4694
rect 4433 -4696 4499 -4680
rect 3847 -4772 3913 -4734
rect 4433 -4730 4449 -4696
rect 4483 -4730 4499 -4696
rect 4433 -4772 4499 -4730
rect 4541 -4700 4593 -4622
rect 4631 -4458 4774 -4456
rect 4808 -4458 4824 -4424
rect 4858 -4440 4892 -4364
rect 5080 -4338 5096 -4304
rect 5130 -4338 5174 -4304
rect 5208 -4338 5224 -4304
rect 5258 -4312 5339 -4296
rect 5490 -4304 5524 -4262
rect 5010 -4372 5044 -4364
rect 5292 -4346 5339 -4312
rect 5010 -4406 5170 -4372
rect 4631 -4490 4766 -4458
rect 4858 -4474 5052 -4440
rect 5086 -4474 5102 -4440
rect 4631 -4598 4673 -4490
rect 4858 -4492 4892 -4474
rect 4631 -4632 4639 -4598
rect 4631 -4648 4673 -4632
rect 4707 -4534 4777 -4524
rect 4707 -4550 4743 -4534
rect 4707 -4584 4735 -4550
rect 4769 -4584 4777 -4568
rect 4707 -4648 4777 -4584
rect 4811 -4526 4892 -4492
rect 4811 -4682 4845 -4526
rect 4959 -4539 5067 -4508
rect 5136 -4524 5170 -4406
rect 5258 -4380 5339 -4346
rect 5292 -4414 5339 -4380
rect 5258 -4448 5339 -4414
rect 5292 -4482 5339 -4448
rect 5258 -4498 5339 -4482
rect 5136 -4530 5225 -4524
rect 4993 -4548 5067 -4539
rect 4879 -4576 4923 -4560
rect 4913 -4610 4923 -4576
rect 4959 -4582 4975 -4573
rect 5009 -4582 5067 -4548
rect 4879 -4616 4923 -4610
rect 5019 -4602 5067 -4582
rect 4879 -4650 4985 -4616
rect 4655 -4696 4845 -4682
rect 4541 -4734 4561 -4700
rect 4595 -4734 4611 -4700
rect 4655 -4730 4671 -4696
rect 4705 -4730 4845 -4696
rect 4655 -4738 4845 -4730
rect 4879 -4700 4917 -4684
rect 4879 -4734 4883 -4700
rect 4951 -4696 4985 -4650
rect 5053 -4636 5067 -4602
rect 5019 -4662 5067 -4636
rect 5101 -4540 5225 -4530
rect 5101 -4574 5175 -4540
rect 5209 -4574 5225 -4540
rect 5101 -4590 5225 -4574
rect 5101 -4625 5166 -4590
rect 5273 -4624 5339 -4498
rect 5101 -4680 5165 -4625
rect 4951 -4714 5101 -4696
rect 5135 -4714 5165 -4680
rect 4951 -4730 5165 -4714
rect 5205 -4657 5239 -4635
rect 4879 -4772 4917 -4734
rect 5205 -4772 5239 -4691
rect 5273 -4658 5289 -4624
rect 5323 -4658 5339 -4624
rect 5273 -4692 5339 -4658
rect 5273 -4726 5289 -4692
rect 5323 -4726 5339 -4692
rect 5377 -4338 5393 -4304
rect 5427 -4338 5443 -4304
rect 5377 -4372 5443 -4338
rect 5377 -4406 5393 -4372
rect 5427 -4406 5443 -4372
rect 5377 -4524 5443 -4406
rect 5672 -4312 5723 -4296
rect 5490 -4372 5524 -4338
rect 5490 -4440 5524 -4406
rect 5490 -4490 5524 -4474
rect 5574 -4340 5625 -4324
rect 5608 -4374 5625 -4340
rect 5574 -4408 5625 -4374
rect 5608 -4442 5625 -4408
rect 5672 -4346 5689 -4312
rect 5672 -4380 5723 -4346
rect 5757 -4328 5823 -4262
rect 5757 -4362 5773 -4328
rect 5807 -4362 5823 -4328
rect 5857 -4312 5891 -4296
rect 5672 -4414 5689 -4380
rect 5857 -4380 5891 -4346
rect 5723 -4414 5822 -4396
rect 5672 -4430 5822 -4414
rect 5574 -4464 5625 -4442
rect 5574 -4500 5742 -4464
rect 5583 -4515 5742 -4500
rect 5377 -4540 5549 -4524
rect 5377 -4574 5515 -4540
rect 5377 -4590 5549 -4574
rect 5583 -4549 5614 -4515
rect 5652 -4540 5742 -4515
rect 5652 -4549 5686 -4540
rect 5583 -4574 5686 -4549
rect 5720 -4574 5742 -4540
rect 5377 -4670 5427 -4590
rect 5583 -4594 5742 -4574
rect 5776 -4525 5822 -4430
rect 5776 -4534 5788 -4525
rect 5810 -4568 5822 -4559
rect 5583 -4630 5625 -4594
rect 5776 -4628 5822 -4568
rect 5574 -4646 5625 -4630
rect 5377 -4704 5393 -4670
rect 5377 -4720 5427 -4704
rect 5490 -4676 5524 -4653
rect 5273 -4734 5339 -4726
rect 5490 -4772 5524 -4710
rect 5608 -4680 5625 -4646
rect 5574 -4736 5625 -4680
rect 5672 -4662 5822 -4628
rect 5672 -4670 5723 -4662
rect 5672 -4704 5689 -4670
rect 5857 -4670 5891 -4432
rect 5925 -4456 5990 -4299
rect 6024 -4304 6074 -4262
rect 6024 -4338 6040 -4304
rect 6024 -4354 6074 -4338
rect 6108 -4312 6158 -4296
rect 6108 -4346 6124 -4312
rect 6108 -4362 6158 -4346
rect 6201 -4306 6337 -4296
rect 6201 -4340 6217 -4306
rect 6251 -4340 6337 -4306
rect 6452 -4314 6518 -4262
rect 6645 -4304 6719 -4262
rect 6201 -4362 6337 -4340
rect 6108 -4388 6142 -4362
rect 6063 -4422 6142 -4388
rect 6176 -4398 6269 -4396
rect 5937 -4479 6029 -4456
rect 5937 -4513 5995 -4479
rect 5937 -4614 6029 -4513
rect 5937 -4648 5961 -4614
rect 5999 -4648 6029 -4614
rect 5937 -4666 6029 -4648
rect 5672 -4720 5723 -4704
rect 5757 -4730 5773 -4696
rect 5807 -4730 5823 -4696
rect 6063 -4694 6097 -4422
rect 6176 -4424 6235 -4398
rect 6210 -4432 6235 -4424
rect 6210 -4458 6269 -4432
rect 6176 -4474 6269 -4458
rect 6131 -4534 6201 -4512
rect 6131 -4568 6143 -4534
rect 6177 -4568 6201 -4534
rect 6131 -4586 6201 -4568
rect 6131 -4620 6154 -4586
rect 6188 -4620 6201 -4586
rect 6131 -4636 6201 -4620
rect 6235 -4592 6269 -4474
rect 6303 -4518 6337 -4362
rect 6371 -4330 6405 -4314
rect 6452 -4348 6468 -4314
rect 6502 -4348 6518 -4314
rect 6552 -4330 6586 -4314
rect 6371 -4382 6405 -4364
rect 6645 -4338 6665 -4304
rect 6699 -4338 6719 -4304
rect 6645 -4354 6719 -4338
rect 6753 -4312 6787 -4296
rect 6552 -4382 6586 -4364
rect 6371 -4416 6586 -4382
rect 6753 -4388 6787 -4346
rect 6834 -4305 7008 -4296
rect 6834 -4339 6850 -4305
rect 6884 -4339 7008 -4305
rect 6834 -4364 7008 -4339
rect 7042 -4304 7092 -4262
rect 7076 -4338 7092 -4304
rect 7196 -4304 7340 -4262
rect 7042 -4354 7092 -4338
rect 7126 -4330 7160 -4314
rect 6675 -4422 6787 -4388
rect 6675 -4450 6709 -4422
rect 6409 -4484 6425 -4450
rect 6459 -4484 6709 -4450
rect 6848 -4432 6859 -4398
rect 6893 -4424 6940 -4398
rect 6848 -4456 6890 -4432
rect 6303 -4538 6641 -4518
rect 6303 -4552 6607 -4538
rect 6235 -4626 6256 -4592
rect 6290 -4626 6306 -4592
rect 6235 -4636 6306 -4626
rect 6340 -4694 6374 -4552
rect 6415 -4602 6511 -4586
rect 6449 -4636 6487 -4602
rect 6545 -4620 6573 -4586
rect 6607 -4588 6641 -4572
rect 6521 -4636 6573 -4620
rect 6675 -4622 6709 -4484
rect 5857 -4720 5891 -4704
rect 5757 -4772 5823 -4730
rect 5963 -4734 5979 -4700
rect 6013 -4734 6029 -4700
rect 6063 -4728 6112 -4694
rect 6146 -4728 6162 -4694
rect 6203 -4728 6219 -4694
rect 6253 -4728 6374 -4694
rect 6549 -4696 6615 -4680
rect 5963 -4772 6029 -4734
rect 6549 -4730 6565 -4696
rect 6599 -4730 6615 -4696
rect 6549 -4772 6615 -4730
rect 6657 -4700 6709 -4622
rect 6747 -4458 6890 -4456
rect 6924 -4458 6940 -4424
rect 6974 -4440 7008 -4364
rect 7196 -4338 7212 -4304
rect 7246 -4338 7290 -4304
rect 7324 -4338 7340 -4304
rect 7374 -4312 7455 -4296
rect 7606 -4304 7640 -4262
rect 7126 -4372 7160 -4364
rect 7408 -4346 7455 -4312
rect 7126 -4406 7286 -4372
rect 6747 -4490 6882 -4458
rect 6974 -4474 7168 -4440
rect 7202 -4474 7218 -4440
rect 6747 -4598 6789 -4490
rect 6974 -4492 7008 -4474
rect 6747 -4632 6755 -4598
rect 6747 -4648 6789 -4632
rect 6823 -4534 6893 -4524
rect 6823 -4550 6859 -4534
rect 6823 -4584 6851 -4550
rect 6885 -4584 6893 -4568
rect 6823 -4648 6893 -4584
rect 6927 -4526 7008 -4492
rect 6927 -4682 6961 -4526
rect 7075 -4539 7183 -4508
rect 7252 -4524 7286 -4406
rect 7374 -4380 7455 -4346
rect 7408 -4414 7455 -4380
rect 7374 -4448 7455 -4414
rect 7408 -4482 7455 -4448
rect 7374 -4498 7455 -4482
rect 7252 -4530 7341 -4524
rect 7109 -4548 7183 -4539
rect 6995 -4576 7039 -4560
rect 7029 -4610 7039 -4576
rect 7075 -4582 7091 -4573
rect 7125 -4582 7183 -4548
rect 6995 -4616 7039 -4610
rect 7135 -4602 7183 -4582
rect 6995 -4650 7101 -4616
rect 6771 -4696 6961 -4682
rect 6657 -4734 6677 -4700
rect 6711 -4734 6727 -4700
rect 6771 -4730 6787 -4696
rect 6821 -4730 6961 -4696
rect 6771 -4738 6961 -4730
rect 6995 -4700 7033 -4684
rect 6995 -4734 6999 -4700
rect 7067 -4696 7101 -4650
rect 7169 -4636 7183 -4602
rect 7135 -4662 7183 -4636
rect 7217 -4540 7341 -4530
rect 7217 -4574 7291 -4540
rect 7325 -4574 7341 -4540
rect 7217 -4590 7341 -4574
rect 7217 -4625 7282 -4590
rect 7389 -4624 7455 -4498
rect 7217 -4680 7281 -4625
rect 7067 -4714 7217 -4696
rect 7251 -4714 7281 -4680
rect 7067 -4730 7281 -4714
rect 7321 -4657 7355 -4635
rect 6995 -4772 7033 -4734
rect 7321 -4772 7355 -4691
rect 7389 -4658 7405 -4624
rect 7439 -4658 7455 -4624
rect 7389 -4692 7455 -4658
rect 7389 -4726 7405 -4692
rect 7439 -4726 7455 -4692
rect 7493 -4338 7509 -4304
rect 7543 -4338 7559 -4304
rect 7493 -4372 7559 -4338
rect 7493 -4406 7509 -4372
rect 7543 -4406 7559 -4372
rect 7493 -4524 7559 -4406
rect 7788 -4312 7839 -4296
rect 7606 -4372 7640 -4338
rect 7606 -4440 7640 -4406
rect 7606 -4490 7640 -4474
rect 7690 -4340 7741 -4324
rect 7724 -4374 7741 -4340
rect 7690 -4408 7741 -4374
rect 7724 -4442 7741 -4408
rect 7788 -4346 7805 -4312
rect 7788 -4380 7839 -4346
rect 7873 -4328 7939 -4262
rect 7873 -4362 7889 -4328
rect 7923 -4362 7939 -4328
rect 7973 -4312 8007 -4296
rect 7788 -4414 7805 -4380
rect 7973 -4380 8007 -4346
rect 7839 -4414 7938 -4396
rect 7788 -4430 7938 -4414
rect 7690 -4464 7741 -4442
rect 7690 -4500 7858 -4464
rect 7699 -4515 7858 -4500
rect 7493 -4540 7665 -4524
rect 7493 -4574 7631 -4540
rect 7493 -4590 7665 -4574
rect 7699 -4549 7730 -4515
rect 7768 -4540 7858 -4515
rect 7768 -4549 7802 -4540
rect 7699 -4574 7802 -4549
rect 7836 -4574 7858 -4540
rect 7493 -4670 7543 -4590
rect 7699 -4594 7858 -4574
rect 7892 -4525 7938 -4430
rect 7892 -4534 7904 -4525
rect 7926 -4568 7938 -4559
rect 7699 -4630 7741 -4594
rect 7892 -4628 7938 -4568
rect 7690 -4646 7741 -4630
rect 7493 -4704 7509 -4670
rect 7493 -4720 7543 -4704
rect 7606 -4676 7640 -4653
rect 7389 -4734 7455 -4726
rect 7606 -4772 7640 -4710
rect 7724 -4680 7741 -4646
rect 7690 -4736 7741 -4680
rect 7788 -4662 7938 -4628
rect 7788 -4670 7839 -4662
rect 7788 -4704 7805 -4670
rect 7973 -4670 8007 -4432
rect 8041 -4456 8106 -4299
rect 8140 -4304 8190 -4262
rect 8140 -4338 8156 -4304
rect 8140 -4354 8190 -4338
rect 8224 -4312 8274 -4296
rect 8224 -4346 8240 -4312
rect 8224 -4362 8274 -4346
rect 8317 -4306 8453 -4296
rect 8317 -4340 8333 -4306
rect 8367 -4340 8453 -4306
rect 8568 -4314 8634 -4262
rect 8761 -4304 8835 -4262
rect 8317 -4362 8453 -4340
rect 8224 -4388 8258 -4362
rect 8179 -4422 8258 -4388
rect 8292 -4398 8385 -4396
rect 8053 -4479 8145 -4456
rect 8053 -4513 8111 -4479
rect 8053 -4614 8145 -4513
rect 8053 -4648 8077 -4614
rect 8115 -4648 8145 -4614
rect 8053 -4666 8145 -4648
rect 7788 -4720 7839 -4704
rect 7873 -4730 7889 -4696
rect 7923 -4730 7939 -4696
rect 8179 -4694 8213 -4422
rect 8292 -4424 8351 -4398
rect 8326 -4432 8351 -4424
rect 8326 -4458 8385 -4432
rect 8292 -4474 8385 -4458
rect 8247 -4534 8317 -4512
rect 8247 -4568 8259 -4534
rect 8293 -4568 8317 -4534
rect 8247 -4586 8317 -4568
rect 8247 -4620 8270 -4586
rect 8304 -4620 8317 -4586
rect 8247 -4636 8317 -4620
rect 8351 -4592 8385 -4474
rect 8419 -4518 8453 -4362
rect 8487 -4330 8521 -4314
rect 8568 -4348 8584 -4314
rect 8618 -4348 8634 -4314
rect 8668 -4330 8702 -4314
rect 8487 -4382 8521 -4364
rect 8761 -4338 8781 -4304
rect 8815 -4338 8835 -4304
rect 8761 -4354 8835 -4338
rect 8869 -4312 8903 -4296
rect 8668 -4382 8702 -4364
rect 8487 -4416 8702 -4382
rect 8869 -4388 8903 -4346
rect 8950 -4305 9124 -4296
rect 8950 -4339 8966 -4305
rect 9000 -4339 9124 -4305
rect 8950 -4364 9124 -4339
rect 9158 -4304 9208 -4262
rect 9192 -4338 9208 -4304
rect 9312 -4304 9456 -4262
rect 9158 -4354 9208 -4338
rect 9242 -4330 9276 -4314
rect 8791 -4422 8903 -4388
rect 8791 -4450 8825 -4422
rect 8525 -4484 8541 -4450
rect 8575 -4484 8825 -4450
rect 8964 -4432 8975 -4398
rect 9009 -4424 9056 -4398
rect 8964 -4456 9006 -4432
rect 8419 -4538 8757 -4518
rect 8419 -4552 8723 -4538
rect 8351 -4626 8372 -4592
rect 8406 -4626 8422 -4592
rect 8351 -4636 8422 -4626
rect 8456 -4694 8490 -4552
rect 8531 -4602 8627 -4586
rect 8565 -4636 8603 -4602
rect 8661 -4620 8689 -4586
rect 8723 -4588 8757 -4572
rect 8637 -4636 8689 -4620
rect 8791 -4622 8825 -4484
rect 7973 -4720 8007 -4704
rect 7873 -4772 7939 -4730
rect 8079 -4734 8095 -4700
rect 8129 -4734 8145 -4700
rect 8179 -4728 8228 -4694
rect 8262 -4728 8278 -4694
rect 8319 -4728 8335 -4694
rect 8369 -4728 8490 -4694
rect 8665 -4696 8731 -4680
rect 8079 -4772 8145 -4734
rect 8665 -4730 8681 -4696
rect 8715 -4730 8731 -4696
rect 8665 -4772 8731 -4730
rect 8773 -4700 8825 -4622
rect 8863 -4458 9006 -4456
rect 9040 -4458 9056 -4424
rect 9090 -4440 9124 -4364
rect 9312 -4338 9328 -4304
rect 9362 -4338 9406 -4304
rect 9440 -4338 9456 -4304
rect 9490 -4312 9571 -4296
rect 9722 -4304 9756 -4262
rect 9242 -4372 9276 -4364
rect 9524 -4346 9571 -4312
rect 9242 -4406 9402 -4372
rect 8863 -4490 8998 -4458
rect 9090 -4474 9284 -4440
rect 9318 -4474 9334 -4440
rect 8863 -4598 8905 -4490
rect 9090 -4492 9124 -4474
rect 8863 -4632 8871 -4598
rect 8863 -4648 8905 -4632
rect 8939 -4534 9009 -4524
rect 8939 -4550 8975 -4534
rect 8939 -4584 8967 -4550
rect 9001 -4584 9009 -4568
rect 8939 -4648 9009 -4584
rect 9043 -4526 9124 -4492
rect 9043 -4682 9077 -4526
rect 9191 -4539 9299 -4508
rect 9368 -4524 9402 -4406
rect 9490 -4380 9571 -4346
rect 9524 -4414 9571 -4380
rect 9490 -4448 9571 -4414
rect 9524 -4482 9571 -4448
rect 9490 -4498 9571 -4482
rect 9368 -4530 9457 -4524
rect 9225 -4548 9299 -4539
rect 9111 -4576 9155 -4560
rect 9145 -4610 9155 -4576
rect 9191 -4582 9207 -4573
rect 9241 -4582 9299 -4548
rect 9111 -4616 9155 -4610
rect 9251 -4602 9299 -4582
rect 9111 -4650 9217 -4616
rect 8887 -4696 9077 -4682
rect 8773 -4734 8793 -4700
rect 8827 -4734 8843 -4700
rect 8887 -4730 8903 -4696
rect 8937 -4730 9077 -4696
rect 8887 -4738 9077 -4730
rect 9111 -4700 9149 -4684
rect 9111 -4734 9115 -4700
rect 9183 -4696 9217 -4650
rect 9285 -4636 9299 -4602
rect 9251 -4662 9299 -4636
rect 9333 -4540 9457 -4530
rect 9333 -4574 9407 -4540
rect 9441 -4574 9457 -4540
rect 9333 -4590 9457 -4574
rect 9333 -4625 9398 -4590
rect 9505 -4624 9571 -4498
rect 9333 -4680 9397 -4625
rect 9183 -4714 9333 -4696
rect 9367 -4714 9397 -4680
rect 9183 -4730 9397 -4714
rect 9437 -4657 9471 -4635
rect 9111 -4772 9149 -4734
rect 9437 -4772 9471 -4691
rect 9505 -4658 9521 -4624
rect 9555 -4658 9571 -4624
rect 9505 -4692 9571 -4658
rect 9505 -4726 9521 -4692
rect 9555 -4726 9571 -4692
rect 9609 -4338 9625 -4304
rect 9659 -4338 9675 -4304
rect 9609 -4372 9675 -4338
rect 9609 -4406 9625 -4372
rect 9659 -4406 9675 -4372
rect 9609 -4524 9675 -4406
rect 9904 -4312 9955 -4296
rect 9722 -4372 9756 -4338
rect 9722 -4440 9756 -4406
rect 9722 -4490 9756 -4474
rect 9806 -4340 9857 -4324
rect 9840 -4374 9857 -4340
rect 9806 -4408 9857 -4374
rect 9840 -4442 9857 -4408
rect 9904 -4346 9921 -4312
rect 9904 -4380 9955 -4346
rect 9989 -4328 10055 -4262
rect 9989 -4362 10005 -4328
rect 10039 -4362 10055 -4328
rect 10089 -4312 10123 -4296
rect 9904 -4414 9921 -4380
rect 10089 -4380 10123 -4346
rect 9955 -4414 10054 -4396
rect 9904 -4430 10054 -4414
rect 9806 -4464 9857 -4442
rect 9806 -4500 9974 -4464
rect 9815 -4515 9974 -4500
rect 9609 -4540 9781 -4524
rect 9609 -4574 9747 -4540
rect 9609 -4590 9781 -4574
rect 9815 -4549 9846 -4515
rect 9884 -4540 9974 -4515
rect 9884 -4549 9918 -4540
rect 9815 -4574 9918 -4549
rect 9952 -4574 9974 -4540
rect 9609 -4670 9659 -4590
rect 9815 -4594 9974 -4574
rect 10008 -4525 10054 -4430
rect 10008 -4534 10020 -4525
rect 10042 -4568 10054 -4559
rect 9815 -4630 9857 -4594
rect 10008 -4628 10054 -4568
rect 9806 -4646 9857 -4630
rect 9609 -4704 9625 -4670
rect 9609 -4720 9659 -4704
rect 9722 -4676 9756 -4653
rect 9505 -4734 9571 -4726
rect 9722 -4772 9756 -4710
rect 9840 -4680 9857 -4646
rect 9806 -4736 9857 -4680
rect 9904 -4662 10054 -4628
rect 9904 -4670 9955 -4662
rect 9904 -4704 9921 -4670
rect 10089 -4670 10123 -4432
rect 10157 -4456 10222 -4299
rect 10256 -4304 10306 -4262
rect 10256 -4338 10272 -4304
rect 10256 -4354 10306 -4338
rect 10340 -4312 10390 -4296
rect 10340 -4346 10356 -4312
rect 10340 -4362 10390 -4346
rect 10433 -4306 10569 -4296
rect 10433 -4340 10449 -4306
rect 10483 -4340 10569 -4306
rect 10684 -4314 10750 -4262
rect 10877 -4304 10951 -4262
rect 10433 -4362 10569 -4340
rect 10340 -4388 10374 -4362
rect 10295 -4422 10374 -4388
rect 10408 -4398 10501 -4396
rect 10169 -4479 10261 -4456
rect 10169 -4513 10227 -4479
rect 10169 -4614 10261 -4513
rect 10169 -4648 10193 -4614
rect 10231 -4648 10261 -4614
rect 10169 -4666 10261 -4648
rect 9904 -4720 9955 -4704
rect 9989 -4730 10005 -4696
rect 10039 -4730 10055 -4696
rect 10295 -4694 10329 -4422
rect 10408 -4424 10467 -4398
rect 10442 -4432 10467 -4424
rect 10442 -4458 10501 -4432
rect 10408 -4474 10501 -4458
rect 10363 -4534 10433 -4512
rect 10363 -4568 10375 -4534
rect 10409 -4568 10433 -4534
rect 10363 -4586 10433 -4568
rect 10363 -4620 10386 -4586
rect 10420 -4620 10433 -4586
rect 10363 -4636 10433 -4620
rect 10467 -4592 10501 -4474
rect 10535 -4518 10569 -4362
rect 10603 -4330 10637 -4314
rect 10684 -4348 10700 -4314
rect 10734 -4348 10750 -4314
rect 10784 -4330 10818 -4314
rect 10603 -4382 10637 -4364
rect 10877 -4338 10897 -4304
rect 10931 -4338 10951 -4304
rect 10877 -4354 10951 -4338
rect 10985 -4312 11019 -4296
rect 10784 -4382 10818 -4364
rect 10603 -4416 10818 -4382
rect 10985 -4388 11019 -4346
rect 11066 -4305 11240 -4296
rect 11066 -4339 11082 -4305
rect 11116 -4339 11240 -4305
rect 11066 -4364 11240 -4339
rect 11274 -4304 11324 -4262
rect 11308 -4338 11324 -4304
rect 11428 -4304 11572 -4262
rect 11274 -4354 11324 -4338
rect 11358 -4330 11392 -4314
rect 10907 -4422 11019 -4388
rect 10907 -4450 10941 -4422
rect 10641 -4484 10657 -4450
rect 10691 -4484 10941 -4450
rect 11080 -4432 11091 -4398
rect 11125 -4424 11172 -4398
rect 11080 -4456 11122 -4432
rect 10535 -4538 10873 -4518
rect 10535 -4552 10839 -4538
rect 10467 -4626 10488 -4592
rect 10522 -4626 10538 -4592
rect 10467 -4636 10538 -4626
rect 10572 -4694 10606 -4552
rect 10647 -4602 10743 -4586
rect 10681 -4636 10719 -4602
rect 10777 -4620 10805 -4586
rect 10839 -4588 10873 -4572
rect 10753 -4636 10805 -4620
rect 10907 -4622 10941 -4484
rect 10089 -4720 10123 -4704
rect 9989 -4772 10055 -4730
rect 10195 -4734 10211 -4700
rect 10245 -4734 10261 -4700
rect 10295 -4728 10344 -4694
rect 10378 -4728 10394 -4694
rect 10435 -4728 10451 -4694
rect 10485 -4728 10606 -4694
rect 10781 -4696 10847 -4680
rect 10195 -4772 10261 -4734
rect 10781 -4730 10797 -4696
rect 10831 -4730 10847 -4696
rect 10781 -4772 10847 -4730
rect 10889 -4700 10941 -4622
rect 10979 -4458 11122 -4456
rect 11156 -4458 11172 -4424
rect 11206 -4440 11240 -4364
rect 11428 -4338 11444 -4304
rect 11478 -4338 11522 -4304
rect 11556 -4338 11572 -4304
rect 11606 -4312 11687 -4296
rect 11838 -4304 11872 -4262
rect 11358 -4372 11392 -4364
rect 11640 -4346 11687 -4312
rect 11358 -4406 11518 -4372
rect 10979 -4490 11114 -4458
rect 11206 -4474 11400 -4440
rect 11434 -4474 11450 -4440
rect 10979 -4598 11021 -4490
rect 11206 -4492 11240 -4474
rect 10979 -4632 10987 -4598
rect 10979 -4648 11021 -4632
rect 11055 -4534 11125 -4524
rect 11055 -4550 11091 -4534
rect 11055 -4584 11083 -4550
rect 11117 -4584 11125 -4568
rect 11055 -4648 11125 -4584
rect 11159 -4526 11240 -4492
rect 11159 -4682 11193 -4526
rect 11307 -4539 11415 -4508
rect 11484 -4524 11518 -4406
rect 11606 -4380 11687 -4346
rect 11640 -4414 11687 -4380
rect 11606 -4448 11687 -4414
rect 11640 -4482 11687 -4448
rect 11606 -4498 11687 -4482
rect 11484 -4530 11573 -4524
rect 11341 -4548 11415 -4539
rect 11227 -4576 11271 -4560
rect 11261 -4610 11271 -4576
rect 11307 -4582 11323 -4573
rect 11357 -4582 11415 -4548
rect 11227 -4616 11271 -4610
rect 11367 -4602 11415 -4582
rect 11227 -4650 11333 -4616
rect 11003 -4696 11193 -4682
rect 10889 -4734 10909 -4700
rect 10943 -4734 10959 -4700
rect 11003 -4730 11019 -4696
rect 11053 -4730 11193 -4696
rect 11003 -4738 11193 -4730
rect 11227 -4700 11265 -4684
rect 11227 -4734 11231 -4700
rect 11299 -4696 11333 -4650
rect 11401 -4636 11415 -4602
rect 11367 -4662 11415 -4636
rect 11449 -4540 11573 -4530
rect 11449 -4574 11523 -4540
rect 11557 -4574 11573 -4540
rect 11449 -4590 11573 -4574
rect 11449 -4625 11514 -4590
rect 11621 -4624 11687 -4498
rect 11449 -4680 11513 -4625
rect 11299 -4714 11449 -4696
rect 11483 -4714 11513 -4680
rect 11299 -4730 11513 -4714
rect 11553 -4657 11587 -4635
rect 11227 -4772 11265 -4734
rect 11553 -4772 11587 -4691
rect 11621 -4658 11637 -4624
rect 11671 -4658 11687 -4624
rect 11621 -4692 11687 -4658
rect 11621 -4726 11637 -4692
rect 11671 -4726 11687 -4692
rect 11725 -4338 11741 -4304
rect 11775 -4338 11791 -4304
rect 11725 -4372 11791 -4338
rect 11725 -4406 11741 -4372
rect 11775 -4406 11791 -4372
rect 11725 -4524 11791 -4406
rect 12020 -4312 12071 -4296
rect 11838 -4372 11872 -4338
rect 11838 -4440 11872 -4406
rect 11838 -4490 11872 -4474
rect 11922 -4340 11973 -4324
rect 11956 -4374 11973 -4340
rect 11922 -4408 11973 -4374
rect 11956 -4442 11973 -4408
rect 12020 -4346 12037 -4312
rect 12020 -4380 12071 -4346
rect 12105 -4328 12171 -4262
rect 12105 -4362 12121 -4328
rect 12155 -4362 12171 -4328
rect 12205 -4312 12239 -4296
rect 12020 -4414 12037 -4380
rect 12205 -4380 12239 -4346
rect 12071 -4414 12170 -4396
rect 12020 -4430 12170 -4414
rect 11922 -4464 11973 -4442
rect 11922 -4500 12090 -4464
rect 11931 -4515 12090 -4500
rect 11725 -4540 11897 -4524
rect 11725 -4574 11863 -4540
rect 11725 -4590 11897 -4574
rect 11931 -4549 11962 -4515
rect 12000 -4540 12090 -4515
rect 12000 -4549 12034 -4540
rect 11931 -4574 12034 -4549
rect 12068 -4574 12090 -4540
rect 11725 -4670 11775 -4590
rect 11931 -4594 12090 -4574
rect 12124 -4525 12170 -4430
rect 12124 -4534 12136 -4525
rect 12158 -4568 12170 -4559
rect 11931 -4630 11973 -4594
rect 12124 -4628 12170 -4568
rect 11922 -4646 11973 -4630
rect 11725 -4704 11741 -4670
rect 11725 -4720 11775 -4704
rect 11838 -4676 11872 -4653
rect 11621 -4734 11687 -4726
rect 11838 -4772 11872 -4710
rect 11956 -4680 11973 -4646
rect 11922 -4736 11973 -4680
rect 12020 -4662 12170 -4628
rect 12020 -4670 12071 -4662
rect 12020 -4704 12037 -4670
rect 12205 -4670 12239 -4432
rect 12273 -4456 12338 -4299
rect 12372 -4304 12422 -4262
rect 12372 -4338 12388 -4304
rect 12372 -4354 12422 -4338
rect 12456 -4312 12506 -4296
rect 12456 -4346 12472 -4312
rect 12456 -4362 12506 -4346
rect 12549 -4306 12685 -4296
rect 12549 -4340 12565 -4306
rect 12599 -4340 12685 -4306
rect 12800 -4314 12866 -4262
rect 12993 -4304 13067 -4262
rect 12549 -4362 12685 -4340
rect 12456 -4388 12490 -4362
rect 12411 -4422 12490 -4388
rect 12524 -4398 12617 -4396
rect 12285 -4479 12377 -4456
rect 12285 -4513 12343 -4479
rect 12285 -4614 12377 -4513
rect 12285 -4648 12309 -4614
rect 12347 -4648 12377 -4614
rect 12285 -4666 12377 -4648
rect 12020 -4720 12071 -4704
rect 12105 -4730 12121 -4696
rect 12155 -4730 12171 -4696
rect 12411 -4694 12445 -4422
rect 12524 -4424 12583 -4398
rect 12558 -4432 12583 -4424
rect 12558 -4458 12617 -4432
rect 12524 -4474 12617 -4458
rect 12479 -4534 12549 -4512
rect 12479 -4568 12491 -4534
rect 12525 -4568 12549 -4534
rect 12479 -4586 12549 -4568
rect 12479 -4620 12502 -4586
rect 12536 -4620 12549 -4586
rect 12479 -4636 12549 -4620
rect 12583 -4592 12617 -4474
rect 12651 -4518 12685 -4362
rect 12719 -4330 12753 -4314
rect 12800 -4348 12816 -4314
rect 12850 -4348 12866 -4314
rect 12900 -4330 12934 -4314
rect 12719 -4382 12753 -4364
rect 12993 -4338 13013 -4304
rect 13047 -4338 13067 -4304
rect 12993 -4354 13067 -4338
rect 13101 -4312 13135 -4296
rect 12900 -4382 12934 -4364
rect 12719 -4416 12934 -4382
rect 13101 -4388 13135 -4346
rect 13182 -4305 13356 -4296
rect 13182 -4339 13198 -4305
rect 13232 -4339 13356 -4305
rect 13182 -4364 13356 -4339
rect 13390 -4304 13440 -4262
rect 13424 -4338 13440 -4304
rect 13544 -4304 13688 -4262
rect 13390 -4354 13440 -4338
rect 13474 -4330 13508 -4314
rect 13023 -4422 13135 -4388
rect 13023 -4450 13057 -4422
rect 12757 -4484 12773 -4450
rect 12807 -4484 13057 -4450
rect 13196 -4432 13207 -4398
rect 13241 -4424 13288 -4398
rect 13196 -4456 13238 -4432
rect 12651 -4538 12989 -4518
rect 12651 -4552 12955 -4538
rect 12583 -4626 12604 -4592
rect 12638 -4626 12654 -4592
rect 12583 -4636 12654 -4626
rect 12688 -4694 12722 -4552
rect 12763 -4602 12859 -4586
rect 12797 -4636 12835 -4602
rect 12893 -4620 12921 -4586
rect 12955 -4588 12989 -4572
rect 12869 -4636 12921 -4620
rect 13023 -4622 13057 -4484
rect 12205 -4720 12239 -4704
rect 12105 -4772 12171 -4730
rect 12311 -4734 12327 -4700
rect 12361 -4734 12377 -4700
rect 12411 -4728 12460 -4694
rect 12494 -4728 12510 -4694
rect 12551 -4728 12567 -4694
rect 12601 -4728 12722 -4694
rect 12897 -4696 12963 -4680
rect 12311 -4772 12377 -4734
rect 12897 -4730 12913 -4696
rect 12947 -4730 12963 -4696
rect 12897 -4772 12963 -4730
rect 13005 -4700 13057 -4622
rect 13095 -4458 13238 -4456
rect 13272 -4458 13288 -4424
rect 13322 -4440 13356 -4364
rect 13544 -4338 13560 -4304
rect 13594 -4338 13638 -4304
rect 13672 -4338 13688 -4304
rect 13722 -4312 13803 -4296
rect 13954 -4304 13988 -4262
rect 13474 -4372 13508 -4364
rect 13756 -4346 13803 -4312
rect 13474 -4406 13634 -4372
rect 13095 -4490 13230 -4458
rect 13322 -4474 13516 -4440
rect 13550 -4474 13566 -4440
rect 13095 -4598 13137 -4490
rect 13322 -4492 13356 -4474
rect 13095 -4632 13103 -4598
rect 13095 -4648 13137 -4632
rect 13171 -4534 13241 -4524
rect 13171 -4550 13207 -4534
rect 13171 -4584 13199 -4550
rect 13233 -4584 13241 -4568
rect 13171 -4648 13241 -4584
rect 13275 -4526 13356 -4492
rect 13275 -4682 13309 -4526
rect 13423 -4539 13531 -4508
rect 13600 -4524 13634 -4406
rect 13722 -4380 13803 -4346
rect 13756 -4414 13803 -4380
rect 13722 -4448 13803 -4414
rect 13756 -4482 13803 -4448
rect 13722 -4498 13803 -4482
rect 13600 -4530 13689 -4524
rect 13457 -4548 13531 -4539
rect 13343 -4576 13387 -4560
rect 13377 -4610 13387 -4576
rect 13423 -4582 13439 -4573
rect 13473 -4582 13531 -4548
rect 13343 -4616 13387 -4610
rect 13483 -4602 13531 -4582
rect 13343 -4650 13449 -4616
rect 13119 -4696 13309 -4682
rect 13005 -4734 13025 -4700
rect 13059 -4734 13075 -4700
rect 13119 -4730 13135 -4696
rect 13169 -4730 13309 -4696
rect 13119 -4738 13309 -4730
rect 13343 -4700 13381 -4684
rect 13343 -4734 13347 -4700
rect 13415 -4696 13449 -4650
rect 13517 -4636 13531 -4602
rect 13483 -4662 13531 -4636
rect 13565 -4540 13689 -4530
rect 13565 -4574 13639 -4540
rect 13673 -4574 13689 -4540
rect 13565 -4590 13689 -4574
rect 13565 -4625 13630 -4590
rect 13737 -4624 13803 -4498
rect 13565 -4680 13629 -4625
rect 13415 -4714 13565 -4696
rect 13599 -4714 13629 -4680
rect 13415 -4730 13629 -4714
rect 13669 -4657 13703 -4635
rect 13343 -4772 13381 -4734
rect 13669 -4772 13703 -4691
rect 13737 -4658 13753 -4624
rect 13787 -4658 13803 -4624
rect 13737 -4692 13803 -4658
rect 13737 -4726 13753 -4692
rect 13787 -4726 13803 -4692
rect 13841 -4338 13857 -4304
rect 13891 -4338 13907 -4304
rect 13841 -4372 13907 -4338
rect 13841 -4406 13857 -4372
rect 13891 -4406 13907 -4372
rect 13841 -4524 13907 -4406
rect 14136 -4312 14187 -4296
rect 13954 -4372 13988 -4338
rect 13954 -4440 13988 -4406
rect 13954 -4490 13988 -4474
rect 14038 -4340 14089 -4324
rect 14072 -4374 14089 -4340
rect 14038 -4408 14089 -4374
rect 14072 -4442 14089 -4408
rect 14136 -4346 14153 -4312
rect 14136 -4380 14187 -4346
rect 14221 -4328 14287 -4262
rect 14221 -4362 14237 -4328
rect 14271 -4362 14287 -4328
rect 14321 -4312 14355 -4296
rect 14136 -4414 14153 -4380
rect 14321 -4380 14355 -4346
rect 14187 -4414 14286 -4396
rect 14136 -4430 14286 -4414
rect 14038 -4464 14089 -4442
rect 14038 -4500 14206 -4464
rect 14047 -4515 14206 -4500
rect 13841 -4540 14013 -4524
rect 13841 -4574 13979 -4540
rect 13841 -4590 14013 -4574
rect 14047 -4549 14078 -4515
rect 14116 -4540 14206 -4515
rect 14116 -4549 14150 -4540
rect 14047 -4574 14150 -4549
rect 14184 -4574 14206 -4540
rect 13841 -4670 13891 -4590
rect 14047 -4594 14206 -4574
rect 14240 -4525 14286 -4430
rect 14240 -4534 14252 -4525
rect 14274 -4568 14286 -4559
rect 14047 -4630 14089 -4594
rect 14240 -4628 14286 -4568
rect 14038 -4646 14089 -4630
rect 13841 -4704 13857 -4670
rect 13841 -4720 13891 -4704
rect 13954 -4676 13988 -4653
rect 13737 -4734 13803 -4726
rect 13954 -4772 13988 -4710
rect 14072 -4680 14089 -4646
rect 14038 -4736 14089 -4680
rect 14136 -4662 14286 -4628
rect 14136 -4670 14187 -4662
rect 14136 -4704 14153 -4670
rect 14321 -4670 14355 -4432
rect 14389 -4456 14454 -4299
rect 14488 -4304 14538 -4262
rect 14488 -4338 14504 -4304
rect 14488 -4354 14538 -4338
rect 14572 -4312 14622 -4296
rect 14572 -4346 14588 -4312
rect 14572 -4362 14622 -4346
rect 14665 -4306 14801 -4296
rect 14665 -4340 14681 -4306
rect 14715 -4340 14801 -4306
rect 14916 -4314 14982 -4262
rect 15109 -4304 15183 -4262
rect 14665 -4362 14801 -4340
rect 14572 -4388 14606 -4362
rect 14527 -4422 14606 -4388
rect 14640 -4398 14733 -4396
rect 14401 -4479 14493 -4456
rect 14401 -4513 14459 -4479
rect 14401 -4614 14493 -4513
rect 14401 -4648 14425 -4614
rect 14463 -4648 14493 -4614
rect 14401 -4666 14493 -4648
rect 14136 -4720 14187 -4704
rect 14221 -4730 14237 -4696
rect 14271 -4730 14287 -4696
rect 14527 -4694 14561 -4422
rect 14640 -4424 14699 -4398
rect 14674 -4432 14699 -4424
rect 14674 -4458 14733 -4432
rect 14640 -4474 14733 -4458
rect 14595 -4534 14665 -4512
rect 14595 -4568 14607 -4534
rect 14641 -4568 14665 -4534
rect 14595 -4586 14665 -4568
rect 14595 -4620 14618 -4586
rect 14652 -4620 14665 -4586
rect 14595 -4636 14665 -4620
rect 14699 -4592 14733 -4474
rect 14767 -4518 14801 -4362
rect 14835 -4330 14869 -4314
rect 14916 -4348 14932 -4314
rect 14966 -4348 14982 -4314
rect 15016 -4330 15050 -4314
rect 14835 -4382 14869 -4364
rect 15109 -4338 15129 -4304
rect 15163 -4338 15183 -4304
rect 15109 -4354 15183 -4338
rect 15217 -4312 15251 -4296
rect 15016 -4382 15050 -4364
rect 14835 -4416 15050 -4382
rect 15217 -4388 15251 -4346
rect 15298 -4305 15472 -4296
rect 15298 -4339 15314 -4305
rect 15348 -4339 15472 -4305
rect 15298 -4364 15472 -4339
rect 15506 -4304 15556 -4262
rect 15540 -4338 15556 -4304
rect 15660 -4304 15804 -4262
rect 15506 -4354 15556 -4338
rect 15590 -4330 15624 -4314
rect 15139 -4422 15251 -4388
rect 15139 -4450 15173 -4422
rect 14873 -4484 14889 -4450
rect 14923 -4484 15173 -4450
rect 15312 -4432 15323 -4398
rect 15357 -4424 15404 -4398
rect 15312 -4456 15354 -4432
rect 14767 -4538 15105 -4518
rect 14767 -4552 15071 -4538
rect 14699 -4626 14720 -4592
rect 14754 -4626 14770 -4592
rect 14699 -4636 14770 -4626
rect 14804 -4694 14838 -4552
rect 14879 -4602 14975 -4586
rect 14913 -4636 14951 -4602
rect 15009 -4620 15037 -4586
rect 15071 -4588 15105 -4572
rect 14985 -4636 15037 -4620
rect 15139 -4622 15173 -4484
rect 14321 -4720 14355 -4704
rect 14221 -4772 14287 -4730
rect 14427 -4734 14443 -4700
rect 14477 -4734 14493 -4700
rect 14527 -4728 14576 -4694
rect 14610 -4728 14626 -4694
rect 14667 -4728 14683 -4694
rect 14717 -4728 14838 -4694
rect 15013 -4696 15079 -4680
rect 14427 -4772 14493 -4734
rect 15013 -4730 15029 -4696
rect 15063 -4730 15079 -4696
rect 15013 -4772 15079 -4730
rect 15121 -4700 15173 -4622
rect 15211 -4458 15354 -4456
rect 15388 -4458 15404 -4424
rect 15438 -4440 15472 -4364
rect 15660 -4338 15676 -4304
rect 15710 -4338 15754 -4304
rect 15788 -4338 15804 -4304
rect 15838 -4312 15919 -4296
rect 16070 -4304 16104 -4262
rect 15590 -4372 15624 -4364
rect 15872 -4346 15919 -4312
rect 15590 -4406 15750 -4372
rect 15211 -4490 15346 -4458
rect 15438 -4474 15632 -4440
rect 15666 -4474 15682 -4440
rect 15211 -4598 15253 -4490
rect 15438 -4492 15472 -4474
rect 15211 -4632 15219 -4598
rect 15211 -4648 15253 -4632
rect 15287 -4534 15357 -4524
rect 15287 -4550 15323 -4534
rect 15287 -4584 15315 -4550
rect 15349 -4584 15357 -4568
rect 15287 -4648 15357 -4584
rect 15391 -4526 15472 -4492
rect 15391 -4682 15425 -4526
rect 15539 -4539 15647 -4508
rect 15716 -4524 15750 -4406
rect 15838 -4380 15919 -4346
rect 15872 -4414 15919 -4380
rect 15838 -4448 15919 -4414
rect 15872 -4482 15919 -4448
rect 15838 -4498 15919 -4482
rect 15716 -4530 15805 -4524
rect 15573 -4548 15647 -4539
rect 15459 -4576 15503 -4560
rect 15493 -4610 15503 -4576
rect 15539 -4582 15555 -4573
rect 15589 -4582 15647 -4548
rect 15459 -4616 15503 -4610
rect 15599 -4602 15647 -4582
rect 15459 -4650 15565 -4616
rect 15235 -4696 15425 -4682
rect 15121 -4734 15141 -4700
rect 15175 -4734 15191 -4700
rect 15235 -4730 15251 -4696
rect 15285 -4730 15425 -4696
rect 15235 -4738 15425 -4730
rect 15459 -4700 15497 -4684
rect 15459 -4734 15463 -4700
rect 15531 -4696 15565 -4650
rect 15633 -4636 15647 -4602
rect 15599 -4662 15647 -4636
rect 15681 -4540 15805 -4530
rect 15681 -4574 15755 -4540
rect 15789 -4574 15805 -4540
rect 15681 -4590 15805 -4574
rect 15681 -4625 15746 -4590
rect 15853 -4624 15919 -4498
rect 15681 -4680 15745 -4625
rect 15531 -4714 15681 -4696
rect 15715 -4714 15745 -4680
rect 15531 -4730 15745 -4714
rect 15785 -4657 15819 -4635
rect 15459 -4772 15497 -4734
rect 15785 -4772 15819 -4691
rect 15853 -4658 15869 -4624
rect 15903 -4658 15919 -4624
rect 15853 -4692 15919 -4658
rect 15853 -4726 15869 -4692
rect 15903 -4726 15919 -4692
rect 15957 -4338 15973 -4304
rect 16007 -4338 16023 -4304
rect 15957 -4372 16023 -4338
rect 15957 -4406 15973 -4372
rect 16007 -4406 16023 -4372
rect 15957 -4524 16023 -4406
rect 16252 -4312 16303 -4296
rect 16070 -4372 16104 -4338
rect 16070 -4440 16104 -4406
rect 16070 -4490 16104 -4474
rect 16154 -4340 16205 -4324
rect 16188 -4374 16205 -4340
rect 16154 -4408 16205 -4374
rect 16188 -4442 16205 -4408
rect 16252 -4346 16269 -4312
rect 16252 -4380 16303 -4346
rect 16337 -4328 16403 -4262
rect 16337 -4362 16353 -4328
rect 16387 -4362 16403 -4328
rect 16437 -4312 16471 -4296
rect 16252 -4414 16269 -4380
rect 16437 -4380 16471 -4346
rect 16303 -4414 16402 -4396
rect 16252 -4430 16402 -4414
rect 16154 -4464 16205 -4442
rect 16154 -4500 16322 -4464
rect 16163 -4515 16322 -4500
rect 15957 -4540 16129 -4524
rect 15957 -4574 16095 -4540
rect 15957 -4590 16129 -4574
rect 16163 -4549 16194 -4515
rect 16232 -4540 16322 -4515
rect 16232 -4549 16266 -4540
rect 16163 -4574 16266 -4549
rect 16300 -4574 16322 -4540
rect 15957 -4670 16007 -4590
rect 16163 -4594 16322 -4574
rect 16356 -4525 16402 -4430
rect 16356 -4534 16368 -4525
rect 16390 -4568 16402 -4559
rect 16163 -4630 16205 -4594
rect 16356 -4628 16402 -4568
rect 16154 -4646 16205 -4630
rect 15957 -4704 15973 -4670
rect 15957 -4720 16007 -4704
rect 16070 -4676 16104 -4653
rect 15853 -4734 15919 -4726
rect 16070 -4772 16104 -4710
rect 16188 -4680 16205 -4646
rect 16154 -4736 16205 -4680
rect 16252 -4662 16402 -4628
rect 16252 -4670 16303 -4662
rect 16252 -4704 16269 -4670
rect 16437 -4670 16471 -4432
rect 16505 -4456 16570 -4299
rect 16604 -4304 16654 -4262
rect 16604 -4338 16620 -4304
rect 16604 -4354 16654 -4338
rect 16688 -4312 16738 -4296
rect 16688 -4346 16704 -4312
rect 16688 -4362 16738 -4346
rect 16781 -4306 16917 -4296
rect 16781 -4340 16797 -4306
rect 16831 -4340 16917 -4306
rect 17032 -4314 17098 -4262
rect 17225 -4304 17299 -4262
rect 16781 -4362 16917 -4340
rect 16688 -4388 16722 -4362
rect 16643 -4422 16722 -4388
rect 16756 -4398 16849 -4396
rect 16517 -4479 16609 -4456
rect 16517 -4513 16575 -4479
rect 16517 -4614 16609 -4513
rect 16517 -4648 16541 -4614
rect 16579 -4648 16609 -4614
rect 16517 -4666 16609 -4648
rect 16252 -4720 16303 -4704
rect 16337 -4730 16353 -4696
rect 16387 -4730 16403 -4696
rect 16643 -4694 16677 -4422
rect 16756 -4424 16815 -4398
rect 16790 -4432 16815 -4424
rect 16790 -4458 16849 -4432
rect 16756 -4474 16849 -4458
rect 16711 -4534 16781 -4512
rect 16711 -4568 16723 -4534
rect 16757 -4568 16781 -4534
rect 16711 -4586 16781 -4568
rect 16711 -4620 16734 -4586
rect 16768 -4620 16781 -4586
rect 16711 -4636 16781 -4620
rect 16815 -4592 16849 -4474
rect 16883 -4518 16917 -4362
rect 16951 -4330 16985 -4314
rect 17032 -4348 17048 -4314
rect 17082 -4348 17098 -4314
rect 17132 -4330 17166 -4314
rect 16951 -4382 16985 -4364
rect 17225 -4338 17245 -4304
rect 17279 -4338 17299 -4304
rect 17225 -4354 17299 -4338
rect 17333 -4312 17367 -4296
rect 17132 -4382 17166 -4364
rect 16951 -4416 17166 -4382
rect 17333 -4388 17367 -4346
rect 17414 -4305 17588 -4296
rect 17414 -4339 17430 -4305
rect 17464 -4339 17588 -4305
rect 17414 -4364 17588 -4339
rect 17622 -4304 17672 -4262
rect 17656 -4338 17672 -4304
rect 17776 -4304 17920 -4262
rect 17622 -4354 17672 -4338
rect 17706 -4330 17740 -4314
rect 17255 -4422 17367 -4388
rect 17255 -4450 17289 -4422
rect 16989 -4484 17005 -4450
rect 17039 -4484 17289 -4450
rect 17428 -4432 17439 -4398
rect 17473 -4424 17520 -4398
rect 17428 -4456 17470 -4432
rect 16883 -4538 17221 -4518
rect 16883 -4552 17187 -4538
rect 16815 -4626 16836 -4592
rect 16870 -4626 16886 -4592
rect 16815 -4636 16886 -4626
rect 16920 -4694 16954 -4552
rect 16995 -4602 17091 -4586
rect 17029 -4636 17067 -4602
rect 17125 -4620 17153 -4586
rect 17187 -4588 17221 -4572
rect 17101 -4636 17153 -4620
rect 17255 -4622 17289 -4484
rect 16437 -4720 16471 -4704
rect 16337 -4772 16403 -4730
rect 16543 -4734 16559 -4700
rect 16593 -4734 16609 -4700
rect 16643 -4728 16692 -4694
rect 16726 -4728 16742 -4694
rect 16783 -4728 16799 -4694
rect 16833 -4728 16954 -4694
rect 17129 -4696 17195 -4680
rect 16543 -4772 16609 -4734
rect 17129 -4730 17145 -4696
rect 17179 -4730 17195 -4696
rect 17129 -4772 17195 -4730
rect 17237 -4700 17289 -4622
rect 17327 -4458 17470 -4456
rect 17504 -4458 17520 -4424
rect 17554 -4440 17588 -4364
rect 17776 -4338 17792 -4304
rect 17826 -4338 17870 -4304
rect 17904 -4338 17920 -4304
rect 17954 -4312 18035 -4296
rect 18186 -4304 18220 -4262
rect 17706 -4372 17740 -4364
rect 17988 -4346 18035 -4312
rect 17706 -4406 17866 -4372
rect 17327 -4490 17462 -4458
rect 17554 -4474 17748 -4440
rect 17782 -4474 17798 -4440
rect 17327 -4598 17369 -4490
rect 17554 -4492 17588 -4474
rect 17327 -4632 17335 -4598
rect 17327 -4648 17369 -4632
rect 17403 -4534 17473 -4524
rect 17403 -4550 17439 -4534
rect 17403 -4584 17431 -4550
rect 17465 -4584 17473 -4568
rect 17403 -4648 17473 -4584
rect 17507 -4526 17588 -4492
rect 17507 -4682 17541 -4526
rect 17655 -4539 17763 -4508
rect 17832 -4524 17866 -4406
rect 17954 -4380 18035 -4346
rect 17988 -4414 18035 -4380
rect 17954 -4448 18035 -4414
rect 17988 -4482 18035 -4448
rect 17954 -4498 18035 -4482
rect 17832 -4530 17921 -4524
rect 17689 -4548 17763 -4539
rect 17575 -4576 17619 -4560
rect 17609 -4610 17619 -4576
rect 17655 -4582 17671 -4573
rect 17705 -4582 17763 -4548
rect 17575 -4616 17619 -4610
rect 17715 -4602 17763 -4582
rect 17575 -4650 17681 -4616
rect 17351 -4696 17541 -4682
rect 17237 -4734 17257 -4700
rect 17291 -4734 17307 -4700
rect 17351 -4730 17367 -4696
rect 17401 -4730 17541 -4696
rect 17351 -4738 17541 -4730
rect 17575 -4700 17613 -4684
rect 17575 -4734 17579 -4700
rect 17647 -4696 17681 -4650
rect 17749 -4636 17763 -4602
rect 17715 -4662 17763 -4636
rect 17797 -4540 17921 -4530
rect 17797 -4574 17871 -4540
rect 17905 -4574 17921 -4540
rect 17797 -4590 17921 -4574
rect 17797 -4625 17862 -4590
rect 17969 -4624 18035 -4498
rect 17797 -4680 17861 -4625
rect 17647 -4714 17797 -4696
rect 17831 -4714 17861 -4680
rect 17647 -4730 17861 -4714
rect 17901 -4657 17935 -4635
rect 17575 -4772 17613 -4734
rect 17901 -4772 17935 -4691
rect 17969 -4658 17985 -4624
rect 18019 -4658 18035 -4624
rect 17969 -4692 18035 -4658
rect 17969 -4726 17985 -4692
rect 18019 -4726 18035 -4692
rect 18073 -4338 18089 -4304
rect 18123 -4338 18139 -4304
rect 18073 -4372 18139 -4338
rect 18073 -4406 18089 -4372
rect 18123 -4406 18139 -4372
rect 18073 -4524 18139 -4406
rect 18368 -4312 18419 -4296
rect 18186 -4372 18220 -4338
rect 18186 -4440 18220 -4406
rect 18186 -4490 18220 -4474
rect 18270 -4340 18321 -4324
rect 18304 -4374 18321 -4340
rect 18270 -4408 18321 -4374
rect 18304 -4442 18321 -4408
rect 18368 -4346 18385 -4312
rect 18368 -4380 18419 -4346
rect 18453 -4328 18519 -4262
rect 18453 -4362 18469 -4328
rect 18503 -4362 18519 -4328
rect 18553 -4312 18587 -4296
rect 18368 -4414 18385 -4380
rect 18553 -4380 18587 -4346
rect 18419 -4414 18518 -4396
rect 18368 -4430 18518 -4414
rect 18270 -4464 18321 -4442
rect 18270 -4500 18438 -4464
rect 18279 -4515 18438 -4500
rect 18073 -4540 18245 -4524
rect 18073 -4574 18211 -4540
rect 18073 -4590 18245 -4574
rect 18279 -4549 18310 -4515
rect 18348 -4540 18438 -4515
rect 18348 -4549 18382 -4540
rect 18279 -4574 18382 -4549
rect 18416 -4574 18438 -4540
rect 18073 -4670 18123 -4590
rect 18279 -4594 18438 -4574
rect 18472 -4525 18518 -4430
rect 18472 -4534 18484 -4525
rect 18506 -4568 18518 -4559
rect 18279 -4630 18321 -4594
rect 18472 -4628 18518 -4568
rect 18270 -4646 18321 -4630
rect 18073 -4704 18089 -4670
rect 18073 -4720 18123 -4704
rect 18186 -4676 18220 -4653
rect 17969 -4734 18035 -4726
rect 18186 -4772 18220 -4710
rect 18304 -4680 18321 -4646
rect 18270 -4736 18321 -4680
rect 18368 -4662 18518 -4628
rect 18368 -4670 18419 -4662
rect 18368 -4704 18385 -4670
rect 18553 -4670 18587 -4432
rect 18621 -4456 18686 -4299
rect 18720 -4304 18770 -4262
rect 18720 -4338 18736 -4304
rect 18720 -4354 18770 -4338
rect 18804 -4312 18854 -4296
rect 18804 -4346 18820 -4312
rect 18804 -4362 18854 -4346
rect 18897 -4306 19033 -4296
rect 18897 -4340 18913 -4306
rect 18947 -4340 19033 -4306
rect 19148 -4314 19214 -4262
rect 19341 -4304 19415 -4262
rect 18897 -4362 19033 -4340
rect 18804 -4388 18838 -4362
rect 18759 -4422 18838 -4388
rect 18872 -4398 18965 -4396
rect 18633 -4479 18725 -4456
rect 18633 -4513 18691 -4479
rect 18633 -4614 18725 -4513
rect 18633 -4648 18657 -4614
rect 18695 -4648 18725 -4614
rect 18633 -4666 18725 -4648
rect 18368 -4720 18419 -4704
rect 18453 -4730 18469 -4696
rect 18503 -4730 18519 -4696
rect 18759 -4694 18793 -4422
rect 18872 -4424 18931 -4398
rect 18906 -4432 18931 -4424
rect 18906 -4458 18965 -4432
rect 18872 -4474 18965 -4458
rect 18827 -4534 18897 -4512
rect 18827 -4568 18839 -4534
rect 18873 -4568 18897 -4534
rect 18827 -4586 18897 -4568
rect 18827 -4620 18850 -4586
rect 18884 -4620 18897 -4586
rect 18827 -4636 18897 -4620
rect 18931 -4592 18965 -4474
rect 18999 -4518 19033 -4362
rect 19067 -4330 19101 -4314
rect 19148 -4348 19164 -4314
rect 19198 -4348 19214 -4314
rect 19248 -4330 19282 -4314
rect 19067 -4382 19101 -4364
rect 19341 -4338 19361 -4304
rect 19395 -4338 19415 -4304
rect 19341 -4354 19415 -4338
rect 19449 -4312 19483 -4296
rect 19248 -4382 19282 -4364
rect 19067 -4416 19282 -4382
rect 19449 -4388 19483 -4346
rect 19530 -4305 19704 -4296
rect 19530 -4339 19546 -4305
rect 19580 -4339 19704 -4305
rect 19530 -4364 19704 -4339
rect 19738 -4304 19788 -4262
rect 19772 -4338 19788 -4304
rect 19892 -4304 20036 -4262
rect 19738 -4354 19788 -4338
rect 19822 -4330 19856 -4314
rect 19371 -4422 19483 -4388
rect 19371 -4450 19405 -4422
rect 19105 -4484 19121 -4450
rect 19155 -4484 19405 -4450
rect 19544 -4432 19555 -4398
rect 19589 -4424 19636 -4398
rect 19544 -4456 19586 -4432
rect 18999 -4538 19337 -4518
rect 18999 -4552 19303 -4538
rect 18931 -4626 18952 -4592
rect 18986 -4626 19002 -4592
rect 18931 -4636 19002 -4626
rect 19036 -4694 19070 -4552
rect 19111 -4602 19207 -4586
rect 19145 -4636 19183 -4602
rect 19241 -4620 19269 -4586
rect 19303 -4588 19337 -4572
rect 19217 -4636 19269 -4620
rect 19371 -4622 19405 -4484
rect 18553 -4720 18587 -4704
rect 18453 -4772 18519 -4730
rect 18659 -4734 18675 -4700
rect 18709 -4734 18725 -4700
rect 18759 -4728 18808 -4694
rect 18842 -4728 18858 -4694
rect 18899 -4728 18915 -4694
rect 18949 -4728 19070 -4694
rect 19245 -4696 19311 -4680
rect 18659 -4772 18725 -4734
rect 19245 -4730 19261 -4696
rect 19295 -4730 19311 -4696
rect 19245 -4772 19311 -4730
rect 19353 -4700 19405 -4622
rect 19443 -4458 19586 -4456
rect 19620 -4458 19636 -4424
rect 19670 -4440 19704 -4364
rect 19892 -4338 19908 -4304
rect 19942 -4338 19986 -4304
rect 20020 -4338 20036 -4304
rect 20070 -4312 20151 -4296
rect 20302 -4304 20336 -4262
rect 19822 -4372 19856 -4364
rect 20104 -4346 20151 -4312
rect 19822 -4406 19982 -4372
rect 19443 -4490 19578 -4458
rect 19670 -4474 19864 -4440
rect 19898 -4474 19914 -4440
rect 19443 -4598 19485 -4490
rect 19670 -4492 19704 -4474
rect 19443 -4632 19451 -4598
rect 19443 -4648 19485 -4632
rect 19519 -4534 19589 -4524
rect 19519 -4550 19555 -4534
rect 19519 -4584 19547 -4550
rect 19581 -4584 19589 -4568
rect 19519 -4648 19589 -4584
rect 19623 -4526 19704 -4492
rect 19623 -4682 19657 -4526
rect 19771 -4539 19879 -4508
rect 19948 -4524 19982 -4406
rect 20070 -4380 20151 -4346
rect 20104 -4414 20151 -4380
rect 20070 -4448 20151 -4414
rect 20104 -4482 20151 -4448
rect 20070 -4498 20151 -4482
rect 19948 -4530 20037 -4524
rect 19805 -4548 19879 -4539
rect 19691 -4576 19735 -4560
rect 19725 -4610 19735 -4576
rect 19771 -4582 19787 -4573
rect 19821 -4582 19879 -4548
rect 19691 -4616 19735 -4610
rect 19831 -4602 19879 -4582
rect 19691 -4650 19797 -4616
rect 19467 -4696 19657 -4682
rect 19353 -4734 19373 -4700
rect 19407 -4734 19423 -4700
rect 19467 -4730 19483 -4696
rect 19517 -4730 19657 -4696
rect 19467 -4738 19657 -4730
rect 19691 -4700 19729 -4684
rect 19691 -4734 19695 -4700
rect 19763 -4696 19797 -4650
rect 19865 -4636 19879 -4602
rect 19831 -4662 19879 -4636
rect 19913 -4540 20037 -4530
rect 19913 -4574 19987 -4540
rect 20021 -4574 20037 -4540
rect 19913 -4590 20037 -4574
rect 19913 -4625 19978 -4590
rect 20085 -4624 20151 -4498
rect 19913 -4680 19977 -4625
rect 19763 -4714 19913 -4696
rect 19947 -4714 19977 -4680
rect 19763 -4730 19977 -4714
rect 20017 -4657 20051 -4635
rect 19691 -4772 19729 -4734
rect 20017 -4772 20051 -4691
rect 20085 -4658 20101 -4624
rect 20135 -4658 20151 -4624
rect 20085 -4692 20151 -4658
rect 20085 -4726 20101 -4692
rect 20135 -4726 20151 -4692
rect 20189 -4338 20205 -4304
rect 20239 -4338 20255 -4304
rect 20189 -4372 20255 -4338
rect 20189 -4406 20205 -4372
rect 20239 -4406 20255 -4372
rect 20189 -4524 20255 -4406
rect 20484 -4312 20535 -4296
rect 20302 -4372 20336 -4338
rect 20302 -4440 20336 -4406
rect 20302 -4490 20336 -4474
rect 20386 -4340 20437 -4324
rect 20420 -4374 20437 -4340
rect 20386 -4408 20437 -4374
rect 20420 -4442 20437 -4408
rect 20484 -4346 20501 -4312
rect 20484 -4380 20535 -4346
rect 20569 -4328 20635 -4262
rect 20569 -4362 20585 -4328
rect 20619 -4362 20635 -4328
rect 20669 -4312 20703 -4296
rect 20484 -4414 20501 -4380
rect 20669 -4380 20703 -4346
rect 20535 -4414 20634 -4396
rect 20484 -4430 20634 -4414
rect 20386 -4464 20437 -4442
rect 20386 -4500 20554 -4464
rect 20395 -4515 20554 -4500
rect 20189 -4540 20361 -4524
rect 20189 -4574 20327 -4540
rect 20189 -4590 20361 -4574
rect 20395 -4549 20426 -4515
rect 20464 -4540 20554 -4515
rect 20464 -4549 20498 -4540
rect 20395 -4574 20498 -4549
rect 20532 -4574 20554 -4540
rect 20189 -4670 20239 -4590
rect 20395 -4594 20554 -4574
rect 20588 -4525 20634 -4430
rect 20588 -4534 20600 -4525
rect 20622 -4568 20634 -4559
rect 20395 -4630 20437 -4594
rect 20588 -4628 20634 -4568
rect 20386 -4646 20437 -4630
rect 20189 -4704 20205 -4670
rect 20189 -4720 20239 -4704
rect 20302 -4676 20336 -4653
rect 20085 -4734 20151 -4726
rect 20302 -4772 20336 -4710
rect 20420 -4680 20437 -4646
rect 20386 -4736 20437 -4680
rect 20484 -4662 20634 -4628
rect 20484 -4670 20535 -4662
rect 20484 -4704 20501 -4670
rect 20669 -4670 20703 -4432
rect 20737 -4456 20802 -4299
rect 20836 -4304 20886 -4262
rect 20836 -4338 20852 -4304
rect 20836 -4354 20886 -4338
rect 20920 -4312 20970 -4296
rect 20920 -4346 20936 -4312
rect 20920 -4362 20970 -4346
rect 21013 -4306 21149 -4296
rect 21013 -4340 21029 -4306
rect 21063 -4340 21149 -4306
rect 21264 -4314 21330 -4262
rect 21457 -4304 21531 -4262
rect 21013 -4362 21149 -4340
rect 20920 -4388 20954 -4362
rect 20875 -4422 20954 -4388
rect 20988 -4398 21081 -4396
rect 20749 -4479 20841 -4456
rect 20749 -4513 20807 -4479
rect 20749 -4614 20841 -4513
rect 20749 -4648 20773 -4614
rect 20811 -4648 20841 -4614
rect 20749 -4666 20841 -4648
rect 20484 -4720 20535 -4704
rect 20569 -4730 20585 -4696
rect 20619 -4730 20635 -4696
rect 20875 -4694 20909 -4422
rect 20988 -4424 21047 -4398
rect 21022 -4432 21047 -4424
rect 21022 -4458 21081 -4432
rect 20988 -4474 21081 -4458
rect 20943 -4534 21013 -4512
rect 20943 -4568 20955 -4534
rect 20989 -4568 21013 -4534
rect 20943 -4586 21013 -4568
rect 20943 -4620 20966 -4586
rect 21000 -4620 21013 -4586
rect 20943 -4636 21013 -4620
rect 21047 -4592 21081 -4474
rect 21115 -4518 21149 -4362
rect 21183 -4330 21217 -4314
rect 21264 -4348 21280 -4314
rect 21314 -4348 21330 -4314
rect 21364 -4330 21398 -4314
rect 21183 -4382 21217 -4364
rect 21457 -4338 21477 -4304
rect 21511 -4338 21531 -4304
rect 21457 -4354 21531 -4338
rect 21565 -4312 21599 -4296
rect 21364 -4382 21398 -4364
rect 21183 -4416 21398 -4382
rect 21565 -4388 21599 -4346
rect 21646 -4305 21820 -4296
rect 21646 -4339 21662 -4305
rect 21696 -4339 21820 -4305
rect 21646 -4364 21820 -4339
rect 21854 -4304 21904 -4262
rect 21888 -4338 21904 -4304
rect 22008 -4304 22152 -4262
rect 21854 -4354 21904 -4338
rect 21938 -4330 21972 -4314
rect 21487 -4422 21599 -4388
rect 21487 -4450 21521 -4422
rect 21221 -4484 21237 -4450
rect 21271 -4484 21521 -4450
rect 21660 -4432 21671 -4398
rect 21705 -4424 21752 -4398
rect 21660 -4456 21702 -4432
rect 21115 -4538 21453 -4518
rect 21115 -4552 21419 -4538
rect 21047 -4626 21068 -4592
rect 21102 -4626 21118 -4592
rect 21047 -4636 21118 -4626
rect 21152 -4694 21186 -4552
rect 21227 -4602 21323 -4586
rect 21261 -4636 21299 -4602
rect 21357 -4620 21385 -4586
rect 21419 -4588 21453 -4572
rect 21333 -4636 21385 -4620
rect 21487 -4622 21521 -4484
rect 20669 -4720 20703 -4704
rect 20569 -4772 20635 -4730
rect 20775 -4734 20791 -4700
rect 20825 -4734 20841 -4700
rect 20875 -4728 20924 -4694
rect 20958 -4728 20974 -4694
rect 21015 -4728 21031 -4694
rect 21065 -4728 21186 -4694
rect 21361 -4696 21427 -4680
rect 20775 -4772 20841 -4734
rect 21361 -4730 21377 -4696
rect 21411 -4730 21427 -4696
rect 21361 -4772 21427 -4730
rect 21469 -4700 21521 -4622
rect 21559 -4458 21702 -4456
rect 21736 -4458 21752 -4424
rect 21786 -4440 21820 -4364
rect 22008 -4338 22024 -4304
rect 22058 -4338 22102 -4304
rect 22136 -4338 22152 -4304
rect 22186 -4312 22267 -4296
rect 22418 -4304 22452 -4262
rect 21938 -4372 21972 -4364
rect 22220 -4346 22267 -4312
rect 21938 -4406 22098 -4372
rect 21559 -4490 21694 -4458
rect 21786 -4474 21980 -4440
rect 22014 -4474 22030 -4440
rect 21559 -4598 21601 -4490
rect 21786 -4492 21820 -4474
rect 21559 -4632 21567 -4598
rect 21559 -4648 21601 -4632
rect 21635 -4534 21705 -4524
rect 21635 -4550 21671 -4534
rect 21635 -4584 21663 -4550
rect 21697 -4584 21705 -4568
rect 21635 -4648 21705 -4584
rect 21739 -4526 21820 -4492
rect 21739 -4682 21773 -4526
rect 21887 -4539 21995 -4508
rect 22064 -4524 22098 -4406
rect 22186 -4380 22267 -4346
rect 22220 -4414 22267 -4380
rect 22186 -4448 22267 -4414
rect 22220 -4482 22267 -4448
rect 22186 -4498 22267 -4482
rect 22064 -4530 22153 -4524
rect 21921 -4548 21995 -4539
rect 21807 -4576 21851 -4560
rect 21841 -4610 21851 -4576
rect 21887 -4582 21903 -4573
rect 21937 -4582 21995 -4548
rect 21807 -4616 21851 -4610
rect 21947 -4602 21995 -4582
rect 21807 -4650 21913 -4616
rect 21583 -4696 21773 -4682
rect 21469 -4734 21489 -4700
rect 21523 -4734 21539 -4700
rect 21583 -4730 21599 -4696
rect 21633 -4730 21773 -4696
rect 21583 -4738 21773 -4730
rect 21807 -4700 21845 -4684
rect 21807 -4734 21811 -4700
rect 21879 -4696 21913 -4650
rect 21981 -4636 21995 -4602
rect 21947 -4662 21995 -4636
rect 22029 -4540 22153 -4530
rect 22029 -4574 22103 -4540
rect 22137 -4574 22153 -4540
rect 22029 -4590 22153 -4574
rect 22029 -4625 22094 -4590
rect 22201 -4624 22267 -4498
rect 22029 -4680 22093 -4625
rect 21879 -4714 22029 -4696
rect 22063 -4714 22093 -4680
rect 21879 -4730 22093 -4714
rect 22133 -4657 22167 -4635
rect 21807 -4772 21845 -4734
rect 22133 -4772 22167 -4691
rect 22201 -4658 22217 -4624
rect 22251 -4658 22267 -4624
rect 22201 -4692 22267 -4658
rect 22201 -4726 22217 -4692
rect 22251 -4726 22267 -4692
rect 22305 -4338 22321 -4304
rect 22355 -4338 22371 -4304
rect 22305 -4372 22371 -4338
rect 22305 -4406 22321 -4372
rect 22355 -4406 22371 -4372
rect 22305 -4524 22371 -4406
rect 22600 -4312 22651 -4296
rect 22418 -4372 22452 -4338
rect 22418 -4440 22452 -4406
rect 22418 -4490 22452 -4474
rect 22502 -4340 22553 -4324
rect 22536 -4374 22553 -4340
rect 22502 -4408 22553 -4374
rect 22536 -4442 22553 -4408
rect 22600 -4346 22617 -4312
rect 22600 -4380 22651 -4346
rect 22685 -4328 22751 -4262
rect 22685 -4362 22701 -4328
rect 22735 -4362 22751 -4328
rect 22785 -4312 22819 -4296
rect 22600 -4414 22617 -4380
rect 22785 -4380 22819 -4346
rect 22651 -4414 22750 -4396
rect 22600 -4430 22750 -4414
rect 22502 -4464 22553 -4442
rect 22502 -4500 22670 -4464
rect 22511 -4515 22670 -4500
rect 22305 -4540 22477 -4524
rect 22305 -4574 22443 -4540
rect 22305 -4590 22477 -4574
rect 22511 -4549 22542 -4515
rect 22580 -4540 22670 -4515
rect 22580 -4549 22614 -4540
rect 22511 -4574 22614 -4549
rect 22648 -4574 22670 -4540
rect 22305 -4670 22355 -4590
rect 22511 -4594 22670 -4574
rect 22704 -4525 22750 -4430
rect 22704 -4534 22716 -4525
rect 22738 -4568 22750 -4559
rect 22511 -4630 22553 -4594
rect 22704 -4628 22750 -4568
rect 22502 -4646 22553 -4630
rect 22305 -4704 22321 -4670
rect 22305 -4720 22355 -4704
rect 22418 -4676 22452 -4653
rect 22201 -4734 22267 -4726
rect 22418 -4772 22452 -4710
rect 22536 -4680 22553 -4646
rect 22502 -4736 22553 -4680
rect 22600 -4662 22750 -4628
rect 22600 -4670 22651 -4662
rect 22600 -4704 22617 -4670
rect 22785 -4670 22819 -4432
rect 22853 -4456 22918 -4299
rect 22952 -4304 23002 -4262
rect 22952 -4338 22968 -4304
rect 22952 -4354 23002 -4338
rect 23036 -4312 23086 -4296
rect 23036 -4346 23052 -4312
rect 23036 -4362 23086 -4346
rect 23129 -4306 23265 -4296
rect 23129 -4340 23145 -4306
rect 23179 -4340 23265 -4306
rect 23380 -4314 23446 -4262
rect 23573 -4304 23647 -4262
rect 23129 -4362 23265 -4340
rect 23036 -4388 23070 -4362
rect 22991 -4422 23070 -4388
rect 23104 -4398 23197 -4396
rect 22865 -4479 22957 -4456
rect 22865 -4513 22923 -4479
rect 22865 -4614 22957 -4513
rect 22865 -4648 22889 -4614
rect 22927 -4648 22957 -4614
rect 22865 -4666 22957 -4648
rect 22600 -4720 22651 -4704
rect 22685 -4730 22701 -4696
rect 22735 -4730 22751 -4696
rect 22991 -4694 23025 -4422
rect 23104 -4424 23163 -4398
rect 23138 -4432 23163 -4424
rect 23138 -4458 23197 -4432
rect 23104 -4474 23197 -4458
rect 23059 -4534 23129 -4512
rect 23059 -4568 23071 -4534
rect 23105 -4568 23129 -4534
rect 23059 -4586 23129 -4568
rect 23059 -4620 23082 -4586
rect 23116 -4620 23129 -4586
rect 23059 -4636 23129 -4620
rect 23163 -4592 23197 -4474
rect 23231 -4518 23265 -4362
rect 23299 -4330 23333 -4314
rect 23380 -4348 23396 -4314
rect 23430 -4348 23446 -4314
rect 23480 -4330 23514 -4314
rect 23299 -4382 23333 -4364
rect 23573 -4338 23593 -4304
rect 23627 -4338 23647 -4304
rect 23573 -4354 23647 -4338
rect 23681 -4312 23715 -4296
rect 23480 -4382 23514 -4364
rect 23299 -4416 23514 -4382
rect 23681 -4388 23715 -4346
rect 23762 -4305 23936 -4296
rect 23762 -4339 23778 -4305
rect 23812 -4339 23936 -4305
rect 23762 -4364 23936 -4339
rect 23970 -4304 24020 -4262
rect 24004 -4338 24020 -4304
rect 24124 -4304 24268 -4262
rect 23970 -4354 24020 -4338
rect 24054 -4330 24088 -4314
rect 23603 -4422 23715 -4388
rect 23603 -4450 23637 -4422
rect 23337 -4484 23353 -4450
rect 23387 -4484 23637 -4450
rect 23776 -4432 23787 -4398
rect 23821 -4424 23868 -4398
rect 23776 -4456 23818 -4432
rect 23231 -4538 23569 -4518
rect 23231 -4552 23535 -4538
rect 23163 -4626 23184 -4592
rect 23218 -4626 23234 -4592
rect 23163 -4636 23234 -4626
rect 23268 -4694 23302 -4552
rect 23343 -4602 23439 -4586
rect 23377 -4636 23415 -4602
rect 23473 -4620 23501 -4586
rect 23535 -4588 23569 -4572
rect 23449 -4636 23501 -4620
rect 23603 -4622 23637 -4484
rect 22785 -4720 22819 -4704
rect 22685 -4772 22751 -4730
rect 22891 -4734 22907 -4700
rect 22941 -4734 22957 -4700
rect 22991 -4728 23040 -4694
rect 23074 -4728 23090 -4694
rect 23131 -4728 23147 -4694
rect 23181 -4728 23302 -4694
rect 23477 -4696 23543 -4680
rect 22891 -4772 22957 -4734
rect 23477 -4730 23493 -4696
rect 23527 -4730 23543 -4696
rect 23477 -4772 23543 -4730
rect 23585 -4700 23637 -4622
rect 23675 -4458 23818 -4456
rect 23852 -4458 23868 -4424
rect 23902 -4440 23936 -4364
rect 24124 -4338 24140 -4304
rect 24174 -4338 24218 -4304
rect 24252 -4338 24268 -4304
rect 24302 -4312 24383 -4296
rect 24534 -4304 24568 -4262
rect 24054 -4372 24088 -4364
rect 24336 -4346 24383 -4312
rect 24054 -4406 24214 -4372
rect 23675 -4490 23810 -4458
rect 23902 -4474 24096 -4440
rect 24130 -4474 24146 -4440
rect 23675 -4598 23717 -4490
rect 23902 -4492 23936 -4474
rect 23675 -4632 23683 -4598
rect 23675 -4648 23717 -4632
rect 23751 -4534 23821 -4524
rect 23751 -4550 23787 -4534
rect 23751 -4584 23779 -4550
rect 23813 -4584 23821 -4568
rect 23751 -4648 23821 -4584
rect 23855 -4526 23936 -4492
rect 23855 -4682 23889 -4526
rect 24003 -4539 24111 -4508
rect 24180 -4524 24214 -4406
rect 24302 -4380 24383 -4346
rect 24336 -4414 24383 -4380
rect 24302 -4448 24383 -4414
rect 24336 -4482 24383 -4448
rect 24302 -4498 24383 -4482
rect 24180 -4530 24269 -4524
rect 24037 -4548 24111 -4539
rect 23923 -4576 23967 -4560
rect 23957 -4610 23967 -4576
rect 24003 -4582 24019 -4573
rect 24053 -4582 24111 -4548
rect 23923 -4616 23967 -4610
rect 24063 -4602 24111 -4582
rect 23923 -4650 24029 -4616
rect 23699 -4696 23889 -4682
rect 23585 -4734 23605 -4700
rect 23639 -4734 23655 -4700
rect 23699 -4730 23715 -4696
rect 23749 -4730 23889 -4696
rect 23699 -4738 23889 -4730
rect 23923 -4700 23961 -4684
rect 23923 -4734 23927 -4700
rect 23995 -4696 24029 -4650
rect 24097 -4636 24111 -4602
rect 24063 -4662 24111 -4636
rect 24145 -4540 24269 -4530
rect 24145 -4574 24219 -4540
rect 24253 -4574 24269 -4540
rect 24145 -4590 24269 -4574
rect 24145 -4625 24210 -4590
rect 24317 -4624 24383 -4498
rect 24145 -4680 24209 -4625
rect 23995 -4714 24145 -4696
rect 24179 -4714 24209 -4680
rect 23995 -4730 24209 -4714
rect 24249 -4657 24283 -4635
rect 23923 -4772 23961 -4734
rect 24249 -4772 24283 -4691
rect 24317 -4658 24333 -4624
rect 24367 -4658 24383 -4624
rect 24317 -4692 24383 -4658
rect 24317 -4726 24333 -4692
rect 24367 -4726 24383 -4692
rect 24421 -4338 24437 -4304
rect 24471 -4338 24487 -4304
rect 24421 -4372 24487 -4338
rect 24421 -4406 24437 -4372
rect 24471 -4406 24487 -4372
rect 24421 -4524 24487 -4406
rect 24716 -4312 24767 -4296
rect 24534 -4372 24568 -4338
rect 24534 -4440 24568 -4406
rect 24534 -4490 24568 -4474
rect 24618 -4340 24669 -4324
rect 24652 -4374 24669 -4340
rect 24618 -4408 24669 -4374
rect 24652 -4442 24669 -4408
rect 24716 -4346 24733 -4312
rect 24716 -4380 24767 -4346
rect 24801 -4328 24867 -4262
rect 24801 -4362 24817 -4328
rect 24851 -4362 24867 -4328
rect 24901 -4312 24935 -4296
rect 24716 -4414 24733 -4380
rect 24901 -4380 24935 -4346
rect 24767 -4414 24866 -4396
rect 24716 -4430 24866 -4414
rect 24618 -4464 24669 -4442
rect 24618 -4500 24786 -4464
rect 24627 -4515 24786 -4500
rect 24421 -4540 24593 -4524
rect 24421 -4574 24559 -4540
rect 24421 -4590 24593 -4574
rect 24627 -4549 24658 -4515
rect 24696 -4540 24786 -4515
rect 24696 -4549 24730 -4540
rect 24627 -4574 24730 -4549
rect 24764 -4574 24786 -4540
rect 24421 -4670 24471 -4590
rect 24627 -4594 24786 -4574
rect 24820 -4525 24866 -4430
rect 24820 -4534 24832 -4525
rect 24854 -4568 24866 -4559
rect 24627 -4630 24669 -4594
rect 24820 -4628 24866 -4568
rect 24618 -4646 24669 -4630
rect 24421 -4704 24437 -4670
rect 24421 -4720 24471 -4704
rect 24534 -4676 24568 -4653
rect 24317 -4734 24383 -4726
rect 24534 -4772 24568 -4710
rect 24652 -4680 24669 -4646
rect 24618 -4736 24669 -4680
rect 24716 -4662 24866 -4628
rect 24716 -4670 24767 -4662
rect 24716 -4704 24733 -4670
rect 24901 -4670 24935 -4432
rect 24969 -4456 25034 -4299
rect 25068 -4304 25118 -4262
rect 25068 -4338 25084 -4304
rect 25068 -4354 25118 -4338
rect 25152 -4312 25202 -4296
rect 25152 -4346 25168 -4312
rect 25152 -4362 25202 -4346
rect 25245 -4306 25381 -4296
rect 25245 -4340 25261 -4306
rect 25295 -4340 25381 -4306
rect 25496 -4314 25562 -4262
rect 25689 -4304 25763 -4262
rect 25245 -4362 25381 -4340
rect 25152 -4388 25186 -4362
rect 25107 -4422 25186 -4388
rect 25220 -4398 25313 -4396
rect 24981 -4479 25073 -4456
rect 24981 -4513 25039 -4479
rect 24981 -4614 25073 -4513
rect 24981 -4648 25005 -4614
rect 25043 -4648 25073 -4614
rect 24981 -4666 25073 -4648
rect 24716 -4720 24767 -4704
rect 24801 -4730 24817 -4696
rect 24851 -4730 24867 -4696
rect 25107 -4694 25141 -4422
rect 25220 -4424 25279 -4398
rect 25254 -4432 25279 -4424
rect 25254 -4458 25313 -4432
rect 25220 -4474 25313 -4458
rect 25175 -4534 25245 -4512
rect 25175 -4568 25187 -4534
rect 25221 -4568 25245 -4534
rect 25175 -4586 25245 -4568
rect 25175 -4620 25198 -4586
rect 25232 -4620 25245 -4586
rect 25175 -4636 25245 -4620
rect 25279 -4592 25313 -4474
rect 25347 -4518 25381 -4362
rect 25415 -4330 25449 -4314
rect 25496 -4348 25512 -4314
rect 25546 -4348 25562 -4314
rect 25596 -4330 25630 -4314
rect 25415 -4382 25449 -4364
rect 25689 -4338 25709 -4304
rect 25743 -4338 25763 -4304
rect 25689 -4354 25763 -4338
rect 25797 -4312 25831 -4296
rect 25596 -4382 25630 -4364
rect 25415 -4416 25630 -4382
rect 25797 -4388 25831 -4346
rect 25878 -4305 26052 -4296
rect 25878 -4339 25894 -4305
rect 25928 -4339 26052 -4305
rect 25878 -4364 26052 -4339
rect 26086 -4304 26136 -4262
rect 26120 -4338 26136 -4304
rect 26240 -4304 26384 -4262
rect 26086 -4354 26136 -4338
rect 26170 -4330 26204 -4314
rect 25719 -4422 25831 -4388
rect 25719 -4450 25753 -4422
rect 25453 -4484 25469 -4450
rect 25503 -4484 25753 -4450
rect 25892 -4432 25903 -4398
rect 25937 -4424 25984 -4398
rect 25892 -4456 25934 -4432
rect 25347 -4538 25685 -4518
rect 25347 -4552 25651 -4538
rect 25279 -4626 25300 -4592
rect 25334 -4626 25350 -4592
rect 25279 -4636 25350 -4626
rect 25384 -4694 25418 -4552
rect 25459 -4602 25555 -4586
rect 25493 -4636 25531 -4602
rect 25589 -4620 25617 -4586
rect 25651 -4588 25685 -4572
rect 25565 -4636 25617 -4620
rect 25719 -4622 25753 -4484
rect 24901 -4720 24935 -4704
rect 24801 -4772 24867 -4730
rect 25007 -4734 25023 -4700
rect 25057 -4734 25073 -4700
rect 25107 -4728 25156 -4694
rect 25190 -4728 25206 -4694
rect 25247 -4728 25263 -4694
rect 25297 -4728 25418 -4694
rect 25593 -4696 25659 -4680
rect 25007 -4772 25073 -4734
rect 25593 -4730 25609 -4696
rect 25643 -4730 25659 -4696
rect 25593 -4772 25659 -4730
rect 25701 -4700 25753 -4622
rect 25791 -4458 25934 -4456
rect 25968 -4458 25984 -4424
rect 26018 -4440 26052 -4364
rect 26240 -4338 26256 -4304
rect 26290 -4338 26334 -4304
rect 26368 -4338 26384 -4304
rect 26418 -4312 26499 -4296
rect 26650 -4304 26684 -4262
rect 26170 -4372 26204 -4364
rect 26452 -4346 26499 -4312
rect 26170 -4406 26330 -4372
rect 25791 -4490 25926 -4458
rect 26018 -4474 26212 -4440
rect 26246 -4474 26262 -4440
rect 25791 -4598 25833 -4490
rect 26018 -4492 26052 -4474
rect 25791 -4632 25799 -4598
rect 25791 -4648 25833 -4632
rect 25867 -4534 25937 -4524
rect 25867 -4550 25903 -4534
rect 25867 -4584 25895 -4550
rect 25929 -4584 25937 -4568
rect 25867 -4648 25937 -4584
rect 25971 -4526 26052 -4492
rect 25971 -4682 26005 -4526
rect 26119 -4539 26227 -4508
rect 26296 -4524 26330 -4406
rect 26418 -4380 26499 -4346
rect 26452 -4414 26499 -4380
rect 26418 -4448 26499 -4414
rect 26452 -4482 26499 -4448
rect 26418 -4498 26499 -4482
rect 26296 -4530 26385 -4524
rect 26153 -4548 26227 -4539
rect 26039 -4576 26083 -4560
rect 26073 -4610 26083 -4576
rect 26119 -4582 26135 -4573
rect 26169 -4582 26227 -4548
rect 26039 -4616 26083 -4610
rect 26179 -4602 26227 -4582
rect 26039 -4650 26145 -4616
rect 25815 -4696 26005 -4682
rect 25701 -4734 25721 -4700
rect 25755 -4734 25771 -4700
rect 25815 -4730 25831 -4696
rect 25865 -4730 26005 -4696
rect 25815 -4738 26005 -4730
rect 26039 -4700 26077 -4684
rect 26039 -4734 26043 -4700
rect 26111 -4696 26145 -4650
rect 26213 -4636 26227 -4602
rect 26179 -4662 26227 -4636
rect 26261 -4540 26385 -4530
rect 26261 -4574 26335 -4540
rect 26369 -4574 26385 -4540
rect 26261 -4590 26385 -4574
rect 26261 -4625 26326 -4590
rect 26433 -4624 26499 -4498
rect 26261 -4680 26325 -4625
rect 26111 -4714 26261 -4696
rect 26295 -4714 26325 -4680
rect 26111 -4730 26325 -4714
rect 26365 -4657 26399 -4635
rect 26039 -4772 26077 -4734
rect 26365 -4772 26399 -4691
rect 26433 -4658 26449 -4624
rect 26483 -4658 26499 -4624
rect 26433 -4692 26499 -4658
rect 26433 -4726 26449 -4692
rect 26483 -4726 26499 -4692
rect 26537 -4338 26553 -4304
rect 26587 -4338 26603 -4304
rect 26537 -4372 26603 -4338
rect 26537 -4406 26553 -4372
rect 26587 -4406 26603 -4372
rect 26537 -4524 26603 -4406
rect 26832 -4312 26883 -4296
rect 26650 -4372 26684 -4338
rect 26650 -4440 26684 -4406
rect 26650 -4490 26684 -4474
rect 26734 -4340 26785 -4324
rect 26768 -4374 26785 -4340
rect 26734 -4408 26785 -4374
rect 26768 -4442 26785 -4408
rect 26832 -4346 26849 -4312
rect 26832 -4380 26883 -4346
rect 26917 -4328 26983 -4262
rect 26917 -4362 26933 -4328
rect 26967 -4362 26983 -4328
rect 27017 -4312 27051 -4296
rect 26832 -4414 26849 -4380
rect 27017 -4380 27051 -4346
rect 26883 -4414 26982 -4396
rect 26832 -4430 26982 -4414
rect 26734 -4464 26785 -4442
rect 26734 -4500 26902 -4464
rect 26743 -4515 26902 -4500
rect 26537 -4540 26709 -4524
rect 26537 -4574 26675 -4540
rect 26537 -4590 26709 -4574
rect 26743 -4549 26774 -4515
rect 26812 -4540 26902 -4515
rect 26812 -4549 26846 -4540
rect 26743 -4574 26846 -4549
rect 26880 -4574 26902 -4540
rect 26537 -4670 26587 -4590
rect 26743 -4594 26902 -4574
rect 26936 -4525 26982 -4430
rect 26936 -4534 26948 -4525
rect 26970 -4568 26982 -4559
rect 26743 -4630 26785 -4594
rect 26936 -4628 26982 -4568
rect 26734 -4646 26785 -4630
rect 26537 -4704 26553 -4670
rect 26537 -4720 26587 -4704
rect 26650 -4676 26684 -4653
rect 26433 -4734 26499 -4726
rect 26650 -4772 26684 -4710
rect 26768 -4680 26785 -4646
rect 26734 -4736 26785 -4680
rect 26832 -4662 26982 -4628
rect 26832 -4670 26883 -4662
rect 26832 -4704 26849 -4670
rect 27017 -4670 27051 -4432
rect 27085 -4456 27150 -4299
rect 27184 -4304 27234 -4262
rect 27184 -4338 27200 -4304
rect 27184 -4354 27234 -4338
rect 27268 -4312 27318 -4296
rect 27268 -4346 27284 -4312
rect 27268 -4362 27318 -4346
rect 27361 -4306 27497 -4296
rect 27361 -4340 27377 -4306
rect 27411 -4340 27497 -4306
rect 27612 -4314 27678 -4262
rect 27805 -4304 27879 -4262
rect 27361 -4362 27497 -4340
rect 27268 -4388 27302 -4362
rect 27223 -4422 27302 -4388
rect 27336 -4398 27429 -4396
rect 27097 -4479 27189 -4456
rect 27097 -4513 27155 -4479
rect 27097 -4614 27189 -4513
rect 27097 -4648 27121 -4614
rect 27159 -4648 27189 -4614
rect 27097 -4666 27189 -4648
rect 26832 -4720 26883 -4704
rect 26917 -4730 26933 -4696
rect 26967 -4730 26983 -4696
rect 27223 -4694 27257 -4422
rect 27336 -4424 27395 -4398
rect 27370 -4432 27395 -4424
rect 27370 -4458 27429 -4432
rect 27336 -4474 27429 -4458
rect 27291 -4534 27361 -4512
rect 27291 -4568 27303 -4534
rect 27337 -4568 27361 -4534
rect 27291 -4586 27361 -4568
rect 27291 -4620 27314 -4586
rect 27348 -4620 27361 -4586
rect 27291 -4636 27361 -4620
rect 27395 -4592 27429 -4474
rect 27463 -4518 27497 -4362
rect 27531 -4330 27565 -4314
rect 27612 -4348 27628 -4314
rect 27662 -4348 27678 -4314
rect 27712 -4330 27746 -4314
rect 27531 -4382 27565 -4364
rect 27805 -4338 27825 -4304
rect 27859 -4338 27879 -4304
rect 27805 -4354 27879 -4338
rect 27913 -4312 27947 -4296
rect 27712 -4382 27746 -4364
rect 27531 -4416 27746 -4382
rect 27913 -4388 27947 -4346
rect 27994 -4305 28168 -4296
rect 27994 -4339 28010 -4305
rect 28044 -4339 28168 -4305
rect 27994 -4364 28168 -4339
rect 28202 -4304 28252 -4262
rect 28236 -4338 28252 -4304
rect 28356 -4304 28500 -4262
rect 28202 -4354 28252 -4338
rect 28286 -4330 28320 -4314
rect 27835 -4422 27947 -4388
rect 27835 -4450 27869 -4422
rect 27569 -4484 27585 -4450
rect 27619 -4484 27869 -4450
rect 28008 -4432 28019 -4398
rect 28053 -4424 28100 -4398
rect 28008 -4456 28050 -4432
rect 27463 -4538 27801 -4518
rect 27463 -4552 27767 -4538
rect 27395 -4626 27416 -4592
rect 27450 -4626 27466 -4592
rect 27395 -4636 27466 -4626
rect 27500 -4694 27534 -4552
rect 27575 -4602 27671 -4586
rect 27609 -4636 27647 -4602
rect 27705 -4620 27733 -4586
rect 27767 -4588 27801 -4572
rect 27681 -4636 27733 -4620
rect 27835 -4622 27869 -4484
rect 27017 -4720 27051 -4704
rect 26917 -4772 26983 -4730
rect 27123 -4734 27139 -4700
rect 27173 -4734 27189 -4700
rect 27223 -4728 27272 -4694
rect 27306 -4728 27322 -4694
rect 27363 -4728 27379 -4694
rect 27413 -4728 27534 -4694
rect 27709 -4696 27775 -4680
rect 27123 -4772 27189 -4734
rect 27709 -4730 27725 -4696
rect 27759 -4730 27775 -4696
rect 27709 -4772 27775 -4730
rect 27817 -4700 27869 -4622
rect 27907 -4458 28050 -4456
rect 28084 -4458 28100 -4424
rect 28134 -4440 28168 -4364
rect 28356 -4338 28372 -4304
rect 28406 -4338 28450 -4304
rect 28484 -4338 28500 -4304
rect 28534 -4312 28615 -4296
rect 28766 -4304 28800 -4262
rect 28286 -4372 28320 -4364
rect 28568 -4346 28615 -4312
rect 28286 -4406 28446 -4372
rect 27907 -4490 28042 -4458
rect 28134 -4474 28328 -4440
rect 28362 -4474 28378 -4440
rect 27907 -4598 27949 -4490
rect 28134 -4492 28168 -4474
rect 27907 -4632 27915 -4598
rect 27907 -4648 27949 -4632
rect 27983 -4534 28053 -4524
rect 27983 -4550 28019 -4534
rect 27983 -4584 28011 -4550
rect 28045 -4584 28053 -4568
rect 27983 -4648 28053 -4584
rect 28087 -4526 28168 -4492
rect 28087 -4682 28121 -4526
rect 28235 -4539 28343 -4508
rect 28412 -4524 28446 -4406
rect 28534 -4380 28615 -4346
rect 28568 -4414 28615 -4380
rect 28534 -4448 28615 -4414
rect 28568 -4482 28615 -4448
rect 28534 -4498 28615 -4482
rect 28412 -4530 28501 -4524
rect 28269 -4548 28343 -4539
rect 28155 -4576 28199 -4560
rect 28189 -4610 28199 -4576
rect 28235 -4582 28251 -4573
rect 28285 -4582 28343 -4548
rect 28155 -4616 28199 -4610
rect 28295 -4602 28343 -4582
rect 28155 -4650 28261 -4616
rect 27931 -4696 28121 -4682
rect 27817 -4734 27837 -4700
rect 27871 -4734 27887 -4700
rect 27931 -4730 27947 -4696
rect 27981 -4730 28121 -4696
rect 27931 -4738 28121 -4730
rect 28155 -4700 28193 -4684
rect 28155 -4734 28159 -4700
rect 28227 -4696 28261 -4650
rect 28329 -4636 28343 -4602
rect 28295 -4662 28343 -4636
rect 28377 -4540 28501 -4530
rect 28377 -4574 28451 -4540
rect 28485 -4574 28501 -4540
rect 28377 -4590 28501 -4574
rect 28377 -4625 28442 -4590
rect 28549 -4624 28615 -4498
rect 28377 -4680 28441 -4625
rect 28227 -4714 28377 -4696
rect 28411 -4714 28441 -4680
rect 28227 -4730 28441 -4714
rect 28481 -4657 28515 -4635
rect 28155 -4772 28193 -4734
rect 28481 -4772 28515 -4691
rect 28549 -4658 28565 -4624
rect 28599 -4658 28615 -4624
rect 28549 -4692 28615 -4658
rect 28549 -4726 28565 -4692
rect 28599 -4726 28615 -4692
rect 28653 -4338 28669 -4304
rect 28703 -4338 28719 -4304
rect 28653 -4372 28719 -4338
rect 28653 -4406 28669 -4372
rect 28703 -4406 28719 -4372
rect 28653 -4524 28719 -4406
rect 28948 -4312 28999 -4296
rect 28766 -4372 28800 -4338
rect 28766 -4440 28800 -4406
rect 28766 -4490 28800 -4474
rect 28850 -4340 28901 -4324
rect 28884 -4374 28901 -4340
rect 28850 -4408 28901 -4374
rect 28884 -4442 28901 -4408
rect 28948 -4346 28965 -4312
rect 28948 -4380 28999 -4346
rect 29033 -4328 29099 -4262
rect 29033 -4362 29049 -4328
rect 29083 -4362 29099 -4328
rect 29133 -4312 29167 -4296
rect 28948 -4414 28965 -4380
rect 29133 -4380 29167 -4346
rect 28999 -4414 29098 -4396
rect 28948 -4430 29098 -4414
rect 28850 -4464 28901 -4442
rect 28850 -4500 29018 -4464
rect 28859 -4515 29018 -4500
rect 28653 -4540 28825 -4524
rect 28653 -4574 28791 -4540
rect 28653 -4590 28825 -4574
rect 28859 -4549 28890 -4515
rect 28928 -4540 29018 -4515
rect 28928 -4549 28962 -4540
rect 28859 -4574 28962 -4549
rect 28996 -4574 29018 -4540
rect 28653 -4670 28703 -4590
rect 28859 -4594 29018 -4574
rect 29052 -4525 29098 -4430
rect 29052 -4534 29064 -4525
rect 29086 -4568 29098 -4559
rect 28859 -4630 28901 -4594
rect 29052 -4628 29098 -4568
rect 28850 -4646 28901 -4630
rect 28653 -4704 28669 -4670
rect 28653 -4720 28703 -4704
rect 28766 -4676 28800 -4653
rect 28549 -4734 28615 -4726
rect 28766 -4772 28800 -4710
rect 28884 -4680 28901 -4646
rect 28850 -4736 28901 -4680
rect 28948 -4662 29098 -4628
rect 28948 -4670 28999 -4662
rect 28948 -4704 28965 -4670
rect 29133 -4670 29167 -4432
rect 29201 -4456 29266 -4299
rect 29300 -4304 29350 -4262
rect 29300 -4338 29316 -4304
rect 29300 -4354 29350 -4338
rect 29384 -4312 29434 -4296
rect 29384 -4346 29400 -4312
rect 29384 -4362 29434 -4346
rect 29477 -4306 29613 -4296
rect 29477 -4340 29493 -4306
rect 29527 -4340 29613 -4306
rect 29728 -4314 29794 -4262
rect 29921 -4304 29995 -4262
rect 29477 -4362 29613 -4340
rect 29384 -4388 29418 -4362
rect 29339 -4422 29418 -4388
rect 29452 -4398 29545 -4396
rect 29213 -4479 29305 -4456
rect 29213 -4513 29271 -4479
rect 29213 -4614 29305 -4513
rect 29213 -4648 29237 -4614
rect 29275 -4648 29305 -4614
rect 29213 -4666 29305 -4648
rect 28948 -4720 28999 -4704
rect 29033 -4730 29049 -4696
rect 29083 -4730 29099 -4696
rect 29339 -4694 29373 -4422
rect 29452 -4424 29511 -4398
rect 29486 -4432 29511 -4424
rect 29486 -4458 29545 -4432
rect 29452 -4474 29545 -4458
rect 29407 -4534 29477 -4512
rect 29407 -4568 29419 -4534
rect 29453 -4568 29477 -4534
rect 29407 -4586 29477 -4568
rect 29407 -4620 29430 -4586
rect 29464 -4620 29477 -4586
rect 29407 -4636 29477 -4620
rect 29511 -4592 29545 -4474
rect 29579 -4518 29613 -4362
rect 29647 -4330 29681 -4314
rect 29728 -4348 29744 -4314
rect 29778 -4348 29794 -4314
rect 29828 -4330 29862 -4314
rect 29647 -4382 29681 -4364
rect 29921 -4338 29941 -4304
rect 29975 -4338 29995 -4304
rect 29921 -4354 29995 -4338
rect 30029 -4312 30063 -4296
rect 29828 -4382 29862 -4364
rect 29647 -4416 29862 -4382
rect 30029 -4388 30063 -4346
rect 30110 -4305 30284 -4296
rect 30110 -4339 30126 -4305
rect 30160 -4339 30284 -4305
rect 30110 -4364 30284 -4339
rect 30318 -4304 30368 -4262
rect 30352 -4338 30368 -4304
rect 30472 -4304 30616 -4262
rect 30318 -4354 30368 -4338
rect 30402 -4330 30436 -4314
rect 29951 -4422 30063 -4388
rect 29951 -4450 29985 -4422
rect 29685 -4484 29701 -4450
rect 29735 -4484 29985 -4450
rect 30124 -4432 30135 -4398
rect 30169 -4424 30216 -4398
rect 30124 -4456 30166 -4432
rect 29579 -4538 29917 -4518
rect 29579 -4552 29883 -4538
rect 29511 -4626 29532 -4592
rect 29566 -4626 29582 -4592
rect 29511 -4636 29582 -4626
rect 29616 -4694 29650 -4552
rect 29691 -4602 29787 -4586
rect 29725 -4636 29763 -4602
rect 29821 -4620 29849 -4586
rect 29883 -4588 29917 -4572
rect 29797 -4636 29849 -4620
rect 29951 -4622 29985 -4484
rect 29133 -4720 29167 -4704
rect 29033 -4772 29099 -4730
rect 29239 -4734 29255 -4700
rect 29289 -4734 29305 -4700
rect 29339 -4728 29388 -4694
rect 29422 -4728 29438 -4694
rect 29479 -4728 29495 -4694
rect 29529 -4728 29650 -4694
rect 29825 -4696 29891 -4680
rect 29239 -4772 29305 -4734
rect 29825 -4730 29841 -4696
rect 29875 -4730 29891 -4696
rect 29825 -4772 29891 -4730
rect 29933 -4700 29985 -4622
rect 30023 -4458 30166 -4456
rect 30200 -4458 30216 -4424
rect 30250 -4440 30284 -4364
rect 30472 -4338 30488 -4304
rect 30522 -4338 30566 -4304
rect 30600 -4338 30616 -4304
rect 30650 -4312 30731 -4296
rect 30882 -4304 30916 -4262
rect 30402 -4372 30436 -4364
rect 30684 -4346 30731 -4312
rect 30402 -4406 30562 -4372
rect 30023 -4490 30158 -4458
rect 30250 -4474 30444 -4440
rect 30478 -4474 30494 -4440
rect 30023 -4598 30065 -4490
rect 30250 -4492 30284 -4474
rect 30023 -4632 30031 -4598
rect 30023 -4648 30065 -4632
rect 30099 -4534 30169 -4524
rect 30099 -4550 30135 -4534
rect 30099 -4584 30127 -4550
rect 30161 -4584 30169 -4568
rect 30099 -4648 30169 -4584
rect 30203 -4526 30284 -4492
rect 30203 -4682 30237 -4526
rect 30351 -4539 30459 -4508
rect 30528 -4524 30562 -4406
rect 30650 -4380 30731 -4346
rect 30684 -4414 30731 -4380
rect 30650 -4448 30731 -4414
rect 30684 -4482 30731 -4448
rect 30650 -4498 30731 -4482
rect 30528 -4530 30617 -4524
rect 30385 -4548 30459 -4539
rect 30271 -4576 30315 -4560
rect 30305 -4610 30315 -4576
rect 30351 -4582 30367 -4573
rect 30401 -4582 30459 -4548
rect 30271 -4616 30315 -4610
rect 30411 -4602 30459 -4582
rect 30271 -4650 30377 -4616
rect 30047 -4696 30237 -4682
rect 29933 -4734 29953 -4700
rect 29987 -4734 30003 -4700
rect 30047 -4730 30063 -4696
rect 30097 -4730 30237 -4696
rect 30047 -4738 30237 -4730
rect 30271 -4700 30309 -4684
rect 30271 -4734 30275 -4700
rect 30343 -4696 30377 -4650
rect 30445 -4636 30459 -4602
rect 30411 -4662 30459 -4636
rect 30493 -4540 30617 -4530
rect 30493 -4574 30567 -4540
rect 30601 -4574 30617 -4540
rect 30493 -4590 30617 -4574
rect 30493 -4625 30558 -4590
rect 30665 -4624 30731 -4498
rect 30493 -4680 30557 -4625
rect 30343 -4714 30493 -4696
rect 30527 -4714 30557 -4680
rect 30343 -4730 30557 -4714
rect 30597 -4657 30631 -4635
rect 30271 -4772 30309 -4734
rect 30597 -4772 30631 -4691
rect 30665 -4658 30681 -4624
rect 30715 -4658 30731 -4624
rect 30665 -4692 30731 -4658
rect 30665 -4726 30681 -4692
rect 30715 -4726 30731 -4692
rect 30769 -4338 30785 -4304
rect 30819 -4338 30835 -4304
rect 30769 -4372 30835 -4338
rect 30769 -4406 30785 -4372
rect 30819 -4406 30835 -4372
rect 30769 -4524 30835 -4406
rect 31064 -4312 31115 -4296
rect 30882 -4372 30916 -4338
rect 30882 -4440 30916 -4406
rect 30882 -4490 30916 -4474
rect 30966 -4340 31017 -4324
rect 31000 -4374 31017 -4340
rect 30966 -4408 31017 -4374
rect 31000 -4442 31017 -4408
rect 31064 -4346 31081 -4312
rect 31064 -4380 31115 -4346
rect 31149 -4328 31215 -4262
rect 31149 -4362 31165 -4328
rect 31199 -4362 31215 -4328
rect 31249 -4312 31283 -4296
rect 31064 -4414 31081 -4380
rect 31249 -4380 31283 -4346
rect 31115 -4414 31214 -4396
rect 31064 -4430 31214 -4414
rect 30966 -4464 31017 -4442
rect 30966 -4500 31134 -4464
rect 30975 -4515 31134 -4500
rect 30769 -4540 30941 -4524
rect 30769 -4574 30907 -4540
rect 30769 -4590 30941 -4574
rect 30975 -4549 31006 -4515
rect 31044 -4540 31134 -4515
rect 31044 -4549 31078 -4540
rect 30975 -4574 31078 -4549
rect 31112 -4574 31134 -4540
rect 30769 -4670 30819 -4590
rect 30975 -4594 31134 -4574
rect 31168 -4525 31214 -4430
rect 31168 -4534 31180 -4525
rect 31202 -4568 31214 -4559
rect 30975 -4630 31017 -4594
rect 31168 -4628 31214 -4568
rect 30966 -4646 31017 -4630
rect 30769 -4704 30785 -4670
rect 30769 -4720 30819 -4704
rect 30882 -4676 30916 -4653
rect 30665 -4734 30731 -4726
rect 30882 -4772 30916 -4710
rect 31000 -4680 31017 -4646
rect 30966 -4736 31017 -4680
rect 31064 -4662 31214 -4628
rect 31064 -4670 31115 -4662
rect 31064 -4704 31081 -4670
rect 31249 -4670 31283 -4432
rect 31317 -4456 31382 -4299
rect 31416 -4304 31466 -4262
rect 31416 -4338 31432 -4304
rect 31416 -4354 31466 -4338
rect 31500 -4312 31550 -4296
rect 31500 -4346 31516 -4312
rect 31500 -4362 31550 -4346
rect 31593 -4306 31729 -4296
rect 31593 -4340 31609 -4306
rect 31643 -4340 31729 -4306
rect 31844 -4314 31910 -4262
rect 32037 -4304 32111 -4262
rect 31593 -4362 31729 -4340
rect 31500 -4388 31534 -4362
rect 31455 -4422 31534 -4388
rect 31568 -4398 31661 -4396
rect 31329 -4479 31421 -4456
rect 31329 -4513 31387 -4479
rect 31329 -4614 31421 -4513
rect 31329 -4648 31353 -4614
rect 31391 -4648 31421 -4614
rect 31329 -4666 31421 -4648
rect 31064 -4720 31115 -4704
rect 31149 -4730 31165 -4696
rect 31199 -4730 31215 -4696
rect 31455 -4694 31489 -4422
rect 31568 -4424 31627 -4398
rect 31602 -4432 31627 -4424
rect 31602 -4458 31661 -4432
rect 31568 -4474 31661 -4458
rect 31523 -4534 31593 -4512
rect 31523 -4568 31535 -4534
rect 31569 -4568 31593 -4534
rect 31523 -4586 31593 -4568
rect 31523 -4620 31546 -4586
rect 31580 -4620 31593 -4586
rect 31523 -4636 31593 -4620
rect 31627 -4592 31661 -4474
rect 31695 -4518 31729 -4362
rect 31763 -4330 31797 -4314
rect 31844 -4348 31860 -4314
rect 31894 -4348 31910 -4314
rect 31944 -4330 31978 -4314
rect 31763 -4382 31797 -4364
rect 32037 -4338 32057 -4304
rect 32091 -4338 32111 -4304
rect 32037 -4354 32111 -4338
rect 32145 -4312 32179 -4296
rect 31944 -4382 31978 -4364
rect 31763 -4416 31978 -4382
rect 32145 -4388 32179 -4346
rect 32226 -4305 32400 -4296
rect 32226 -4339 32242 -4305
rect 32276 -4339 32400 -4305
rect 32226 -4364 32400 -4339
rect 32434 -4304 32484 -4262
rect 32468 -4338 32484 -4304
rect 32588 -4304 32732 -4262
rect 32434 -4354 32484 -4338
rect 32518 -4330 32552 -4314
rect 32067 -4422 32179 -4388
rect 32067 -4450 32101 -4422
rect 31801 -4484 31817 -4450
rect 31851 -4484 32101 -4450
rect 32240 -4432 32251 -4398
rect 32285 -4424 32332 -4398
rect 32240 -4456 32282 -4432
rect 31695 -4538 32033 -4518
rect 31695 -4552 31999 -4538
rect 31627 -4626 31648 -4592
rect 31682 -4626 31698 -4592
rect 31627 -4636 31698 -4626
rect 31732 -4694 31766 -4552
rect 31807 -4602 31903 -4586
rect 31841 -4636 31879 -4602
rect 31937 -4620 31965 -4586
rect 31999 -4588 32033 -4572
rect 31913 -4636 31965 -4620
rect 32067 -4622 32101 -4484
rect 31249 -4720 31283 -4704
rect 31149 -4772 31215 -4730
rect 31355 -4734 31371 -4700
rect 31405 -4734 31421 -4700
rect 31455 -4728 31504 -4694
rect 31538 -4728 31554 -4694
rect 31595 -4728 31611 -4694
rect 31645 -4728 31766 -4694
rect 31941 -4696 32007 -4680
rect 31355 -4772 31421 -4734
rect 31941 -4730 31957 -4696
rect 31991 -4730 32007 -4696
rect 31941 -4772 32007 -4730
rect 32049 -4700 32101 -4622
rect 32139 -4458 32282 -4456
rect 32316 -4458 32332 -4424
rect 32366 -4440 32400 -4364
rect 32588 -4338 32604 -4304
rect 32638 -4338 32682 -4304
rect 32716 -4338 32732 -4304
rect 32766 -4312 32847 -4296
rect 32998 -4304 33032 -4262
rect 32518 -4372 32552 -4364
rect 32800 -4346 32847 -4312
rect 32518 -4406 32678 -4372
rect 32139 -4490 32274 -4458
rect 32366 -4474 32560 -4440
rect 32594 -4474 32610 -4440
rect 32139 -4598 32181 -4490
rect 32366 -4492 32400 -4474
rect 32139 -4632 32147 -4598
rect 32139 -4648 32181 -4632
rect 32215 -4534 32285 -4524
rect 32215 -4550 32251 -4534
rect 32215 -4584 32243 -4550
rect 32277 -4584 32285 -4568
rect 32215 -4648 32285 -4584
rect 32319 -4526 32400 -4492
rect 32319 -4682 32353 -4526
rect 32467 -4539 32575 -4508
rect 32644 -4524 32678 -4406
rect 32766 -4380 32847 -4346
rect 32800 -4414 32847 -4380
rect 32766 -4448 32847 -4414
rect 32800 -4482 32847 -4448
rect 32766 -4498 32847 -4482
rect 32644 -4530 32733 -4524
rect 32501 -4548 32575 -4539
rect 32387 -4576 32431 -4560
rect 32421 -4610 32431 -4576
rect 32467 -4582 32483 -4573
rect 32517 -4582 32575 -4548
rect 32387 -4616 32431 -4610
rect 32527 -4602 32575 -4582
rect 32387 -4650 32493 -4616
rect 32163 -4696 32353 -4682
rect 32049 -4734 32069 -4700
rect 32103 -4734 32119 -4700
rect 32163 -4730 32179 -4696
rect 32213 -4730 32353 -4696
rect 32163 -4738 32353 -4730
rect 32387 -4700 32425 -4684
rect 32387 -4734 32391 -4700
rect 32459 -4696 32493 -4650
rect 32561 -4636 32575 -4602
rect 32527 -4662 32575 -4636
rect 32609 -4540 32733 -4530
rect 32609 -4574 32683 -4540
rect 32717 -4574 32733 -4540
rect 32609 -4590 32733 -4574
rect 32609 -4625 32674 -4590
rect 32781 -4624 32847 -4498
rect 32609 -4680 32673 -4625
rect 32459 -4714 32609 -4696
rect 32643 -4714 32673 -4680
rect 32459 -4730 32673 -4714
rect 32713 -4657 32747 -4635
rect 32387 -4772 32425 -4734
rect 32713 -4772 32747 -4691
rect 32781 -4658 32797 -4624
rect 32831 -4658 32847 -4624
rect 32781 -4692 32847 -4658
rect 32781 -4726 32797 -4692
rect 32831 -4726 32847 -4692
rect 32885 -4338 32901 -4304
rect 32935 -4338 32951 -4304
rect 32885 -4372 32951 -4338
rect 32885 -4406 32901 -4372
rect 32935 -4406 32951 -4372
rect 32885 -4524 32951 -4406
rect 32998 -4372 33032 -4338
rect 32998 -4440 33032 -4406
rect 32998 -4490 33032 -4474
rect 33082 -4340 33133 -4324
rect 33116 -4374 33133 -4340
rect 33082 -4408 33133 -4374
rect 33116 -4442 33133 -4408
rect 33082 -4464 33133 -4442
rect 33082 -4500 33162 -4464
rect 33091 -4515 33162 -4500
rect 32885 -4540 33057 -4524
rect 32885 -4574 33023 -4540
rect 32885 -4590 33057 -4574
rect 33091 -4549 33122 -4515
rect 33160 -4549 33162 -4515
rect 32885 -4670 32935 -4590
rect 33091 -4594 33162 -4549
rect 33091 -4630 33133 -4594
rect 33082 -4646 33133 -4630
rect 32885 -4704 32901 -4670
rect 32885 -4720 32935 -4704
rect 32998 -4676 33032 -4653
rect 32781 -4734 32847 -4726
rect 32998 -4772 33032 -4710
rect 33116 -4680 33133 -4646
rect 33082 -4736 33133 -4680
rect -9158 -4830 -9129 -4772
rect -9095 -4830 -9037 -4772
rect -9003 -4830 -8945 -4772
rect -8911 -4830 -8853 -4772
rect -8819 -4830 -8761 -4772
rect -8727 -4830 -8669 -4772
rect -8635 -4830 -8577 -4772
rect -8543 -4830 -8485 -4772
rect -8451 -4830 -8393 -4772
rect -8359 -4830 -8301 -4772
rect -8267 -4830 -8209 -4772
rect -8175 -4830 -8117 -4772
rect -8083 -4830 -8025 -4772
rect -7991 -4830 -7933 -4772
rect -7899 -4830 -7841 -4772
rect -7807 -4830 -7749 -4772
rect -7715 -4830 -7657 -4772
rect -7623 -4830 -7565 -4772
rect -7531 -4830 -7473 -4772
rect -7439 -4830 -7381 -4772
rect -7347 -4830 -7289 -4772
rect -7255 -4830 -7197 -4772
rect -7163 -4830 -7105 -4772
rect -7071 -4830 -7013 -4772
rect -6979 -4830 -6921 -4772
rect -6887 -4830 -6829 -4772
rect -6795 -4830 -6737 -4772
rect -6703 -4830 -6645 -4772
rect -6611 -4830 -6553 -4772
rect -6519 -4830 -6461 -4772
rect -6427 -4830 -6369 -4772
rect -6335 -4830 -6277 -4772
rect -6243 -4830 -6185 -4772
rect -6151 -4830 -6093 -4772
rect -6059 -4830 -6001 -4772
rect -5967 -4830 -5909 -4772
rect -5875 -4830 -5817 -4772
rect -5783 -4830 -5725 -4772
rect -5691 -4830 -5633 -4772
rect -5599 -4830 -5541 -4772
rect -5507 -4830 -5449 -4772
rect -5415 -4830 -5357 -4772
rect -5323 -4830 -5265 -4772
rect -5231 -4830 -5173 -4772
rect -5139 -4830 -5081 -4772
rect -5047 -4830 -4989 -4772
rect -4955 -4830 -4897 -4772
rect -4863 -4830 -4805 -4772
rect -4771 -4830 -4713 -4772
rect -4679 -4830 -4621 -4772
rect -4587 -4830 -4529 -4772
rect -4495 -4830 -4437 -4772
rect -4403 -4830 -4345 -4772
rect -4311 -4830 -4253 -4772
rect -4219 -4830 -4161 -4772
rect -4127 -4830 -4069 -4772
rect -4035 -4830 -3977 -4772
rect -3943 -4830 -3885 -4772
rect -3851 -4830 -3793 -4772
rect -3759 -4830 -3701 -4772
rect -3667 -4830 -3609 -4772
rect -3575 -4830 -3517 -4772
rect -3483 -4830 -3425 -4772
rect -3391 -4830 -3333 -4772
rect -3299 -4830 -3241 -4772
rect -3207 -4830 -3149 -4772
rect -3115 -4830 -3057 -4772
rect -3023 -4830 -2965 -4772
rect -2931 -4830 -2873 -4772
rect -2839 -4830 -2781 -4772
rect -2747 -4830 -2689 -4772
rect -2655 -4830 -2597 -4772
rect -2563 -4830 -2505 -4772
rect -2471 -4830 -2413 -4772
rect -2379 -4830 -2321 -4772
rect -2287 -4830 -2229 -4772
rect -2195 -4830 -2137 -4772
rect -2103 -4830 -2045 -4772
rect -2011 -4830 -1953 -4772
rect -1919 -4830 -1861 -4772
rect -1827 -4830 -1769 -4772
rect -1735 -4830 -1677 -4772
rect -1643 -4830 -1585 -4772
rect -1551 -4830 -1493 -4772
rect -1459 -4830 -1401 -4772
rect -1367 -4830 -1309 -4772
rect -1275 -4830 -1217 -4772
rect -1183 -4830 -1125 -4772
rect -1091 -4830 -1033 -4772
rect -999 -4830 -941 -4772
rect -907 -4830 -849 -4772
rect -815 -4830 -757 -4772
rect -723 -4830 -665 -4772
rect -631 -4830 -573 -4772
rect -539 -4830 -481 -4772
rect -447 -4830 -389 -4772
rect -355 -4830 -297 -4772
rect -263 -4830 -205 -4772
rect -171 -4830 -113 -4772
rect -79 -4830 -21 -4772
rect 13 -4830 71 -4772
rect 105 -4830 163 -4772
rect 197 -4830 255 -4772
rect 289 -4830 347 -4772
rect 381 -4830 439 -4772
rect 473 -4830 531 -4772
rect 565 -4830 623 -4772
rect 657 -4830 715 -4772
rect 749 -4830 807 -4772
rect 841 -4830 899 -4772
rect 933 -4830 991 -4772
rect 1025 -4830 1083 -4772
rect 1117 -4830 1175 -4772
rect 1209 -4830 1267 -4772
rect 1301 -4830 1359 -4772
rect 1393 -4830 1451 -4772
rect 1485 -4830 1543 -4772
rect 1577 -4830 1635 -4772
rect 1669 -4830 1727 -4772
rect 1761 -4830 1819 -4772
rect 1853 -4830 1911 -4772
rect 1945 -4830 2003 -4772
rect 2037 -4830 2095 -4772
rect 2129 -4830 2187 -4772
rect 2221 -4830 2279 -4772
rect 2313 -4830 2371 -4772
rect 2405 -4830 2463 -4772
rect 2497 -4830 2555 -4772
rect 2589 -4830 2647 -4772
rect 2681 -4830 2739 -4772
rect 2773 -4830 2831 -4772
rect 2865 -4830 2923 -4772
rect 2957 -4830 3015 -4772
rect 3049 -4830 3107 -4772
rect 3141 -4830 3199 -4772
rect 3233 -4830 3291 -4772
rect 3325 -4830 3383 -4772
rect 3417 -4830 3475 -4772
rect 3509 -4830 3567 -4772
rect 3601 -4830 3659 -4772
rect 3693 -4830 3751 -4772
rect 3785 -4830 3843 -4772
rect 3877 -4830 3935 -4772
rect 3969 -4830 4027 -4772
rect 4061 -4830 4119 -4772
rect 4153 -4830 4211 -4772
rect 4245 -4830 4303 -4772
rect 4337 -4830 4395 -4772
rect 4429 -4830 4487 -4772
rect 4521 -4830 4579 -4772
rect 4613 -4830 4671 -4772
rect 4705 -4830 4763 -4772
rect 4797 -4830 4855 -4772
rect 4889 -4830 4947 -4772
rect 4981 -4830 5039 -4772
rect 5073 -4830 5131 -4772
rect 5165 -4830 5223 -4772
rect 5257 -4830 5315 -4772
rect 5349 -4830 5407 -4772
rect 5441 -4830 5499 -4772
rect 5533 -4830 5591 -4772
rect 5625 -4830 5683 -4772
rect 5717 -4830 5775 -4772
rect 5809 -4830 5867 -4772
rect 5901 -4830 5959 -4772
rect 5993 -4830 6051 -4772
rect 6085 -4830 6143 -4772
rect 6177 -4830 6235 -4772
rect 6269 -4830 6327 -4772
rect 6361 -4830 6419 -4772
rect 6453 -4830 6511 -4772
rect 6545 -4830 6603 -4772
rect 6637 -4830 6695 -4772
rect 6729 -4830 6787 -4772
rect 6821 -4830 6879 -4772
rect 6913 -4830 6971 -4772
rect 7005 -4830 7063 -4772
rect 7097 -4830 7155 -4772
rect 7189 -4830 7247 -4772
rect 7281 -4830 7339 -4772
rect 7373 -4830 7431 -4772
rect 7465 -4830 7523 -4772
rect 7557 -4830 7615 -4772
rect 7649 -4830 7707 -4772
rect 7741 -4830 7799 -4772
rect 7833 -4830 7891 -4772
rect 7925 -4830 7983 -4772
rect 8017 -4830 8075 -4772
rect 8109 -4830 8167 -4772
rect 8201 -4830 8259 -4772
rect 8293 -4830 8351 -4772
rect 8385 -4830 8443 -4772
rect 8477 -4830 8535 -4772
rect 8569 -4830 8627 -4772
rect 8661 -4830 8719 -4772
rect 8753 -4830 8811 -4772
rect 8845 -4830 8903 -4772
rect 8937 -4830 8995 -4772
rect 9029 -4830 9087 -4772
rect 9121 -4830 9179 -4772
rect 9213 -4830 9271 -4772
rect 9305 -4830 9363 -4772
rect 9397 -4830 9455 -4772
rect 9489 -4830 9547 -4772
rect 9581 -4830 9639 -4772
rect 9673 -4830 9731 -4772
rect 9765 -4830 9823 -4772
rect 9857 -4830 9915 -4772
rect 9949 -4830 10007 -4772
rect 10041 -4830 10099 -4772
rect 10133 -4830 10191 -4772
rect 10225 -4830 10283 -4772
rect 10317 -4830 10375 -4772
rect 10409 -4830 10467 -4772
rect 10501 -4830 10559 -4772
rect 10593 -4830 10651 -4772
rect 10685 -4830 10743 -4772
rect 10777 -4830 10835 -4772
rect 10869 -4830 10927 -4772
rect 10961 -4830 11019 -4772
rect 11053 -4830 11111 -4772
rect 11145 -4830 11203 -4772
rect 11237 -4830 11295 -4772
rect 11329 -4830 11387 -4772
rect 11421 -4830 11479 -4772
rect 11513 -4830 11571 -4772
rect 11605 -4830 11663 -4772
rect 11697 -4830 11755 -4772
rect 11789 -4830 11847 -4772
rect 11881 -4830 11939 -4772
rect 11973 -4830 12031 -4772
rect 12065 -4830 12123 -4772
rect 12157 -4830 12215 -4772
rect 12249 -4830 12307 -4772
rect 12341 -4830 12399 -4772
rect 12433 -4830 12491 -4772
rect 12525 -4830 12583 -4772
rect 12617 -4830 12675 -4772
rect 12709 -4830 12767 -4772
rect 12801 -4830 12859 -4772
rect 12893 -4830 12951 -4772
rect 12985 -4830 13043 -4772
rect 13077 -4830 13135 -4772
rect 13169 -4830 13227 -4772
rect 13261 -4830 13319 -4772
rect 13353 -4830 13411 -4772
rect 13445 -4830 13503 -4772
rect 13537 -4830 13595 -4772
rect 13629 -4830 13687 -4772
rect 13721 -4830 13779 -4772
rect 13813 -4830 13871 -4772
rect 13905 -4830 13963 -4772
rect 13997 -4830 14055 -4772
rect 14089 -4830 14147 -4772
rect 14181 -4830 14239 -4772
rect 14273 -4830 14331 -4772
rect 14365 -4830 14423 -4772
rect 14457 -4830 14515 -4772
rect 14549 -4830 14607 -4772
rect 14641 -4830 14699 -4772
rect 14733 -4830 14791 -4772
rect 14825 -4830 14883 -4772
rect 14917 -4830 14975 -4772
rect 15009 -4830 15067 -4772
rect 15101 -4830 15159 -4772
rect 15193 -4830 15251 -4772
rect 15285 -4830 15343 -4772
rect 15377 -4830 15435 -4772
rect 15469 -4830 15527 -4772
rect 15561 -4830 15619 -4772
rect 15653 -4830 15711 -4772
rect 15745 -4830 15803 -4772
rect 15837 -4830 15895 -4772
rect 15929 -4830 15987 -4772
rect 16021 -4830 16079 -4772
rect 16113 -4830 16171 -4772
rect 16205 -4830 16263 -4772
rect 16297 -4830 16355 -4772
rect 16389 -4830 16447 -4772
rect 16481 -4830 16539 -4772
rect 16573 -4830 16631 -4772
rect 16665 -4830 16723 -4772
rect 16757 -4830 16815 -4772
rect 16849 -4830 16907 -4772
rect 16941 -4830 16999 -4772
rect 17033 -4830 17091 -4772
rect 17125 -4830 17183 -4772
rect 17217 -4830 17275 -4772
rect 17309 -4830 17367 -4772
rect 17401 -4830 17459 -4772
rect 17493 -4830 17551 -4772
rect 17585 -4830 17643 -4772
rect 17677 -4830 17735 -4772
rect 17769 -4830 17827 -4772
rect 17861 -4830 17919 -4772
rect 17953 -4830 18011 -4772
rect 18045 -4830 18103 -4772
rect 18137 -4830 18195 -4772
rect 18229 -4830 18287 -4772
rect 18321 -4830 18379 -4772
rect 18413 -4830 18471 -4772
rect 18505 -4830 18563 -4772
rect 18597 -4830 18655 -4772
rect 18689 -4830 18747 -4772
rect 18781 -4830 18839 -4772
rect 18873 -4830 18931 -4772
rect 18965 -4830 19023 -4772
rect 19057 -4830 19115 -4772
rect 19149 -4830 19207 -4772
rect 19241 -4830 19299 -4772
rect 19333 -4830 19391 -4772
rect 19425 -4830 19483 -4772
rect 19517 -4830 19575 -4772
rect 19609 -4830 19667 -4772
rect 19701 -4830 19759 -4772
rect 19793 -4830 19851 -4772
rect 19885 -4830 19943 -4772
rect 19977 -4830 20035 -4772
rect 20069 -4830 20127 -4772
rect 20161 -4830 20219 -4772
rect 20253 -4830 20311 -4772
rect 20345 -4830 20403 -4772
rect 20437 -4830 20495 -4772
rect 20529 -4830 20587 -4772
rect 20621 -4830 20679 -4772
rect 20713 -4830 20771 -4772
rect 20805 -4830 20863 -4772
rect 20897 -4830 20955 -4772
rect 20989 -4830 21047 -4772
rect 21081 -4830 21139 -4772
rect 21173 -4830 21231 -4772
rect 21265 -4830 21323 -4772
rect 21357 -4830 21415 -4772
rect 21449 -4830 21507 -4772
rect 21541 -4830 21599 -4772
rect 21633 -4830 21691 -4772
rect 21725 -4830 21783 -4772
rect 21817 -4830 21875 -4772
rect 21909 -4830 21967 -4772
rect 22001 -4830 22059 -4772
rect 22093 -4830 22151 -4772
rect 22185 -4830 22243 -4772
rect 22277 -4830 22335 -4772
rect 22369 -4830 22427 -4772
rect 22461 -4830 22519 -4772
rect 22553 -4830 22611 -4772
rect 22645 -4830 22703 -4772
rect 22737 -4830 22795 -4772
rect 22829 -4830 22887 -4772
rect 22921 -4830 22979 -4772
rect 23013 -4830 23071 -4772
rect 23105 -4830 23163 -4772
rect 23197 -4830 23255 -4772
rect 23289 -4830 23347 -4772
rect 23381 -4830 23439 -4772
rect 23473 -4830 23531 -4772
rect 23565 -4830 23623 -4772
rect 23657 -4830 23715 -4772
rect 23749 -4830 23807 -4772
rect 23841 -4830 23899 -4772
rect 23933 -4830 23991 -4772
rect 24025 -4830 24083 -4772
rect 24117 -4830 24175 -4772
rect 24209 -4830 24267 -4772
rect 24301 -4830 24359 -4772
rect 24393 -4830 24451 -4772
rect 24485 -4830 24543 -4772
rect 24577 -4830 24635 -4772
rect 24669 -4830 24727 -4772
rect 24761 -4830 24819 -4772
rect 24853 -4830 24911 -4772
rect 24945 -4830 25003 -4772
rect 25037 -4830 25095 -4772
rect 25129 -4830 25187 -4772
rect 25221 -4830 25279 -4772
rect 25313 -4830 25371 -4772
rect 25405 -4830 25463 -4772
rect 25497 -4830 25555 -4772
rect 25589 -4830 25647 -4772
rect 25681 -4830 25739 -4772
rect 25773 -4830 25831 -4772
rect 25865 -4830 25923 -4772
rect 25957 -4830 26015 -4772
rect 26049 -4830 26107 -4772
rect 26141 -4830 26199 -4772
rect 26233 -4830 26291 -4772
rect 26325 -4830 26383 -4772
rect 26417 -4830 26475 -4772
rect 26509 -4830 26567 -4772
rect 26601 -4830 26659 -4772
rect 26693 -4830 26751 -4772
rect 26785 -4830 26843 -4772
rect 26877 -4830 26935 -4772
rect 26969 -4830 27027 -4772
rect 27061 -4830 27119 -4772
rect 27153 -4830 27211 -4772
rect 27245 -4830 27303 -4772
rect 27337 -4830 27395 -4772
rect 27429 -4830 27487 -4772
rect 27521 -4830 27579 -4772
rect 27613 -4830 27671 -4772
rect 27705 -4830 27763 -4772
rect 27797 -4830 27855 -4772
rect 27889 -4830 27947 -4772
rect 27981 -4830 28039 -4772
rect 28073 -4830 28131 -4772
rect 28165 -4830 28223 -4772
rect 28257 -4830 28315 -4772
rect 28349 -4830 28407 -4772
rect 28441 -4830 28499 -4772
rect 28533 -4830 28591 -4772
rect 28625 -4830 28683 -4772
rect 28717 -4830 28775 -4772
rect 28809 -4830 28867 -4772
rect 28901 -4830 28959 -4772
rect 28993 -4830 29051 -4772
rect 29085 -4830 29143 -4772
rect 29177 -4830 29235 -4772
rect 29269 -4830 29327 -4772
rect 29361 -4830 29419 -4772
rect 29453 -4830 29511 -4772
rect 29545 -4830 29603 -4772
rect 29637 -4830 29695 -4772
rect 29729 -4830 29787 -4772
rect 29821 -4830 29879 -4772
rect 29913 -4830 29971 -4772
rect 30005 -4830 30063 -4772
rect 30097 -4830 30155 -4772
rect 30189 -4830 30247 -4772
rect 30281 -4830 30339 -4772
rect 30373 -4830 30431 -4772
rect 30465 -4830 30523 -4772
rect 30557 -4830 30615 -4772
rect 30649 -4830 30707 -4772
rect 30741 -4830 30799 -4772
rect 30833 -4830 30891 -4772
rect 30925 -4830 30983 -4772
rect 31017 -4830 31075 -4772
rect 31109 -4830 31167 -4772
rect 31201 -4830 31259 -4772
rect 31293 -4830 31351 -4772
rect 31385 -4830 31443 -4772
rect 31477 -4830 31535 -4772
rect 31569 -4830 31627 -4772
rect 31661 -4830 31719 -4772
rect 31753 -4830 31811 -4772
rect 31845 -4830 31903 -4772
rect 31937 -4830 31995 -4772
rect 32029 -4830 32087 -4772
rect 32121 -4830 32179 -4772
rect 32213 -4830 32271 -4772
rect 32305 -4830 32363 -4772
rect 32397 -4830 32455 -4772
rect 32489 -4830 32547 -4772
rect 32581 -4830 32639 -4772
rect 32673 -4830 32731 -4772
rect 32765 -4830 32823 -4772
rect 32857 -4830 32915 -4772
rect 32949 -4830 33007 -4772
rect 33041 -4830 33099 -4772
rect 33133 -4830 33162 -4772
rect -9158 -4846 33162 -4830
rect 4472 -7243 21243 -7011
rect 4472 -7271 21244 -7243
rect 4475 -7513 7623 -7271
rect 4475 -7551 5796 -7513
rect 6018 -7515 6068 -7513
rect 4415 -7585 4431 -7551
rect 4369 -7635 4403 -7619
rect 4369 -9027 4403 -9011
rect 4475 -9061 5796 -7585
rect 6290 -7551 7623 -7513
rect 7657 -7585 7673 -7551
rect 6010 -7635 6080 -7613
rect 6010 -7655 6027 -7635
rect 4415 -9095 4431 -9061
rect 4369 -9145 4403 -9129
rect 4369 -10537 4403 -10521
rect 4475 -10571 5796 -9095
rect 4415 -10605 4431 -10571
rect 4369 -10655 4403 -10639
rect 4369 -12047 4403 -12031
rect 4475 -12081 5796 -10605
rect 4415 -12115 4431 -12081
rect 4369 -12165 4403 -12149
rect 4369 -13557 4403 -13541
rect 4475 -13591 5796 -12115
rect 4415 -13625 4431 -13591
rect 4369 -13675 4403 -13659
rect 4369 -15067 4403 -15051
rect 4475 -15101 5796 -13625
rect 4415 -15135 4431 -15101
rect 4369 -15185 4403 -15169
rect 4369 -16577 4403 -16561
rect 4475 -16611 5796 -15135
rect 4415 -16645 4431 -16611
rect 4369 -16695 4403 -16679
rect 4369 -18087 4403 -18071
rect 4475 -18121 5796 -16645
rect 4415 -18155 4431 -18121
rect 4369 -18205 4403 -18189
rect 4369 -19597 4403 -19581
rect 4475 -19631 5796 -18155
rect 4415 -19665 4431 -19631
rect 4369 -19715 4403 -19699
rect 4369 -21107 4403 -21091
rect 4475 -21141 5796 -19665
rect 4415 -21175 4431 -21141
rect 4369 -21225 4403 -21209
rect 4369 -22617 4403 -22601
rect 4475 -22651 5796 -21175
rect 4415 -22685 4431 -22651
rect 4369 -22735 4403 -22719
rect 4369 -24127 4403 -24111
rect 4475 -24161 5796 -22685
rect 4415 -24195 4431 -24161
rect 4369 -24245 4403 -24229
rect 4369 -25637 4403 -25621
rect 4475 -25671 5796 -24195
rect 4415 -25705 4431 -25671
rect 4475 -25721 5796 -25705
rect 6018 -9011 6027 -7655
rect 6061 -7655 6080 -7635
rect 6061 -9011 6068 -7655
rect 6018 -9145 6068 -9011
rect 6018 -10521 6027 -9145
rect 6061 -10521 6068 -9145
rect 6018 -10655 6068 -10521
rect 6018 -12031 6027 -10655
rect 6061 -12031 6068 -10655
rect 6018 -12165 6068 -12031
rect 6018 -13541 6027 -12165
rect 6061 -13541 6068 -12165
rect 6018 -13675 6068 -13541
rect 6018 -15051 6027 -13675
rect 6061 -15051 6068 -13675
rect 6018 -15185 6068 -15051
rect 6018 -16561 6027 -15185
rect 6061 -16561 6068 -15185
rect 6018 -16695 6068 -16561
rect 6018 -18071 6027 -16695
rect 6061 -18071 6068 -16695
rect 6018 -18205 6068 -18071
rect 6018 -19581 6027 -18205
rect 6061 -19581 6068 -18205
rect 6018 -19715 6068 -19581
rect 6018 -21091 6027 -19715
rect 6061 -21091 6068 -19715
rect 6018 -21225 6068 -21091
rect 6018 -22601 6027 -21225
rect 6061 -22601 6068 -21225
rect 6018 -22735 6068 -22601
rect 6018 -24111 6027 -22735
rect 6061 -24111 6068 -22735
rect 6018 -24245 6068 -24111
rect 6018 -25621 6027 -24245
rect 6061 -25621 6068 -24245
rect 6018 -25721 6068 -25621
rect 6290 -7671 7623 -7585
rect 7685 -7635 7719 -7619
rect 6290 -9061 7619 -7671
rect 7685 -9027 7719 -9011
rect 7657 -9095 7673 -9061
rect 6290 -10571 7619 -9095
rect 7685 -9145 7719 -9129
rect 7685 -10537 7719 -10521
rect 7657 -10605 7673 -10571
rect 6290 -12081 7619 -10605
rect 7685 -10655 7719 -10639
rect 7685 -12047 7719 -12031
rect 7657 -12115 7673 -12081
rect 6290 -13591 7619 -12115
rect 7685 -12165 7719 -12149
rect 7685 -13557 7719 -13541
rect 7657 -13625 7673 -13591
rect 6290 -15101 7619 -13625
rect 7685 -13675 7719 -13659
rect 7685 -15067 7719 -15051
rect 7657 -15135 7673 -15101
rect 6290 -16611 7619 -15135
rect 7685 -15185 7719 -15169
rect 7685 -16577 7719 -16561
rect 7657 -16645 7673 -16611
rect 6290 -18121 7619 -16645
rect 7685 -16695 7719 -16679
rect 7685 -18087 7719 -18071
rect 7657 -18155 7673 -18121
rect 6290 -19631 7619 -18155
rect 7685 -18205 7719 -18189
rect 7685 -19597 7719 -19581
rect 7657 -19665 7673 -19631
rect 6290 -21141 7619 -19665
rect 7685 -19715 7719 -19699
rect 7685 -21107 7719 -21091
rect 7657 -21175 7673 -21141
rect 6290 -22651 7619 -21175
rect 7685 -21225 7719 -21209
rect 7685 -22617 7719 -22601
rect 7657 -22685 7673 -22651
rect 6290 -24161 7619 -22685
rect 7685 -22735 7719 -22719
rect 7685 -24127 7719 -24111
rect 7657 -24195 7673 -24161
rect 6290 -25671 7619 -24195
rect 7685 -24245 7719 -24229
rect 7685 -25637 7719 -25621
rect 7657 -25705 7673 -25671
rect 6290 -25721 7619 -25705
rect 8470 -8121 8792 -7271
rect 10028 -7379 14010 -7370
rect 10028 -7474 10166 -7379
rect 10794 -7383 14010 -7379
rect 10794 -7474 12946 -7383
rect 10028 -7478 12946 -7474
rect 13574 -7478 14010 -7383
rect 10028 -7540 14010 -7478
rect 14722 -7502 15816 -7501
rect 10032 -7541 12195 -7540
rect 12916 -7541 14010 -7540
rect 10032 -7542 11101 -7541
rect 9372 -7559 9425 -7558
rect 9372 -7594 9702 -7559
rect 9372 -7628 9516 -7594
rect 9550 -7628 9702 -7594
rect 9372 -7673 9702 -7628
rect 10032 -7665 10085 -7542
rect 10160 -7628 10176 -7594
rect 10210 -7628 10226 -7594
rect 10630 -7603 10646 -7594
rect 10501 -7628 10646 -7603
rect 10680 -7603 10696 -7594
rect 11095 -7595 12462 -7578
rect 10680 -7628 10831 -7603
rect 10032 -7673 10086 -7665
rect 9373 -7683 9702 -7673
rect 9373 -7719 9388 -7683
rect 9422 -7687 9702 -7683
rect 9422 -7719 9645 -7687
rect 9373 -7723 9645 -7719
rect 9679 -7723 9702 -7687
rect 9373 -7757 9702 -7723
rect 9373 -7793 9387 -7757
rect 9421 -7793 9645 -7757
rect 9679 -7793 9702 -7757
rect 9373 -7830 9702 -7793
rect 9373 -7866 9387 -7830
rect 9421 -7866 9644 -7830
rect 9678 -7866 9702 -7830
rect 9373 -7922 9702 -7866
rect 10033 -7683 10086 -7673
rect 10033 -7719 10048 -7683
rect 10082 -7719 10086 -7683
rect 10033 -7757 10086 -7719
rect 10033 -7793 10047 -7757
rect 10081 -7793 10086 -7757
rect 10033 -7830 10086 -7793
rect 10033 -7866 10047 -7830
rect 10081 -7866 10086 -7830
rect 10033 -7899 10086 -7866
rect 10300 -7687 10360 -7671
rect 10300 -7723 10305 -7687
rect 10339 -7723 10360 -7687
rect 10300 -7757 10360 -7723
rect 10300 -7793 10305 -7757
rect 10339 -7793 10360 -7757
rect 10300 -7830 10360 -7793
rect 10300 -7866 10304 -7830
rect 10338 -7866 10360 -7830
rect 10300 -7877 10360 -7866
rect 10501 -7683 10831 -7628
rect 10501 -7719 10518 -7683
rect 10552 -7687 10831 -7683
rect 10552 -7719 10775 -7687
rect 10501 -7723 10775 -7719
rect 10809 -7723 10831 -7687
rect 10501 -7757 10831 -7723
rect 10501 -7793 10517 -7757
rect 10551 -7793 10775 -7757
rect 10809 -7793 10831 -7757
rect 10501 -7830 10831 -7793
rect 10501 -7866 10517 -7830
rect 10551 -7866 10774 -7830
rect 10808 -7866 10831 -7830
rect 10501 -7877 10831 -7866
rect 11095 -7629 11249 -7595
rect 11283 -7629 11507 -7595
rect 11541 -7629 11765 -7595
rect 11799 -7629 12023 -7595
rect 12057 -7629 12281 -7595
rect 12315 -7629 12462 -7595
rect 11095 -7687 12462 -7629
rect 11095 -7723 11120 -7687
rect 11154 -7723 11378 -7687
rect 11412 -7723 11636 -7687
rect 11670 -7723 11894 -7687
rect 11928 -7723 12152 -7687
rect 12186 -7723 12410 -7687
rect 12444 -7723 12462 -7687
rect 11095 -7758 12462 -7723
rect 11095 -7794 11120 -7758
rect 11154 -7794 11378 -7758
rect 11412 -7794 11636 -7758
rect 11670 -7794 11894 -7758
rect 11928 -7794 12152 -7758
rect 12186 -7794 12410 -7758
rect 12444 -7794 12462 -7758
rect 11095 -7829 12462 -7794
rect 11095 -7865 11120 -7829
rect 11154 -7865 11378 -7829
rect 11412 -7865 11636 -7829
rect 11670 -7865 11894 -7829
rect 11928 -7865 12152 -7829
rect 12186 -7865 12410 -7829
rect 12444 -7865 12462 -7829
rect 9373 -7956 9516 -7922
rect 9550 -7956 9702 -7922
rect 10160 -7956 10176 -7922
rect 10210 -7956 10226 -7922
rect 9373 -8002 9702 -7956
rect 10300 -8121 10362 -7877
rect 10501 -7922 10832 -7877
rect 10501 -7956 10646 -7922
rect 10680 -7956 10832 -7922
rect 10501 -8001 10832 -7956
rect 11095 -7923 12462 -7865
rect 12916 -7687 12976 -7541
rect 13048 -7629 13064 -7595
rect 13098 -7629 13114 -7595
rect 13306 -7629 13322 -7595
rect 13356 -7629 13372 -7595
rect 12916 -7723 12935 -7687
rect 12969 -7723 12976 -7687
rect 12916 -7758 12976 -7723
rect 12916 -7794 12935 -7758
rect 12969 -7794 12976 -7758
rect 12916 -7829 12976 -7794
rect 12916 -7865 12935 -7829
rect 12969 -7865 12976 -7829
rect 12916 -7900 12976 -7865
rect 13184 -7687 13235 -7657
rect 13184 -7723 13193 -7687
rect 13227 -7723 13235 -7687
rect 13184 -7758 13235 -7723
rect 13184 -7794 13193 -7758
rect 13227 -7794 13235 -7758
rect 13184 -7829 13235 -7794
rect 13184 -7865 13193 -7829
rect 13227 -7865 13235 -7829
rect 11095 -7957 11249 -7923
rect 11283 -7957 11507 -7923
rect 11541 -7957 11765 -7923
rect 11799 -7957 12023 -7923
rect 12057 -7957 12281 -7923
rect 12315 -7957 12462 -7923
rect 13048 -7957 13064 -7923
rect 13098 -7957 13114 -7923
rect 11095 -7982 12462 -7957
rect 11369 -8001 11420 -7982
rect 11886 -8001 11937 -7982
rect 12402 -8001 12453 -7982
rect 10501 -8047 10831 -8001
rect 13184 -8014 13235 -7865
rect 13442 -7687 13493 -7541
rect 13564 -7629 13580 -7595
rect 13614 -7629 13630 -7595
rect 13822 -7629 13838 -7595
rect 13872 -7629 13888 -7595
rect 13442 -7723 13451 -7687
rect 13485 -7723 13493 -7687
rect 13442 -7758 13493 -7723
rect 13442 -7794 13451 -7758
rect 13485 -7794 13493 -7758
rect 13442 -7829 13493 -7794
rect 13442 -7865 13451 -7829
rect 13485 -7865 13493 -7829
rect 13442 -7896 13493 -7865
rect 13701 -7687 13752 -7655
rect 13958 -7670 14010 -7541
rect 14721 -7595 16080 -7502
rect 14080 -7629 14096 -7595
rect 14130 -7629 14146 -7595
rect 14721 -7629 14870 -7595
rect 14904 -7629 15128 -7595
rect 15162 -7629 15386 -7595
rect 15420 -7629 15644 -7595
rect 15678 -7629 15902 -7595
rect 15936 -7629 16080 -7595
rect 13701 -7723 13709 -7687
rect 13743 -7723 13752 -7687
rect 13701 -7758 13752 -7723
rect 13701 -7794 13709 -7758
rect 13743 -7794 13752 -7758
rect 13701 -7829 13752 -7794
rect 13701 -7865 13709 -7829
rect 13743 -7865 13752 -7829
rect 13306 -7957 13322 -7923
rect 13356 -7957 13372 -7923
rect 13564 -7957 13580 -7923
rect 13614 -7957 13630 -7923
rect 13701 -8013 13752 -7865
rect 13959 -7687 14010 -7670
rect 13959 -7723 13967 -7687
rect 14001 -7723 14010 -7687
rect 13959 -7758 14010 -7723
rect 13959 -7794 13967 -7758
rect 14001 -7794 14010 -7758
rect 13959 -7829 14010 -7794
rect 13959 -7865 13967 -7829
rect 14001 -7865 14010 -7829
rect 13959 -7896 14010 -7865
rect 14217 -7687 14268 -7656
rect 14217 -7723 14225 -7687
rect 14259 -7723 14268 -7687
rect 14217 -7758 14268 -7723
rect 14217 -7794 14225 -7758
rect 14259 -7794 14268 -7758
rect 14217 -7829 14268 -7794
rect 14217 -7865 14225 -7829
rect 14259 -7865 14268 -7829
rect 13822 -7957 13838 -7923
rect 13872 -7957 13888 -7923
rect 14080 -7957 14096 -7923
rect 14130 -7957 14146 -7923
rect 13701 -8014 13761 -8013
rect 14217 -8014 14268 -7865
rect 13184 -8121 14268 -8014
rect 14721 -7687 16080 -7629
rect 14721 -7723 14741 -7687
rect 14775 -7723 14999 -7687
rect 15033 -7723 15257 -7687
rect 15291 -7723 15515 -7687
rect 15549 -7723 15773 -7687
rect 15807 -7723 16031 -7687
rect 16065 -7723 16080 -7687
rect 14721 -7758 16080 -7723
rect 14721 -7794 14741 -7758
rect 14775 -7794 14999 -7758
rect 15033 -7794 15257 -7758
rect 15291 -7794 15515 -7758
rect 15549 -7794 15773 -7758
rect 15807 -7794 16031 -7758
rect 16065 -7794 16080 -7758
rect 14721 -7829 16080 -7794
rect 14721 -7865 14741 -7829
rect 14775 -7865 14999 -7829
rect 15033 -7865 15257 -7829
rect 15291 -7865 15515 -7829
rect 15549 -7865 15773 -7829
rect 15807 -7865 16031 -7829
rect 16065 -7865 16080 -7829
rect 14721 -7923 16080 -7865
rect 14721 -7957 14870 -7923
rect 14904 -7957 15128 -7923
rect 15162 -7957 15386 -7923
rect 15420 -7957 15644 -7923
rect 15678 -7957 15902 -7923
rect 15936 -7957 16080 -7923
rect 14721 -8064 16080 -7957
rect 16818 -8121 17140 -7271
rect 18096 -7505 21244 -7271
rect 8470 -8123 16480 -8121
rect 16516 -8123 17140 -8121
rect 8470 -8329 17140 -8123
rect 8470 -8331 8792 -8329
rect 8480 -8521 8642 -8331
rect 8479 -8535 8642 -8521
rect 8479 -8859 8641 -8535
rect 9312 -8561 9584 -8531
rect 9664 -8557 9728 -8329
rect 12332 -8521 12396 -8329
rect 9312 -8599 9408 -8561
rect 9474 -8599 9584 -8561
rect 8484 -9367 8634 -8859
rect 9312 -8685 9584 -8599
rect 9312 -8687 9516 -8685
rect 9312 -8723 9330 -8687
rect 9368 -8721 9516 -8687
rect 9554 -8721 9584 -8685
rect 9368 -8723 9584 -8721
rect 9312 -8759 9584 -8723
rect 9665 -8687 9727 -8557
rect 10698 -8561 10970 -8531
rect 10044 -8602 10060 -8568
rect 10214 -8602 10230 -8568
rect 10698 -8599 10794 -8561
rect 10860 -8599 10970 -8561
rect 9665 -8721 9691 -8687
rect 9725 -8721 9727 -8687
rect 9665 -8792 9727 -8721
rect 10549 -8687 10594 -8671
rect 10583 -8721 10594 -8687
rect 10044 -8840 10060 -8806
rect 10214 -8840 10230 -8806
rect 10549 -8949 10594 -8721
rect 10698 -8685 10970 -8599
rect 10698 -8687 10902 -8685
rect 10698 -8723 10716 -8687
rect 10754 -8721 10902 -8687
rect 10940 -8721 10970 -8685
rect 10754 -8723 10970 -8721
rect 10698 -8759 10970 -8723
rect 11068 -8561 11340 -8531
rect 11068 -8599 11164 -8561
rect 11230 -8599 11340 -8561
rect 11068 -8685 11340 -8599
rect 11068 -8687 11272 -8685
rect 11068 -8723 11086 -8687
rect 11124 -8721 11272 -8687
rect 11310 -8721 11340 -8685
rect 11124 -8723 11340 -8721
rect 11068 -8759 11340 -8723
rect 11490 -8561 11762 -8531
rect 11490 -8599 11586 -8561
rect 11652 -8599 11762 -8561
rect 11490 -8685 11762 -8599
rect 11490 -8687 11694 -8685
rect 11490 -8723 11508 -8687
rect 11546 -8721 11694 -8687
rect 11732 -8721 11762 -8685
rect 11546 -8723 11762 -8721
rect 11490 -8759 11762 -8723
rect 11912 -8561 12184 -8531
rect 12332 -8533 12397 -8521
rect 11912 -8599 12008 -8561
rect 12074 -8599 12184 -8561
rect 11912 -8685 12184 -8599
rect 11912 -8687 12116 -8685
rect 11912 -8723 11930 -8687
rect 11968 -8721 12116 -8687
rect 12154 -8721 12184 -8685
rect 11968 -8723 12184 -8721
rect 11912 -8759 12184 -8723
rect 12335 -8687 12397 -8533
rect 13412 -8561 13684 -8531
rect 12714 -8602 12730 -8568
rect 12884 -8602 12900 -8568
rect 13412 -8599 13508 -8561
rect 13574 -8599 13684 -8561
rect 12335 -8721 12361 -8687
rect 12395 -8721 12397 -8687
rect 12335 -8792 12397 -8721
rect 13219 -8687 13264 -8671
rect 13253 -8721 13264 -8687
rect 12714 -8840 12730 -8806
rect 12884 -8840 12900 -8806
rect 13219 -8931 13264 -8721
rect 13412 -8685 13684 -8599
rect 13412 -8687 13616 -8685
rect 13412 -8723 13430 -8687
rect 13468 -8721 13616 -8687
rect 13654 -8721 13684 -8685
rect 13468 -8723 13684 -8721
rect 13412 -8759 13684 -8723
rect 13782 -8561 14054 -8531
rect 13782 -8599 13878 -8561
rect 13944 -8599 14054 -8561
rect 13782 -8685 14054 -8599
rect 13782 -8687 13986 -8685
rect 13782 -8723 13800 -8687
rect 13838 -8721 13986 -8687
rect 14024 -8721 14054 -8685
rect 13838 -8723 14054 -8721
rect 13782 -8759 14054 -8723
rect 14204 -8561 14476 -8531
rect 14204 -8599 14300 -8561
rect 14366 -8599 14476 -8561
rect 14204 -8685 14476 -8599
rect 14204 -8687 14408 -8685
rect 14204 -8723 14222 -8687
rect 14260 -8721 14408 -8687
rect 14446 -8721 14476 -8685
rect 14260 -8723 14476 -8721
rect 14204 -8759 14476 -8723
rect 14626 -8561 14898 -8531
rect 14626 -8599 14722 -8561
rect 14788 -8599 14898 -8561
rect 14626 -8685 14898 -8599
rect 14626 -8687 14830 -8685
rect 14626 -8723 14644 -8687
rect 14682 -8721 14830 -8687
rect 14868 -8721 14898 -8685
rect 14682 -8723 14898 -8721
rect 14626 -8759 14898 -8723
rect 14998 -8549 15062 -8329
rect 16062 -8331 17140 -8329
rect 16062 -8333 16374 -8331
rect 16818 -8337 17140 -8331
rect 16982 -8529 17138 -8337
rect 14998 -8686 15060 -8549
rect 16066 -8561 16338 -8531
rect 15377 -8601 15393 -8567
rect 15547 -8601 15563 -8567
rect 16066 -8599 16162 -8561
rect 16228 -8599 16338 -8561
rect 16982 -8567 17139 -8529
rect 14998 -8720 15024 -8686
rect 15058 -8720 15060 -8686
rect 14998 -8791 15060 -8720
rect 15882 -8686 15927 -8670
rect 15916 -8720 15927 -8686
rect 15377 -8839 15393 -8805
rect 15547 -8839 15563 -8805
rect 10548 -8953 10594 -8949
rect 8479 -9476 8634 -9367
rect 10548 -9355 10593 -8953
rect 13218 -9355 13264 -8931
rect 15882 -8953 15927 -8720
rect 16066 -8685 16338 -8599
rect 16066 -8687 16270 -8685
rect 16066 -8723 16084 -8687
rect 16122 -8721 16270 -8687
rect 16308 -8721 16338 -8685
rect 16122 -8723 16338 -8721
rect 16066 -8759 16338 -8723
rect 10548 -9366 12889 -9355
rect 10548 -9445 12755 -9366
rect 12850 -9445 12889 -9366
rect 10548 -9460 12889 -9445
rect 10548 -9462 11219 -9460
rect 12626 -9461 12889 -9460
rect 13218 -9366 15547 -9355
rect 13218 -9445 15428 -9366
rect 15523 -9445 15547 -9366
rect 13218 -9460 15547 -9445
rect 13218 -9462 13894 -9460
rect 15299 -9461 15547 -9460
rect 15881 -9356 15927 -8953
rect 16983 -8958 17139 -8567
rect 16987 -9123 17137 -8958
rect 16640 -9253 16854 -9207
rect 16640 -9356 16664 -9253
rect 15881 -9431 16664 -9356
rect 16832 -9431 16854 -9253
rect 15881 -9461 16854 -9431
rect 8484 -13373 8634 -9476
rect 9226 -9598 9242 -9564
rect 9276 -9598 9292 -9564
rect 9484 -9598 9500 -9564
rect 9534 -9598 9550 -9564
rect 9742 -9598 9758 -9564
rect 9792 -9598 9808 -9564
rect 10000 -9598 10016 -9564
rect 10050 -9598 10066 -9564
rect 10258 -9598 10274 -9564
rect 10308 -9598 10324 -9564
rect 10516 -9598 10532 -9564
rect 10566 -9598 10582 -9564
rect 10774 -9598 10790 -9564
rect 10824 -9598 10840 -9564
rect 11032 -9598 11048 -9564
rect 11082 -9598 11098 -9564
rect 9107 -9648 9152 -9604
rect 9107 -9684 9113 -9648
rect 9147 -9684 9152 -9648
rect 9107 -9718 9152 -9684
rect 9107 -9754 9113 -9718
rect 9147 -9754 9152 -9718
rect 9107 -9788 9152 -9754
rect 9107 -9824 9113 -9788
rect 9147 -9824 9152 -9788
rect 9107 -10066 9152 -9824
rect 9365 -9648 9410 -9604
rect 9365 -9684 9371 -9648
rect 9405 -9684 9410 -9648
rect 9365 -9718 9410 -9684
rect 9365 -9754 9371 -9718
rect 9405 -9754 9410 -9718
rect 9365 -9788 9410 -9754
rect 9365 -9824 9371 -9788
rect 9405 -9824 9410 -9788
rect 9226 -9908 9242 -9874
rect 9276 -9908 9292 -9874
rect 9226 -10016 9242 -9982
rect 9276 -10016 9292 -9982
rect 9107 -10102 9113 -10066
rect 9147 -10102 9152 -10066
rect 9107 -10136 9152 -10102
rect 9107 -10172 9113 -10136
rect 9147 -10172 9152 -10136
rect 9107 -10206 9152 -10172
rect 9107 -10242 9113 -10206
rect 9147 -10242 9152 -10206
rect 9107 -10484 9152 -10242
rect 9365 -10066 9410 -9824
rect 9622 -9648 9667 -9604
rect 9622 -9684 9629 -9648
rect 9663 -9684 9667 -9648
rect 9622 -9718 9667 -9684
rect 9622 -9754 9629 -9718
rect 9663 -9754 9667 -9718
rect 9622 -9789 9667 -9754
rect 9622 -9825 9629 -9789
rect 9663 -9825 9667 -9789
rect 9484 -9908 9500 -9874
rect 9534 -9908 9550 -9874
rect 9484 -10016 9500 -9982
rect 9534 -10016 9550 -9982
rect 9365 -10102 9371 -10066
rect 9405 -10102 9410 -10066
rect 9365 -10136 9410 -10102
rect 9365 -10172 9371 -10136
rect 9405 -10172 9410 -10136
rect 9365 -10206 9410 -10172
rect 9365 -10242 9371 -10206
rect 9405 -10242 9410 -10206
rect 9226 -10326 9242 -10292
rect 9276 -10326 9292 -10292
rect 9226 -10434 9242 -10400
rect 9276 -10434 9292 -10400
rect 9107 -10520 9113 -10484
rect 9147 -10520 9152 -10484
rect 9107 -10554 9152 -10520
rect 9107 -10590 9113 -10554
rect 9147 -10590 9152 -10554
rect 9107 -10624 9152 -10590
rect 9107 -10660 9113 -10624
rect 9147 -10660 9152 -10624
rect 9107 -10902 9152 -10660
rect 9365 -10484 9410 -10242
rect 9622 -10066 9667 -9825
rect 9882 -9648 9927 -9604
rect 9882 -9684 9887 -9648
rect 9921 -9684 9927 -9648
rect 9882 -9718 9927 -9684
rect 9882 -9754 9887 -9718
rect 9921 -9754 9927 -9718
rect 9882 -9788 9927 -9754
rect 9882 -9824 9887 -9788
rect 9921 -9824 9927 -9788
rect 9742 -9908 9758 -9874
rect 9792 -9908 9808 -9874
rect 9742 -10016 9758 -9982
rect 9792 -10016 9808 -9982
rect 9622 -10102 9629 -10066
rect 9663 -10102 9667 -10066
rect 9622 -10136 9667 -10102
rect 9622 -10172 9629 -10136
rect 9663 -10172 9667 -10136
rect 9622 -10207 9667 -10172
rect 9622 -10243 9629 -10207
rect 9663 -10243 9667 -10207
rect 9484 -10326 9500 -10292
rect 9534 -10326 9550 -10292
rect 9484 -10434 9500 -10400
rect 9534 -10434 9550 -10400
rect 9365 -10520 9371 -10484
rect 9405 -10520 9410 -10484
rect 9365 -10554 9410 -10520
rect 9365 -10590 9371 -10554
rect 9405 -10590 9410 -10554
rect 9365 -10624 9410 -10590
rect 9365 -10660 9371 -10624
rect 9405 -10660 9410 -10624
rect 9226 -10744 9242 -10710
rect 9276 -10744 9292 -10710
rect 9226 -10852 9242 -10818
rect 9276 -10852 9292 -10818
rect 9107 -10938 9113 -10902
rect 9147 -10938 9152 -10902
rect 9107 -10972 9152 -10938
rect 9107 -11008 9113 -10972
rect 9147 -11008 9152 -10972
rect 9107 -11042 9152 -11008
rect 9107 -11078 9113 -11042
rect 9147 -11078 9152 -11042
rect 9107 -11320 9152 -11078
rect 9365 -10902 9410 -10660
rect 9622 -10484 9667 -10243
rect 9882 -10066 9927 -9824
rect 10140 -9648 10185 -9604
rect 10140 -9684 10145 -9648
rect 10179 -9684 10185 -9648
rect 10140 -9718 10185 -9684
rect 10140 -9754 10145 -9718
rect 10179 -9754 10185 -9718
rect 10140 -9788 10185 -9754
rect 10140 -9824 10145 -9788
rect 10179 -9824 10185 -9788
rect 10000 -9908 10016 -9874
rect 10050 -9908 10066 -9874
rect 10000 -10016 10016 -9982
rect 10050 -10016 10066 -9982
rect 9882 -10102 9887 -10066
rect 9921 -10102 9927 -10066
rect 9882 -10136 9927 -10102
rect 9882 -10172 9887 -10136
rect 9921 -10172 9927 -10136
rect 9882 -10206 9927 -10172
rect 9882 -10242 9887 -10206
rect 9921 -10242 9927 -10206
rect 9742 -10326 9758 -10292
rect 9792 -10326 9808 -10292
rect 9742 -10434 9758 -10400
rect 9792 -10434 9808 -10400
rect 9622 -10520 9629 -10484
rect 9663 -10520 9667 -10484
rect 9622 -10554 9667 -10520
rect 9622 -10590 9629 -10554
rect 9663 -10590 9667 -10554
rect 9622 -10625 9667 -10590
rect 9622 -10661 9629 -10625
rect 9663 -10661 9667 -10625
rect 9484 -10744 9500 -10710
rect 9534 -10744 9550 -10710
rect 9484 -10852 9500 -10818
rect 9534 -10852 9550 -10818
rect 9365 -10938 9371 -10902
rect 9405 -10938 9410 -10902
rect 9365 -10972 9410 -10938
rect 9365 -11008 9371 -10972
rect 9405 -11008 9410 -10972
rect 9365 -11042 9410 -11008
rect 9365 -11078 9371 -11042
rect 9405 -11078 9410 -11042
rect 9226 -11162 9242 -11128
rect 9276 -11162 9292 -11128
rect 9226 -11270 9242 -11236
rect 9276 -11270 9292 -11236
rect 9107 -11356 9113 -11320
rect 9147 -11356 9152 -11320
rect 9107 -11390 9152 -11356
rect 9107 -11426 9113 -11390
rect 9147 -11426 9152 -11390
rect 9107 -11460 9152 -11426
rect 9107 -11496 9113 -11460
rect 9147 -11496 9152 -11460
rect 9107 -11738 9152 -11496
rect 9365 -11320 9410 -11078
rect 9622 -10902 9667 -10661
rect 9882 -10484 9927 -10242
rect 10140 -10066 10185 -9824
rect 10397 -9648 10442 -9604
rect 10397 -9684 10403 -9648
rect 10437 -9684 10442 -9648
rect 10397 -9718 10442 -9684
rect 10397 -9754 10403 -9718
rect 10437 -9754 10442 -9718
rect 10397 -9788 10442 -9754
rect 10397 -9824 10403 -9788
rect 10437 -9824 10442 -9788
rect 10258 -9908 10274 -9874
rect 10308 -9908 10324 -9874
rect 10258 -10016 10274 -9982
rect 10308 -10016 10324 -9982
rect 10140 -10102 10145 -10066
rect 10179 -10102 10185 -10066
rect 10140 -10136 10185 -10102
rect 10140 -10172 10145 -10136
rect 10179 -10172 10185 -10136
rect 10140 -10206 10185 -10172
rect 10140 -10242 10145 -10206
rect 10179 -10242 10185 -10206
rect 10000 -10326 10016 -10292
rect 10050 -10326 10066 -10292
rect 10000 -10434 10016 -10400
rect 10050 -10434 10066 -10400
rect 9882 -10520 9887 -10484
rect 9921 -10520 9927 -10484
rect 9882 -10554 9927 -10520
rect 9882 -10590 9887 -10554
rect 9921 -10590 9927 -10554
rect 9882 -10624 9927 -10590
rect 9882 -10660 9887 -10624
rect 9921 -10660 9927 -10624
rect 9742 -10744 9758 -10710
rect 9792 -10744 9808 -10710
rect 9742 -10852 9758 -10818
rect 9792 -10852 9808 -10818
rect 9622 -10938 9629 -10902
rect 9663 -10938 9667 -10902
rect 9622 -10972 9667 -10938
rect 9622 -11008 9629 -10972
rect 9663 -11008 9667 -10972
rect 9622 -11043 9667 -11008
rect 9622 -11079 9629 -11043
rect 9663 -11079 9667 -11043
rect 9484 -11162 9500 -11128
rect 9534 -11162 9550 -11128
rect 9484 -11270 9500 -11236
rect 9534 -11270 9550 -11236
rect 9365 -11356 9371 -11320
rect 9405 -11356 9410 -11320
rect 9365 -11390 9410 -11356
rect 9365 -11426 9371 -11390
rect 9405 -11426 9410 -11390
rect 9365 -11460 9410 -11426
rect 9365 -11496 9371 -11460
rect 9405 -11496 9410 -11460
rect 9226 -11580 9242 -11546
rect 9276 -11580 9292 -11546
rect 9226 -11688 9242 -11654
rect 9276 -11688 9292 -11654
rect 9107 -11774 9113 -11738
rect 9147 -11774 9152 -11738
rect 9107 -11808 9152 -11774
rect 9107 -11844 9113 -11808
rect 9147 -11844 9152 -11808
rect 9107 -11878 9152 -11844
rect 9107 -11914 9113 -11878
rect 9147 -11914 9152 -11878
rect 9107 -12156 9152 -11914
rect 9365 -11738 9410 -11496
rect 9622 -11320 9667 -11079
rect 9882 -10902 9927 -10660
rect 10140 -10484 10185 -10242
rect 10397 -10066 10442 -9824
rect 10654 -9648 10699 -9604
rect 10654 -9684 10661 -9648
rect 10695 -9684 10699 -9648
rect 10654 -9718 10699 -9684
rect 10654 -9754 10661 -9718
rect 10695 -9754 10699 -9718
rect 10654 -9788 10699 -9754
rect 10654 -9824 10661 -9788
rect 10695 -9824 10699 -9788
rect 10516 -9908 10532 -9874
rect 10566 -9908 10582 -9874
rect 10516 -10016 10532 -9982
rect 10566 -10016 10582 -9982
rect 10397 -10102 10403 -10066
rect 10437 -10102 10442 -10066
rect 10397 -10136 10442 -10102
rect 10397 -10172 10403 -10136
rect 10437 -10172 10442 -10136
rect 10397 -10206 10442 -10172
rect 10397 -10242 10403 -10206
rect 10437 -10242 10442 -10206
rect 10258 -10326 10274 -10292
rect 10308 -10326 10324 -10292
rect 10258 -10434 10274 -10400
rect 10308 -10434 10324 -10400
rect 10140 -10520 10145 -10484
rect 10179 -10520 10185 -10484
rect 10140 -10554 10185 -10520
rect 10140 -10590 10145 -10554
rect 10179 -10590 10185 -10554
rect 10140 -10624 10185 -10590
rect 10140 -10660 10145 -10624
rect 10179 -10660 10185 -10624
rect 10000 -10744 10016 -10710
rect 10050 -10744 10066 -10710
rect 10000 -10852 10016 -10818
rect 10050 -10852 10066 -10818
rect 9882 -10938 9887 -10902
rect 9921 -10938 9927 -10902
rect 9882 -10972 9927 -10938
rect 9882 -11008 9887 -10972
rect 9921 -11008 9927 -10972
rect 9882 -11042 9927 -11008
rect 9882 -11078 9887 -11042
rect 9921 -11078 9927 -11042
rect 9742 -11162 9758 -11128
rect 9792 -11162 9808 -11128
rect 9742 -11270 9758 -11236
rect 9792 -11270 9808 -11236
rect 9622 -11356 9629 -11320
rect 9663 -11356 9667 -11320
rect 9622 -11390 9667 -11356
rect 9622 -11426 9629 -11390
rect 9663 -11426 9667 -11390
rect 9622 -11461 9667 -11426
rect 9622 -11497 9629 -11461
rect 9663 -11497 9667 -11461
rect 9484 -11580 9500 -11546
rect 9534 -11580 9550 -11546
rect 9484 -11688 9500 -11654
rect 9534 -11688 9550 -11654
rect 9365 -11774 9371 -11738
rect 9405 -11774 9410 -11738
rect 9365 -11808 9410 -11774
rect 9365 -11844 9371 -11808
rect 9405 -11844 9410 -11808
rect 9365 -11878 9410 -11844
rect 9365 -11914 9371 -11878
rect 9405 -11914 9410 -11878
rect 9226 -11998 9242 -11964
rect 9276 -11998 9292 -11964
rect 9226 -12106 9242 -12072
rect 9276 -12106 9292 -12072
rect 9107 -12192 9113 -12156
rect 9147 -12192 9152 -12156
rect 9107 -12226 9152 -12192
rect 9107 -12262 9113 -12226
rect 9147 -12262 9152 -12226
rect 9107 -12296 9152 -12262
rect 9107 -12332 9113 -12296
rect 9147 -12332 9152 -12296
rect 9107 -12574 9152 -12332
rect 9365 -12156 9410 -11914
rect 9622 -11738 9667 -11497
rect 9882 -11320 9927 -11078
rect 10140 -10902 10185 -10660
rect 10397 -10484 10442 -10242
rect 10654 -10066 10699 -9824
rect 10913 -9648 10958 -9604
rect 10913 -9684 10919 -9648
rect 10953 -9684 10958 -9648
rect 10913 -9718 10958 -9684
rect 10913 -9754 10919 -9718
rect 10953 -9754 10958 -9718
rect 10913 -9788 10958 -9754
rect 10913 -9824 10919 -9788
rect 10953 -9824 10958 -9788
rect 10774 -9908 10790 -9874
rect 10824 -9908 10840 -9874
rect 10774 -10016 10790 -9982
rect 10824 -10016 10840 -9982
rect 10654 -10102 10661 -10066
rect 10695 -10102 10699 -10066
rect 10654 -10136 10699 -10102
rect 10654 -10172 10661 -10136
rect 10695 -10172 10699 -10136
rect 10654 -10206 10699 -10172
rect 10654 -10242 10661 -10206
rect 10695 -10242 10699 -10206
rect 10516 -10326 10532 -10292
rect 10566 -10326 10582 -10292
rect 10516 -10434 10532 -10400
rect 10566 -10434 10582 -10400
rect 10397 -10520 10403 -10484
rect 10437 -10520 10442 -10484
rect 10397 -10554 10442 -10520
rect 10397 -10590 10403 -10554
rect 10437 -10590 10442 -10554
rect 10397 -10624 10442 -10590
rect 10397 -10660 10403 -10624
rect 10437 -10660 10442 -10624
rect 10258 -10744 10274 -10710
rect 10308 -10744 10324 -10710
rect 10258 -10852 10274 -10818
rect 10308 -10852 10324 -10818
rect 10140 -10938 10145 -10902
rect 10179 -10938 10185 -10902
rect 10140 -10972 10185 -10938
rect 10140 -11008 10145 -10972
rect 10179 -11008 10185 -10972
rect 10140 -11042 10185 -11008
rect 10140 -11078 10145 -11042
rect 10179 -11078 10185 -11042
rect 10000 -11162 10016 -11128
rect 10050 -11162 10066 -11128
rect 10000 -11270 10016 -11236
rect 10050 -11270 10066 -11236
rect 9882 -11356 9887 -11320
rect 9921 -11356 9927 -11320
rect 9882 -11390 9927 -11356
rect 9882 -11426 9887 -11390
rect 9921 -11426 9927 -11390
rect 9882 -11460 9927 -11426
rect 9882 -11496 9887 -11460
rect 9921 -11496 9927 -11460
rect 9742 -11580 9758 -11546
rect 9792 -11580 9808 -11546
rect 9742 -11688 9758 -11654
rect 9792 -11688 9808 -11654
rect 9622 -11774 9629 -11738
rect 9663 -11774 9667 -11738
rect 9622 -11808 9667 -11774
rect 9622 -11844 9629 -11808
rect 9663 -11844 9667 -11808
rect 9622 -11879 9667 -11844
rect 9622 -11915 9629 -11879
rect 9663 -11915 9667 -11879
rect 9484 -11998 9500 -11964
rect 9534 -11998 9550 -11964
rect 9484 -12106 9500 -12072
rect 9534 -12106 9550 -12072
rect 9365 -12192 9371 -12156
rect 9405 -12192 9410 -12156
rect 9365 -12226 9410 -12192
rect 9365 -12262 9371 -12226
rect 9405 -12262 9410 -12226
rect 9365 -12296 9410 -12262
rect 9365 -12332 9371 -12296
rect 9405 -12332 9410 -12296
rect 9226 -12416 9242 -12382
rect 9276 -12416 9292 -12382
rect 9365 -12450 9410 -12332
rect 9622 -12156 9667 -11915
rect 9882 -11738 9927 -11496
rect 10140 -11320 10185 -11078
rect 10397 -10902 10442 -10660
rect 10654 -10484 10699 -10242
rect 10913 -10066 10958 -9824
rect 11171 -9648 11216 -9462
rect 11896 -9598 11912 -9564
rect 11946 -9598 11962 -9564
rect 12154 -9598 12170 -9564
rect 12204 -9598 12220 -9564
rect 12412 -9598 12428 -9564
rect 12462 -9598 12478 -9564
rect 12670 -9598 12686 -9564
rect 12720 -9598 12736 -9564
rect 12928 -9598 12944 -9564
rect 12978 -9598 12994 -9564
rect 13186 -9598 13202 -9564
rect 13236 -9598 13252 -9564
rect 13444 -9598 13460 -9564
rect 13494 -9598 13510 -9564
rect 13702 -9598 13718 -9564
rect 13752 -9598 13768 -9564
rect 11171 -9684 11177 -9648
rect 11211 -9684 11216 -9648
rect 11171 -9718 11216 -9684
rect 11171 -9754 11177 -9718
rect 11211 -9754 11216 -9718
rect 11171 -9788 11216 -9754
rect 11171 -9824 11177 -9788
rect 11211 -9824 11216 -9788
rect 11032 -9908 11048 -9874
rect 11082 -9908 11098 -9874
rect 11032 -10016 11048 -9982
rect 11082 -10016 11098 -9982
rect 10913 -10102 10919 -10066
rect 10953 -10102 10958 -10066
rect 10913 -10136 10958 -10102
rect 10913 -10172 10919 -10136
rect 10953 -10172 10958 -10136
rect 10913 -10206 10958 -10172
rect 10913 -10242 10919 -10206
rect 10953 -10242 10958 -10206
rect 10774 -10326 10790 -10292
rect 10824 -10326 10840 -10292
rect 10774 -10434 10790 -10400
rect 10824 -10434 10840 -10400
rect 10654 -10520 10661 -10484
rect 10695 -10520 10699 -10484
rect 10654 -10554 10699 -10520
rect 10654 -10590 10661 -10554
rect 10695 -10590 10699 -10554
rect 10654 -10624 10699 -10590
rect 10654 -10660 10661 -10624
rect 10695 -10660 10699 -10624
rect 10516 -10744 10532 -10710
rect 10566 -10744 10582 -10710
rect 10516 -10852 10532 -10818
rect 10566 -10852 10582 -10818
rect 10397 -10938 10403 -10902
rect 10437 -10938 10442 -10902
rect 10397 -10972 10442 -10938
rect 10397 -11008 10403 -10972
rect 10437 -11008 10442 -10972
rect 10397 -11042 10442 -11008
rect 10397 -11078 10403 -11042
rect 10437 -11078 10442 -11042
rect 10258 -11162 10274 -11128
rect 10308 -11162 10324 -11128
rect 10258 -11270 10274 -11236
rect 10308 -11270 10324 -11236
rect 10140 -11356 10145 -11320
rect 10179 -11356 10185 -11320
rect 10140 -11390 10185 -11356
rect 10140 -11426 10145 -11390
rect 10179 -11426 10185 -11390
rect 10140 -11460 10185 -11426
rect 10140 -11496 10145 -11460
rect 10179 -11496 10185 -11460
rect 10000 -11580 10016 -11546
rect 10050 -11580 10066 -11546
rect 10000 -11688 10016 -11654
rect 10050 -11688 10066 -11654
rect 9882 -11774 9887 -11738
rect 9921 -11774 9927 -11738
rect 9882 -11808 9927 -11774
rect 9882 -11844 9887 -11808
rect 9921 -11844 9927 -11808
rect 9882 -11878 9927 -11844
rect 9882 -11914 9887 -11878
rect 9921 -11914 9927 -11878
rect 9742 -11998 9758 -11964
rect 9792 -11998 9808 -11964
rect 9742 -12106 9758 -12072
rect 9792 -12106 9808 -12072
rect 9622 -12192 9629 -12156
rect 9663 -12192 9667 -12156
rect 9622 -12226 9667 -12192
rect 9622 -12262 9629 -12226
rect 9663 -12262 9667 -12226
rect 9622 -12297 9667 -12262
rect 9622 -12333 9629 -12297
rect 9663 -12333 9667 -12297
rect 9484 -12416 9500 -12382
rect 9534 -12416 9550 -12382
rect 9622 -12450 9667 -12333
rect 9882 -12156 9927 -11914
rect 10140 -11738 10185 -11496
rect 10397 -11320 10442 -11078
rect 10654 -10902 10699 -10660
rect 10913 -10484 10958 -10242
rect 11171 -10066 11216 -9824
rect 11171 -10102 11177 -10066
rect 11211 -10102 11216 -10066
rect 11171 -10136 11216 -10102
rect 11171 -10172 11177 -10136
rect 11211 -10172 11216 -10136
rect 11171 -10206 11216 -10172
rect 11171 -10242 11177 -10206
rect 11211 -10242 11216 -10206
rect 11032 -10326 11048 -10292
rect 11082 -10326 11098 -10292
rect 11032 -10434 11048 -10400
rect 11082 -10434 11098 -10400
rect 10913 -10520 10919 -10484
rect 10953 -10520 10958 -10484
rect 10913 -10554 10958 -10520
rect 10913 -10590 10919 -10554
rect 10953 -10590 10958 -10554
rect 10913 -10624 10958 -10590
rect 10913 -10660 10919 -10624
rect 10953 -10660 10958 -10624
rect 10774 -10744 10790 -10710
rect 10824 -10744 10840 -10710
rect 10774 -10852 10790 -10818
rect 10824 -10852 10840 -10818
rect 10654 -10938 10661 -10902
rect 10695 -10938 10699 -10902
rect 10654 -10972 10699 -10938
rect 10654 -11008 10661 -10972
rect 10695 -11008 10699 -10972
rect 10654 -11042 10699 -11008
rect 10654 -11078 10661 -11042
rect 10695 -11078 10699 -11042
rect 10516 -11162 10532 -11128
rect 10566 -11162 10582 -11128
rect 10516 -11270 10532 -11236
rect 10566 -11270 10582 -11236
rect 10397 -11356 10403 -11320
rect 10437 -11356 10442 -11320
rect 10397 -11390 10442 -11356
rect 10397 -11426 10403 -11390
rect 10437 -11426 10442 -11390
rect 10397 -11460 10442 -11426
rect 10397 -11496 10403 -11460
rect 10437 -11496 10442 -11460
rect 10258 -11580 10274 -11546
rect 10308 -11580 10324 -11546
rect 10258 -11688 10274 -11654
rect 10308 -11688 10324 -11654
rect 10140 -11774 10145 -11738
rect 10179 -11774 10185 -11738
rect 10140 -11808 10185 -11774
rect 10140 -11844 10145 -11808
rect 10179 -11844 10185 -11808
rect 10140 -11878 10185 -11844
rect 10140 -11914 10145 -11878
rect 10179 -11914 10185 -11878
rect 10000 -11998 10016 -11964
rect 10050 -11998 10066 -11964
rect 10000 -12106 10016 -12072
rect 10050 -12106 10066 -12072
rect 9882 -12192 9887 -12156
rect 9921 -12192 9927 -12156
rect 9882 -12226 9927 -12192
rect 9882 -12262 9887 -12226
rect 9921 -12262 9927 -12226
rect 9882 -12296 9927 -12262
rect 9882 -12332 9887 -12296
rect 9921 -12332 9927 -12296
rect 9742 -12416 9758 -12382
rect 9792 -12416 9808 -12382
rect 9882 -12450 9927 -12332
rect 10140 -12156 10185 -11914
rect 10397 -11738 10442 -11496
rect 10654 -11320 10699 -11078
rect 10913 -10902 10958 -10660
rect 11171 -10484 11216 -10242
rect 11171 -10520 11177 -10484
rect 11211 -10520 11216 -10484
rect 11171 -10554 11216 -10520
rect 11171 -10590 11177 -10554
rect 11211 -10590 11216 -10554
rect 11171 -10624 11216 -10590
rect 11171 -10660 11177 -10624
rect 11211 -10660 11216 -10624
rect 11032 -10744 11048 -10710
rect 11082 -10744 11098 -10710
rect 11032 -10852 11048 -10818
rect 11082 -10852 11098 -10818
rect 10913 -10938 10919 -10902
rect 10953 -10938 10958 -10902
rect 10913 -10972 10958 -10938
rect 10913 -11008 10919 -10972
rect 10953 -11008 10958 -10972
rect 10913 -11042 10958 -11008
rect 10913 -11078 10919 -11042
rect 10953 -11078 10958 -11042
rect 10774 -11162 10790 -11128
rect 10824 -11162 10840 -11128
rect 10774 -11270 10790 -11236
rect 10824 -11270 10840 -11236
rect 10654 -11356 10661 -11320
rect 10695 -11356 10699 -11320
rect 10654 -11390 10699 -11356
rect 10654 -11426 10661 -11390
rect 10695 -11426 10699 -11390
rect 10654 -11460 10699 -11426
rect 10654 -11496 10661 -11460
rect 10695 -11496 10699 -11460
rect 10516 -11580 10532 -11546
rect 10566 -11580 10582 -11546
rect 10516 -11688 10532 -11654
rect 10566 -11688 10582 -11654
rect 10397 -11774 10403 -11738
rect 10437 -11774 10442 -11738
rect 10397 -11808 10442 -11774
rect 10397 -11844 10403 -11808
rect 10437 -11844 10442 -11808
rect 10397 -11878 10442 -11844
rect 10397 -11914 10403 -11878
rect 10437 -11914 10442 -11878
rect 10258 -11998 10274 -11964
rect 10308 -11998 10324 -11964
rect 10258 -12106 10274 -12072
rect 10308 -12106 10324 -12072
rect 10140 -12192 10145 -12156
rect 10179 -12192 10185 -12156
rect 10140 -12226 10185 -12192
rect 10140 -12262 10145 -12226
rect 10179 -12262 10185 -12226
rect 10140 -12296 10185 -12262
rect 10140 -12332 10145 -12296
rect 10179 -12332 10185 -12296
rect 10000 -12416 10016 -12382
rect 10050 -12416 10066 -12382
rect 10140 -12450 10185 -12332
rect 10397 -12156 10442 -11914
rect 10654 -11738 10699 -11496
rect 10913 -11320 10958 -11078
rect 11171 -10902 11216 -10660
rect 11171 -10938 11177 -10902
rect 11211 -10938 11216 -10902
rect 11171 -10972 11216 -10938
rect 11171 -11008 11177 -10972
rect 11211 -11008 11216 -10972
rect 11171 -11042 11216 -11008
rect 11171 -11078 11177 -11042
rect 11211 -11078 11216 -11042
rect 11032 -11162 11048 -11128
rect 11082 -11162 11098 -11128
rect 11032 -11270 11048 -11236
rect 11082 -11270 11098 -11236
rect 10913 -11356 10919 -11320
rect 10953 -11356 10958 -11320
rect 10913 -11390 10958 -11356
rect 10913 -11426 10919 -11390
rect 10953 -11426 10958 -11390
rect 10913 -11460 10958 -11426
rect 10913 -11496 10919 -11460
rect 10953 -11496 10958 -11460
rect 10774 -11580 10790 -11546
rect 10824 -11580 10840 -11546
rect 10774 -11688 10790 -11654
rect 10824 -11688 10840 -11654
rect 10654 -11774 10661 -11738
rect 10695 -11774 10699 -11738
rect 10654 -11808 10699 -11774
rect 10654 -11844 10661 -11808
rect 10695 -11844 10699 -11808
rect 10654 -11878 10699 -11844
rect 10654 -11914 10661 -11878
rect 10695 -11914 10699 -11878
rect 10516 -11998 10532 -11964
rect 10566 -11998 10582 -11964
rect 10516 -12106 10532 -12072
rect 10566 -12106 10582 -12072
rect 10397 -12192 10403 -12156
rect 10437 -12192 10442 -12156
rect 10397 -12226 10442 -12192
rect 10397 -12262 10403 -12226
rect 10437 -12262 10442 -12226
rect 10397 -12296 10442 -12262
rect 10397 -12332 10403 -12296
rect 10437 -12332 10442 -12296
rect 10258 -12416 10274 -12382
rect 10308 -12416 10324 -12382
rect 10397 -12450 10442 -12332
rect 10654 -12156 10699 -11914
rect 10913 -11738 10958 -11496
rect 11171 -11320 11216 -11078
rect 11171 -11356 11177 -11320
rect 11211 -11356 11216 -11320
rect 11171 -11390 11216 -11356
rect 11171 -11426 11177 -11390
rect 11211 -11426 11216 -11390
rect 11171 -11460 11216 -11426
rect 11171 -11496 11177 -11460
rect 11211 -11496 11216 -11460
rect 11032 -11580 11048 -11546
rect 11082 -11580 11098 -11546
rect 11032 -11688 11048 -11654
rect 11082 -11688 11098 -11654
rect 10913 -11774 10919 -11738
rect 10953 -11774 10958 -11738
rect 10913 -11808 10958 -11774
rect 10913 -11844 10919 -11808
rect 10953 -11844 10958 -11808
rect 10913 -11878 10958 -11844
rect 10913 -11914 10919 -11878
rect 10953 -11914 10958 -11878
rect 10774 -11998 10790 -11964
rect 10824 -11998 10840 -11964
rect 10774 -12106 10790 -12072
rect 10824 -12106 10840 -12072
rect 10654 -12192 10661 -12156
rect 10695 -12192 10699 -12156
rect 10654 -12226 10699 -12192
rect 10654 -12262 10661 -12226
rect 10695 -12262 10699 -12226
rect 10654 -12296 10699 -12262
rect 10654 -12332 10661 -12296
rect 10695 -12332 10699 -12296
rect 10516 -12416 10532 -12382
rect 10566 -12416 10582 -12382
rect 10654 -12450 10699 -12332
rect 10913 -12156 10958 -11914
rect 11171 -11738 11216 -11496
rect 11171 -11774 11177 -11738
rect 11211 -11774 11216 -11738
rect 11171 -11808 11216 -11774
rect 11171 -11844 11177 -11808
rect 11211 -11844 11216 -11808
rect 11171 -11878 11216 -11844
rect 11171 -11914 11177 -11878
rect 11211 -11914 11216 -11878
rect 11032 -11998 11048 -11964
rect 11082 -11998 11098 -11964
rect 11032 -12106 11048 -12072
rect 11082 -12106 11098 -12072
rect 10913 -12192 10919 -12156
rect 10953 -12192 10958 -12156
rect 10913 -12226 10958 -12192
rect 10913 -12262 10919 -12226
rect 10953 -12262 10958 -12226
rect 10913 -12296 10958 -12262
rect 10913 -12332 10919 -12296
rect 10953 -12332 10958 -12296
rect 10774 -12416 10790 -12382
rect 10824 -12416 10840 -12382
rect 10913 -12450 10958 -12332
rect 11171 -12156 11216 -11914
rect 11171 -12192 11177 -12156
rect 11211 -12192 11216 -12156
rect 11171 -12226 11216 -12192
rect 11171 -12262 11177 -12226
rect 11211 -12262 11216 -12226
rect 11171 -12296 11216 -12262
rect 11171 -12332 11177 -12296
rect 11211 -12332 11216 -12296
rect 11032 -12416 11048 -12382
rect 11082 -12416 11098 -12382
rect 11171 -12450 11216 -12332
rect 11777 -9648 11822 -9604
rect 11777 -9684 11783 -9648
rect 11817 -9684 11822 -9648
rect 11777 -9718 11822 -9684
rect 11777 -9754 11783 -9718
rect 11817 -9754 11822 -9718
rect 11777 -9788 11822 -9754
rect 11777 -9824 11783 -9788
rect 11817 -9824 11822 -9788
rect 11777 -10066 11822 -9824
rect 12035 -9648 12080 -9604
rect 12035 -9684 12041 -9648
rect 12075 -9684 12080 -9648
rect 12035 -9718 12080 -9684
rect 12035 -9754 12041 -9718
rect 12075 -9754 12080 -9718
rect 12035 -9788 12080 -9754
rect 12035 -9824 12041 -9788
rect 12075 -9824 12080 -9788
rect 11896 -9908 11912 -9874
rect 11946 -9908 11962 -9874
rect 11896 -10016 11912 -9982
rect 11946 -10016 11962 -9982
rect 11777 -10102 11783 -10066
rect 11817 -10102 11822 -10066
rect 11777 -10136 11822 -10102
rect 11777 -10172 11783 -10136
rect 11817 -10172 11822 -10136
rect 11777 -10206 11822 -10172
rect 11777 -10242 11783 -10206
rect 11817 -10242 11822 -10206
rect 11777 -10484 11822 -10242
rect 12035 -10066 12080 -9824
rect 12292 -9648 12337 -9604
rect 12292 -9684 12299 -9648
rect 12333 -9684 12337 -9648
rect 12292 -9718 12337 -9684
rect 12292 -9754 12299 -9718
rect 12333 -9754 12337 -9718
rect 12292 -9789 12337 -9754
rect 12292 -9825 12299 -9789
rect 12333 -9825 12337 -9789
rect 12154 -9908 12170 -9874
rect 12204 -9908 12220 -9874
rect 12154 -10016 12170 -9982
rect 12204 -10016 12220 -9982
rect 12035 -10102 12041 -10066
rect 12075 -10102 12080 -10066
rect 12035 -10136 12080 -10102
rect 12035 -10172 12041 -10136
rect 12075 -10172 12080 -10136
rect 12035 -10206 12080 -10172
rect 12035 -10242 12041 -10206
rect 12075 -10242 12080 -10206
rect 11896 -10326 11912 -10292
rect 11946 -10326 11962 -10292
rect 11896 -10434 11912 -10400
rect 11946 -10434 11962 -10400
rect 11777 -10520 11783 -10484
rect 11817 -10520 11822 -10484
rect 11777 -10554 11822 -10520
rect 11777 -10590 11783 -10554
rect 11817 -10590 11822 -10554
rect 11777 -10624 11822 -10590
rect 11777 -10660 11783 -10624
rect 11817 -10660 11822 -10624
rect 11777 -10902 11822 -10660
rect 12035 -10484 12080 -10242
rect 12292 -10066 12337 -9825
rect 12552 -9648 12597 -9604
rect 12552 -9684 12557 -9648
rect 12591 -9684 12597 -9648
rect 12552 -9718 12597 -9684
rect 12552 -9754 12557 -9718
rect 12591 -9754 12597 -9718
rect 12552 -9788 12597 -9754
rect 12552 -9824 12557 -9788
rect 12591 -9824 12597 -9788
rect 12412 -9908 12428 -9874
rect 12462 -9908 12478 -9874
rect 12412 -10016 12428 -9982
rect 12462 -10016 12478 -9982
rect 12292 -10102 12299 -10066
rect 12333 -10102 12337 -10066
rect 12292 -10136 12337 -10102
rect 12292 -10172 12299 -10136
rect 12333 -10172 12337 -10136
rect 12292 -10207 12337 -10172
rect 12292 -10243 12299 -10207
rect 12333 -10243 12337 -10207
rect 12154 -10326 12170 -10292
rect 12204 -10326 12220 -10292
rect 12154 -10434 12170 -10400
rect 12204 -10434 12220 -10400
rect 12035 -10520 12041 -10484
rect 12075 -10520 12080 -10484
rect 12035 -10554 12080 -10520
rect 12035 -10590 12041 -10554
rect 12075 -10590 12080 -10554
rect 12035 -10624 12080 -10590
rect 12035 -10660 12041 -10624
rect 12075 -10660 12080 -10624
rect 11896 -10744 11912 -10710
rect 11946 -10744 11962 -10710
rect 11896 -10852 11912 -10818
rect 11946 -10852 11962 -10818
rect 11777 -10938 11783 -10902
rect 11817 -10938 11822 -10902
rect 11777 -10972 11822 -10938
rect 11777 -11008 11783 -10972
rect 11817 -11008 11822 -10972
rect 11777 -11042 11822 -11008
rect 11777 -11078 11783 -11042
rect 11817 -11078 11822 -11042
rect 11777 -11320 11822 -11078
rect 12035 -10902 12080 -10660
rect 12292 -10484 12337 -10243
rect 12552 -10066 12597 -9824
rect 12810 -9648 12855 -9604
rect 12810 -9684 12815 -9648
rect 12849 -9684 12855 -9648
rect 12810 -9718 12855 -9684
rect 12810 -9754 12815 -9718
rect 12849 -9754 12855 -9718
rect 12810 -9788 12855 -9754
rect 12810 -9824 12815 -9788
rect 12849 -9824 12855 -9788
rect 12670 -9908 12686 -9874
rect 12720 -9908 12736 -9874
rect 12670 -10016 12686 -9982
rect 12720 -10016 12736 -9982
rect 12552 -10102 12557 -10066
rect 12591 -10102 12597 -10066
rect 12552 -10136 12597 -10102
rect 12552 -10172 12557 -10136
rect 12591 -10172 12597 -10136
rect 12552 -10206 12597 -10172
rect 12552 -10242 12557 -10206
rect 12591 -10242 12597 -10206
rect 12412 -10326 12428 -10292
rect 12462 -10326 12478 -10292
rect 12412 -10434 12428 -10400
rect 12462 -10434 12478 -10400
rect 12292 -10520 12299 -10484
rect 12333 -10520 12337 -10484
rect 12292 -10554 12337 -10520
rect 12292 -10590 12299 -10554
rect 12333 -10590 12337 -10554
rect 12292 -10625 12337 -10590
rect 12292 -10661 12299 -10625
rect 12333 -10661 12337 -10625
rect 12154 -10744 12170 -10710
rect 12204 -10744 12220 -10710
rect 12154 -10852 12170 -10818
rect 12204 -10852 12220 -10818
rect 12035 -10938 12041 -10902
rect 12075 -10938 12080 -10902
rect 12035 -10972 12080 -10938
rect 12035 -11008 12041 -10972
rect 12075 -11008 12080 -10972
rect 12035 -11042 12080 -11008
rect 12035 -11078 12041 -11042
rect 12075 -11078 12080 -11042
rect 11896 -11162 11912 -11128
rect 11946 -11162 11962 -11128
rect 11896 -11270 11912 -11236
rect 11946 -11270 11962 -11236
rect 11777 -11356 11783 -11320
rect 11817 -11356 11822 -11320
rect 11777 -11390 11822 -11356
rect 11777 -11426 11783 -11390
rect 11817 -11426 11822 -11390
rect 11777 -11460 11822 -11426
rect 11777 -11496 11783 -11460
rect 11817 -11496 11822 -11460
rect 11777 -11738 11822 -11496
rect 12035 -11320 12080 -11078
rect 12292 -10902 12337 -10661
rect 12552 -10484 12597 -10242
rect 12810 -10066 12855 -9824
rect 13067 -9648 13112 -9604
rect 13067 -9684 13073 -9648
rect 13107 -9684 13112 -9648
rect 13067 -9718 13112 -9684
rect 13067 -9754 13073 -9718
rect 13107 -9754 13112 -9718
rect 13067 -9788 13112 -9754
rect 13067 -9824 13073 -9788
rect 13107 -9824 13112 -9788
rect 12928 -9908 12944 -9874
rect 12978 -9908 12994 -9874
rect 12928 -10016 12944 -9982
rect 12978 -10016 12994 -9982
rect 12810 -10102 12815 -10066
rect 12849 -10102 12855 -10066
rect 12810 -10136 12855 -10102
rect 12810 -10172 12815 -10136
rect 12849 -10172 12855 -10136
rect 12810 -10206 12855 -10172
rect 12810 -10242 12815 -10206
rect 12849 -10242 12855 -10206
rect 12670 -10326 12686 -10292
rect 12720 -10326 12736 -10292
rect 12670 -10434 12686 -10400
rect 12720 -10434 12736 -10400
rect 12552 -10520 12557 -10484
rect 12591 -10520 12597 -10484
rect 12552 -10554 12597 -10520
rect 12552 -10590 12557 -10554
rect 12591 -10590 12597 -10554
rect 12552 -10624 12597 -10590
rect 12552 -10660 12557 -10624
rect 12591 -10660 12597 -10624
rect 12412 -10744 12428 -10710
rect 12462 -10744 12478 -10710
rect 12412 -10852 12428 -10818
rect 12462 -10852 12478 -10818
rect 12292 -10938 12299 -10902
rect 12333 -10938 12337 -10902
rect 12292 -10972 12337 -10938
rect 12292 -11008 12299 -10972
rect 12333 -11008 12337 -10972
rect 12292 -11043 12337 -11008
rect 12292 -11079 12299 -11043
rect 12333 -11079 12337 -11043
rect 12154 -11162 12170 -11128
rect 12204 -11162 12220 -11128
rect 12154 -11270 12170 -11236
rect 12204 -11270 12220 -11236
rect 12035 -11356 12041 -11320
rect 12075 -11356 12080 -11320
rect 12035 -11390 12080 -11356
rect 12035 -11426 12041 -11390
rect 12075 -11426 12080 -11390
rect 12035 -11460 12080 -11426
rect 12035 -11496 12041 -11460
rect 12075 -11496 12080 -11460
rect 11896 -11580 11912 -11546
rect 11946 -11580 11962 -11546
rect 11896 -11688 11912 -11654
rect 11946 -11688 11962 -11654
rect 11777 -11774 11783 -11738
rect 11817 -11774 11822 -11738
rect 11777 -11808 11822 -11774
rect 11777 -11844 11783 -11808
rect 11817 -11844 11822 -11808
rect 11777 -11878 11822 -11844
rect 11777 -11914 11783 -11878
rect 11817 -11914 11822 -11878
rect 11777 -12156 11822 -11914
rect 12035 -11738 12080 -11496
rect 12292 -11320 12337 -11079
rect 12552 -10902 12597 -10660
rect 12810 -10484 12855 -10242
rect 13067 -10066 13112 -9824
rect 13324 -9648 13369 -9604
rect 13324 -9684 13331 -9648
rect 13365 -9684 13369 -9648
rect 13324 -9718 13369 -9684
rect 13324 -9754 13331 -9718
rect 13365 -9754 13369 -9718
rect 13324 -9788 13369 -9754
rect 13324 -9824 13331 -9788
rect 13365 -9824 13369 -9788
rect 13186 -9908 13202 -9874
rect 13236 -9908 13252 -9874
rect 13186 -10016 13202 -9982
rect 13236 -10016 13252 -9982
rect 13067 -10102 13073 -10066
rect 13107 -10102 13112 -10066
rect 13067 -10136 13112 -10102
rect 13067 -10172 13073 -10136
rect 13107 -10172 13112 -10136
rect 13067 -10206 13112 -10172
rect 13067 -10242 13073 -10206
rect 13107 -10242 13112 -10206
rect 12928 -10326 12944 -10292
rect 12978 -10326 12994 -10292
rect 12928 -10434 12944 -10400
rect 12978 -10434 12994 -10400
rect 12810 -10520 12815 -10484
rect 12849 -10520 12855 -10484
rect 12810 -10554 12855 -10520
rect 12810 -10590 12815 -10554
rect 12849 -10590 12855 -10554
rect 12810 -10624 12855 -10590
rect 12810 -10660 12815 -10624
rect 12849 -10660 12855 -10624
rect 12670 -10744 12686 -10710
rect 12720 -10744 12736 -10710
rect 12670 -10852 12686 -10818
rect 12720 -10852 12736 -10818
rect 12552 -10938 12557 -10902
rect 12591 -10938 12597 -10902
rect 12552 -10972 12597 -10938
rect 12552 -11008 12557 -10972
rect 12591 -11008 12597 -10972
rect 12552 -11042 12597 -11008
rect 12552 -11078 12557 -11042
rect 12591 -11078 12597 -11042
rect 12412 -11162 12428 -11128
rect 12462 -11162 12478 -11128
rect 12412 -11270 12428 -11236
rect 12462 -11270 12478 -11236
rect 12292 -11356 12299 -11320
rect 12333 -11356 12337 -11320
rect 12292 -11390 12337 -11356
rect 12292 -11426 12299 -11390
rect 12333 -11426 12337 -11390
rect 12292 -11461 12337 -11426
rect 12292 -11497 12299 -11461
rect 12333 -11497 12337 -11461
rect 12154 -11580 12170 -11546
rect 12204 -11580 12220 -11546
rect 12154 -11688 12170 -11654
rect 12204 -11688 12220 -11654
rect 12035 -11774 12041 -11738
rect 12075 -11774 12080 -11738
rect 12035 -11808 12080 -11774
rect 12035 -11844 12041 -11808
rect 12075 -11844 12080 -11808
rect 12035 -11878 12080 -11844
rect 12035 -11914 12041 -11878
rect 12075 -11914 12080 -11878
rect 11896 -11998 11912 -11964
rect 11946 -11998 11962 -11964
rect 11896 -12106 11912 -12072
rect 11946 -12106 11962 -12072
rect 11777 -12192 11783 -12156
rect 11817 -12192 11822 -12156
rect 11777 -12226 11822 -12192
rect 11777 -12262 11783 -12226
rect 11817 -12262 11822 -12226
rect 11777 -12296 11822 -12262
rect 11777 -12332 11783 -12296
rect 11817 -12332 11822 -12296
rect 11777 -12574 11822 -12332
rect 12035 -12156 12080 -11914
rect 12292 -11738 12337 -11497
rect 12552 -11320 12597 -11078
rect 12810 -10902 12855 -10660
rect 13067 -10484 13112 -10242
rect 13324 -10066 13369 -9824
rect 13583 -9648 13628 -9604
rect 13583 -9684 13589 -9648
rect 13623 -9684 13628 -9648
rect 13583 -9718 13628 -9684
rect 13583 -9754 13589 -9718
rect 13623 -9754 13628 -9718
rect 13583 -9788 13628 -9754
rect 13583 -9824 13589 -9788
rect 13623 -9824 13628 -9788
rect 13444 -9908 13460 -9874
rect 13494 -9908 13510 -9874
rect 13444 -10016 13460 -9982
rect 13494 -10016 13510 -9982
rect 13324 -10102 13331 -10066
rect 13365 -10102 13369 -10066
rect 13324 -10136 13369 -10102
rect 13324 -10172 13331 -10136
rect 13365 -10172 13369 -10136
rect 13324 -10206 13369 -10172
rect 13324 -10242 13331 -10206
rect 13365 -10242 13369 -10206
rect 13186 -10326 13202 -10292
rect 13236 -10326 13252 -10292
rect 13186 -10434 13202 -10400
rect 13236 -10434 13252 -10400
rect 13067 -10520 13073 -10484
rect 13107 -10520 13112 -10484
rect 13067 -10554 13112 -10520
rect 13067 -10590 13073 -10554
rect 13107 -10590 13112 -10554
rect 13067 -10624 13112 -10590
rect 13067 -10660 13073 -10624
rect 13107 -10660 13112 -10624
rect 12928 -10744 12944 -10710
rect 12978 -10744 12994 -10710
rect 12928 -10852 12944 -10818
rect 12978 -10852 12994 -10818
rect 12810 -10938 12815 -10902
rect 12849 -10938 12855 -10902
rect 12810 -10972 12855 -10938
rect 12810 -11008 12815 -10972
rect 12849 -11008 12855 -10972
rect 12810 -11042 12855 -11008
rect 12810 -11078 12815 -11042
rect 12849 -11078 12855 -11042
rect 12670 -11162 12686 -11128
rect 12720 -11162 12736 -11128
rect 12670 -11270 12686 -11236
rect 12720 -11270 12736 -11236
rect 12552 -11356 12557 -11320
rect 12591 -11356 12597 -11320
rect 12552 -11390 12597 -11356
rect 12552 -11426 12557 -11390
rect 12591 -11426 12597 -11390
rect 12552 -11460 12597 -11426
rect 12552 -11496 12557 -11460
rect 12591 -11496 12597 -11460
rect 12412 -11580 12428 -11546
rect 12462 -11580 12478 -11546
rect 12412 -11688 12428 -11654
rect 12462 -11688 12478 -11654
rect 12292 -11774 12299 -11738
rect 12333 -11774 12337 -11738
rect 12292 -11808 12337 -11774
rect 12292 -11844 12299 -11808
rect 12333 -11844 12337 -11808
rect 12292 -11879 12337 -11844
rect 12292 -11915 12299 -11879
rect 12333 -11915 12337 -11879
rect 12154 -11998 12170 -11964
rect 12204 -11998 12220 -11964
rect 12154 -12106 12170 -12072
rect 12204 -12106 12220 -12072
rect 12035 -12192 12041 -12156
rect 12075 -12192 12080 -12156
rect 12035 -12226 12080 -12192
rect 12035 -12262 12041 -12226
rect 12075 -12262 12080 -12226
rect 12035 -12296 12080 -12262
rect 12035 -12332 12041 -12296
rect 12075 -12332 12080 -12296
rect 11896 -12416 11912 -12382
rect 11946 -12416 11962 -12382
rect 12035 -12450 12080 -12332
rect 12292 -12156 12337 -11915
rect 12552 -11738 12597 -11496
rect 12810 -11320 12855 -11078
rect 13067 -10902 13112 -10660
rect 13324 -10484 13369 -10242
rect 13583 -10066 13628 -9824
rect 13841 -9648 13886 -9462
rect 16500 -9463 16549 -9461
rect 14559 -9597 14575 -9563
rect 14609 -9597 14625 -9563
rect 14817 -9597 14833 -9563
rect 14867 -9597 14883 -9563
rect 15075 -9597 15091 -9563
rect 15125 -9597 15141 -9563
rect 15333 -9597 15349 -9563
rect 15383 -9597 15399 -9563
rect 15591 -9597 15607 -9563
rect 15641 -9597 15657 -9563
rect 15849 -9597 15865 -9563
rect 15899 -9597 15915 -9563
rect 16107 -9597 16123 -9563
rect 16157 -9597 16173 -9563
rect 16365 -9597 16381 -9563
rect 16415 -9597 16431 -9563
rect 13841 -9684 13847 -9648
rect 13881 -9684 13886 -9648
rect 13841 -9718 13886 -9684
rect 13841 -9754 13847 -9718
rect 13881 -9754 13886 -9718
rect 13841 -9788 13886 -9754
rect 13841 -9824 13847 -9788
rect 13881 -9824 13886 -9788
rect 13702 -9908 13718 -9874
rect 13752 -9908 13768 -9874
rect 13702 -10016 13718 -9982
rect 13752 -10016 13768 -9982
rect 13583 -10102 13589 -10066
rect 13623 -10102 13628 -10066
rect 13583 -10136 13628 -10102
rect 13583 -10172 13589 -10136
rect 13623 -10172 13628 -10136
rect 13583 -10206 13628 -10172
rect 13583 -10242 13589 -10206
rect 13623 -10242 13628 -10206
rect 13444 -10326 13460 -10292
rect 13494 -10326 13510 -10292
rect 13444 -10434 13460 -10400
rect 13494 -10434 13510 -10400
rect 13324 -10520 13331 -10484
rect 13365 -10520 13369 -10484
rect 13324 -10554 13369 -10520
rect 13324 -10590 13331 -10554
rect 13365 -10590 13369 -10554
rect 13324 -10624 13369 -10590
rect 13324 -10660 13331 -10624
rect 13365 -10660 13369 -10624
rect 13186 -10744 13202 -10710
rect 13236 -10744 13252 -10710
rect 13186 -10852 13202 -10818
rect 13236 -10852 13252 -10818
rect 13067 -10938 13073 -10902
rect 13107 -10938 13112 -10902
rect 13067 -10972 13112 -10938
rect 13067 -11008 13073 -10972
rect 13107 -11008 13112 -10972
rect 13067 -11042 13112 -11008
rect 13067 -11078 13073 -11042
rect 13107 -11078 13112 -11042
rect 12928 -11162 12944 -11128
rect 12978 -11162 12994 -11128
rect 12928 -11270 12944 -11236
rect 12978 -11270 12994 -11236
rect 12810 -11356 12815 -11320
rect 12849 -11356 12855 -11320
rect 12810 -11390 12855 -11356
rect 12810 -11426 12815 -11390
rect 12849 -11426 12855 -11390
rect 12810 -11460 12855 -11426
rect 12810 -11496 12815 -11460
rect 12849 -11496 12855 -11460
rect 12670 -11580 12686 -11546
rect 12720 -11580 12736 -11546
rect 12670 -11688 12686 -11654
rect 12720 -11688 12736 -11654
rect 12552 -11774 12557 -11738
rect 12591 -11774 12597 -11738
rect 12552 -11808 12597 -11774
rect 12552 -11844 12557 -11808
rect 12591 -11844 12597 -11808
rect 12552 -11878 12597 -11844
rect 12552 -11914 12557 -11878
rect 12591 -11914 12597 -11878
rect 12412 -11998 12428 -11964
rect 12462 -11998 12478 -11964
rect 12412 -12106 12428 -12072
rect 12462 -12106 12478 -12072
rect 12292 -12192 12299 -12156
rect 12333 -12192 12337 -12156
rect 12292 -12226 12337 -12192
rect 12292 -12262 12299 -12226
rect 12333 -12262 12337 -12226
rect 12292 -12297 12337 -12262
rect 12292 -12333 12299 -12297
rect 12333 -12333 12337 -12297
rect 12154 -12416 12170 -12382
rect 12204 -12416 12220 -12382
rect 12292 -12450 12337 -12333
rect 12552 -12156 12597 -11914
rect 12810 -11738 12855 -11496
rect 13067 -11320 13112 -11078
rect 13324 -10902 13369 -10660
rect 13583 -10484 13628 -10242
rect 13841 -10066 13886 -9824
rect 13841 -10102 13847 -10066
rect 13881 -10102 13886 -10066
rect 13841 -10136 13886 -10102
rect 13841 -10172 13847 -10136
rect 13881 -10172 13886 -10136
rect 13841 -10206 13886 -10172
rect 13841 -10242 13847 -10206
rect 13881 -10242 13886 -10206
rect 13702 -10326 13718 -10292
rect 13752 -10326 13768 -10292
rect 13702 -10434 13718 -10400
rect 13752 -10434 13768 -10400
rect 13583 -10520 13589 -10484
rect 13623 -10520 13628 -10484
rect 13583 -10554 13628 -10520
rect 13583 -10590 13589 -10554
rect 13623 -10590 13628 -10554
rect 13583 -10624 13628 -10590
rect 13583 -10660 13589 -10624
rect 13623 -10660 13628 -10624
rect 13444 -10744 13460 -10710
rect 13494 -10744 13510 -10710
rect 13444 -10852 13460 -10818
rect 13494 -10852 13510 -10818
rect 13324 -10938 13331 -10902
rect 13365 -10938 13369 -10902
rect 13324 -10972 13369 -10938
rect 13324 -11008 13331 -10972
rect 13365 -11008 13369 -10972
rect 13324 -11042 13369 -11008
rect 13324 -11078 13331 -11042
rect 13365 -11078 13369 -11042
rect 13186 -11162 13202 -11128
rect 13236 -11162 13252 -11128
rect 13186 -11270 13202 -11236
rect 13236 -11270 13252 -11236
rect 13067 -11356 13073 -11320
rect 13107 -11356 13112 -11320
rect 13067 -11390 13112 -11356
rect 13067 -11426 13073 -11390
rect 13107 -11426 13112 -11390
rect 13067 -11460 13112 -11426
rect 13067 -11496 13073 -11460
rect 13107 -11496 13112 -11460
rect 12928 -11580 12944 -11546
rect 12978 -11580 12994 -11546
rect 12928 -11688 12944 -11654
rect 12978 -11688 12994 -11654
rect 12810 -11774 12815 -11738
rect 12849 -11774 12855 -11738
rect 12810 -11808 12855 -11774
rect 12810 -11844 12815 -11808
rect 12849 -11844 12855 -11808
rect 12810 -11878 12855 -11844
rect 12810 -11914 12815 -11878
rect 12849 -11914 12855 -11878
rect 12670 -11998 12686 -11964
rect 12720 -11998 12736 -11964
rect 12670 -12106 12686 -12072
rect 12720 -12106 12736 -12072
rect 12552 -12192 12557 -12156
rect 12591 -12192 12597 -12156
rect 12552 -12226 12597 -12192
rect 12552 -12262 12557 -12226
rect 12591 -12262 12597 -12226
rect 12552 -12296 12597 -12262
rect 12552 -12332 12557 -12296
rect 12591 -12332 12597 -12296
rect 12412 -12416 12428 -12382
rect 12462 -12416 12478 -12382
rect 12552 -12450 12597 -12332
rect 12810 -12156 12855 -11914
rect 13067 -11738 13112 -11496
rect 13324 -11320 13369 -11078
rect 13583 -10902 13628 -10660
rect 13841 -10484 13886 -10242
rect 13841 -10520 13847 -10484
rect 13881 -10520 13886 -10484
rect 13841 -10554 13886 -10520
rect 13841 -10590 13847 -10554
rect 13881 -10590 13886 -10554
rect 13841 -10624 13886 -10590
rect 13841 -10660 13847 -10624
rect 13881 -10660 13886 -10624
rect 13702 -10744 13718 -10710
rect 13752 -10744 13768 -10710
rect 13702 -10852 13718 -10818
rect 13752 -10852 13768 -10818
rect 13583 -10938 13589 -10902
rect 13623 -10938 13628 -10902
rect 13583 -10972 13628 -10938
rect 13583 -11008 13589 -10972
rect 13623 -11008 13628 -10972
rect 13583 -11042 13628 -11008
rect 13583 -11078 13589 -11042
rect 13623 -11078 13628 -11042
rect 13444 -11162 13460 -11128
rect 13494 -11162 13510 -11128
rect 13444 -11270 13460 -11236
rect 13494 -11270 13510 -11236
rect 13324 -11356 13331 -11320
rect 13365 -11356 13369 -11320
rect 13324 -11390 13369 -11356
rect 13324 -11426 13331 -11390
rect 13365 -11426 13369 -11390
rect 13324 -11460 13369 -11426
rect 13324 -11496 13331 -11460
rect 13365 -11496 13369 -11460
rect 13186 -11580 13202 -11546
rect 13236 -11580 13252 -11546
rect 13186 -11688 13202 -11654
rect 13236 -11688 13252 -11654
rect 13067 -11774 13073 -11738
rect 13107 -11774 13112 -11738
rect 13067 -11808 13112 -11774
rect 13067 -11844 13073 -11808
rect 13107 -11844 13112 -11808
rect 13067 -11878 13112 -11844
rect 13067 -11914 13073 -11878
rect 13107 -11914 13112 -11878
rect 12928 -11998 12944 -11964
rect 12978 -11998 12994 -11964
rect 12928 -12106 12944 -12072
rect 12978 -12106 12994 -12072
rect 12810 -12192 12815 -12156
rect 12849 -12192 12855 -12156
rect 12810 -12226 12855 -12192
rect 12810 -12262 12815 -12226
rect 12849 -12262 12855 -12226
rect 12810 -12296 12855 -12262
rect 12810 -12332 12815 -12296
rect 12849 -12332 12855 -12296
rect 12670 -12416 12686 -12382
rect 12720 -12416 12736 -12382
rect 12810 -12450 12855 -12332
rect 13067 -12156 13112 -11914
rect 13324 -11738 13369 -11496
rect 13583 -11320 13628 -11078
rect 13841 -10902 13886 -10660
rect 13841 -10938 13847 -10902
rect 13881 -10938 13886 -10902
rect 13841 -10972 13886 -10938
rect 13841 -11008 13847 -10972
rect 13881 -11008 13886 -10972
rect 13841 -11042 13886 -11008
rect 13841 -11078 13847 -11042
rect 13881 -11078 13886 -11042
rect 13702 -11162 13718 -11128
rect 13752 -11162 13768 -11128
rect 13702 -11270 13718 -11236
rect 13752 -11270 13768 -11236
rect 13583 -11356 13589 -11320
rect 13623 -11356 13628 -11320
rect 13583 -11390 13628 -11356
rect 13583 -11426 13589 -11390
rect 13623 -11426 13628 -11390
rect 13583 -11460 13628 -11426
rect 13583 -11496 13589 -11460
rect 13623 -11496 13628 -11460
rect 13444 -11580 13460 -11546
rect 13494 -11580 13510 -11546
rect 13444 -11688 13460 -11654
rect 13494 -11688 13510 -11654
rect 13324 -11774 13331 -11738
rect 13365 -11774 13369 -11738
rect 13324 -11808 13369 -11774
rect 13324 -11844 13331 -11808
rect 13365 -11844 13369 -11808
rect 13324 -11878 13369 -11844
rect 13324 -11914 13331 -11878
rect 13365 -11914 13369 -11878
rect 13186 -11998 13202 -11964
rect 13236 -11998 13252 -11964
rect 13186 -12106 13202 -12072
rect 13236 -12106 13252 -12072
rect 13067 -12192 13073 -12156
rect 13107 -12192 13112 -12156
rect 13067 -12226 13112 -12192
rect 13067 -12262 13073 -12226
rect 13107 -12262 13112 -12226
rect 13067 -12296 13112 -12262
rect 13067 -12332 13073 -12296
rect 13107 -12332 13112 -12296
rect 12928 -12416 12944 -12382
rect 12978 -12416 12994 -12382
rect 13067 -12450 13112 -12332
rect 13324 -12156 13369 -11914
rect 13583 -11738 13628 -11496
rect 13841 -11320 13886 -11078
rect 13841 -11356 13847 -11320
rect 13881 -11356 13886 -11320
rect 13841 -11390 13886 -11356
rect 13841 -11426 13847 -11390
rect 13881 -11426 13886 -11390
rect 13841 -11460 13886 -11426
rect 13841 -11496 13847 -11460
rect 13881 -11496 13886 -11460
rect 13702 -11580 13718 -11546
rect 13752 -11580 13768 -11546
rect 13702 -11688 13718 -11654
rect 13752 -11688 13768 -11654
rect 13583 -11774 13589 -11738
rect 13623 -11774 13628 -11738
rect 13583 -11808 13628 -11774
rect 13583 -11844 13589 -11808
rect 13623 -11844 13628 -11808
rect 13583 -11878 13628 -11844
rect 13583 -11914 13589 -11878
rect 13623 -11914 13628 -11878
rect 13444 -11998 13460 -11964
rect 13494 -11998 13510 -11964
rect 13444 -12106 13460 -12072
rect 13494 -12106 13510 -12072
rect 13324 -12192 13331 -12156
rect 13365 -12192 13369 -12156
rect 13324 -12226 13369 -12192
rect 13324 -12262 13331 -12226
rect 13365 -12262 13369 -12226
rect 13324 -12296 13369 -12262
rect 13324 -12332 13331 -12296
rect 13365 -12332 13369 -12296
rect 13186 -12416 13202 -12382
rect 13236 -12416 13252 -12382
rect 13324 -12450 13369 -12332
rect 13583 -12156 13628 -11914
rect 13841 -11738 13886 -11496
rect 13841 -11774 13847 -11738
rect 13881 -11774 13886 -11738
rect 13841 -11808 13886 -11774
rect 13841 -11844 13847 -11808
rect 13881 -11844 13886 -11808
rect 13841 -11878 13886 -11844
rect 13841 -11914 13847 -11878
rect 13881 -11914 13886 -11878
rect 13702 -11998 13718 -11964
rect 13752 -11998 13768 -11964
rect 13702 -12106 13718 -12072
rect 13752 -12106 13768 -12072
rect 13583 -12192 13589 -12156
rect 13623 -12192 13628 -12156
rect 13583 -12226 13628 -12192
rect 13583 -12262 13589 -12226
rect 13623 -12262 13628 -12226
rect 13583 -12296 13628 -12262
rect 13583 -12332 13589 -12296
rect 13623 -12332 13628 -12296
rect 13444 -12416 13460 -12382
rect 13494 -12416 13510 -12382
rect 13583 -12450 13628 -12332
rect 13841 -12156 13886 -11914
rect 13841 -12192 13847 -12156
rect 13881 -12192 13886 -12156
rect 13841 -12226 13886 -12192
rect 13841 -12262 13847 -12226
rect 13881 -12262 13886 -12226
rect 13841 -12296 13886 -12262
rect 13841 -12332 13847 -12296
rect 13881 -12332 13886 -12296
rect 13702 -12416 13718 -12382
rect 13752 -12416 13768 -12382
rect 13841 -12450 13886 -12332
rect 14440 -9647 14485 -9603
rect 14440 -9683 14446 -9647
rect 14480 -9683 14485 -9647
rect 14440 -9717 14485 -9683
rect 14440 -9753 14446 -9717
rect 14480 -9753 14485 -9717
rect 14440 -9787 14485 -9753
rect 14440 -9823 14446 -9787
rect 14480 -9823 14485 -9787
rect 14440 -10065 14485 -9823
rect 14698 -9647 14743 -9603
rect 14698 -9683 14704 -9647
rect 14738 -9683 14743 -9647
rect 14698 -9717 14743 -9683
rect 14698 -9753 14704 -9717
rect 14738 -9753 14743 -9717
rect 14698 -9787 14743 -9753
rect 14698 -9823 14704 -9787
rect 14738 -9823 14743 -9787
rect 14559 -9907 14575 -9873
rect 14609 -9907 14625 -9873
rect 14559 -10015 14575 -9981
rect 14609 -10015 14625 -9981
rect 14440 -10101 14446 -10065
rect 14480 -10101 14485 -10065
rect 14440 -10135 14485 -10101
rect 14440 -10171 14446 -10135
rect 14480 -10171 14485 -10135
rect 14440 -10205 14485 -10171
rect 14440 -10241 14446 -10205
rect 14480 -10241 14485 -10205
rect 14440 -10483 14485 -10241
rect 14698 -10065 14743 -9823
rect 14955 -9647 15000 -9603
rect 14955 -9683 14962 -9647
rect 14996 -9683 15000 -9647
rect 14955 -9717 15000 -9683
rect 14955 -9753 14962 -9717
rect 14996 -9753 15000 -9717
rect 14955 -9788 15000 -9753
rect 14955 -9824 14962 -9788
rect 14996 -9824 15000 -9788
rect 14817 -9907 14833 -9873
rect 14867 -9907 14883 -9873
rect 14817 -10015 14833 -9981
rect 14867 -10015 14883 -9981
rect 14698 -10101 14704 -10065
rect 14738 -10101 14743 -10065
rect 14698 -10135 14743 -10101
rect 14698 -10171 14704 -10135
rect 14738 -10171 14743 -10135
rect 14698 -10205 14743 -10171
rect 14698 -10241 14704 -10205
rect 14738 -10241 14743 -10205
rect 14559 -10325 14575 -10291
rect 14609 -10325 14625 -10291
rect 14559 -10433 14575 -10399
rect 14609 -10433 14625 -10399
rect 14440 -10519 14446 -10483
rect 14480 -10519 14485 -10483
rect 14440 -10553 14485 -10519
rect 14440 -10589 14446 -10553
rect 14480 -10589 14485 -10553
rect 14440 -10623 14485 -10589
rect 14440 -10659 14446 -10623
rect 14480 -10659 14485 -10623
rect 14440 -10901 14485 -10659
rect 14698 -10483 14743 -10241
rect 14955 -10065 15000 -9824
rect 15215 -9647 15260 -9603
rect 15215 -9683 15220 -9647
rect 15254 -9683 15260 -9647
rect 15215 -9717 15260 -9683
rect 15215 -9753 15220 -9717
rect 15254 -9753 15260 -9717
rect 15215 -9787 15260 -9753
rect 15215 -9823 15220 -9787
rect 15254 -9823 15260 -9787
rect 15075 -9907 15091 -9873
rect 15125 -9907 15141 -9873
rect 15075 -10015 15091 -9981
rect 15125 -10015 15141 -9981
rect 14955 -10101 14962 -10065
rect 14996 -10101 15000 -10065
rect 14955 -10135 15000 -10101
rect 14955 -10171 14962 -10135
rect 14996 -10171 15000 -10135
rect 14955 -10206 15000 -10171
rect 14955 -10242 14962 -10206
rect 14996 -10242 15000 -10206
rect 14817 -10325 14833 -10291
rect 14867 -10325 14883 -10291
rect 14817 -10433 14833 -10399
rect 14867 -10433 14883 -10399
rect 14698 -10519 14704 -10483
rect 14738 -10519 14743 -10483
rect 14698 -10553 14743 -10519
rect 14698 -10589 14704 -10553
rect 14738 -10589 14743 -10553
rect 14698 -10623 14743 -10589
rect 14698 -10659 14704 -10623
rect 14738 -10659 14743 -10623
rect 14559 -10743 14575 -10709
rect 14609 -10743 14625 -10709
rect 14559 -10851 14575 -10817
rect 14609 -10851 14625 -10817
rect 14440 -10937 14446 -10901
rect 14480 -10937 14485 -10901
rect 14440 -10971 14485 -10937
rect 14440 -11007 14446 -10971
rect 14480 -11007 14485 -10971
rect 14440 -11041 14485 -11007
rect 14440 -11077 14446 -11041
rect 14480 -11077 14485 -11041
rect 14440 -11319 14485 -11077
rect 14698 -10901 14743 -10659
rect 14955 -10483 15000 -10242
rect 15215 -10065 15260 -9823
rect 15473 -9647 15518 -9603
rect 15473 -9683 15478 -9647
rect 15512 -9683 15518 -9647
rect 15473 -9717 15518 -9683
rect 15473 -9753 15478 -9717
rect 15512 -9753 15518 -9717
rect 15473 -9787 15518 -9753
rect 15473 -9823 15478 -9787
rect 15512 -9823 15518 -9787
rect 15333 -9907 15349 -9873
rect 15383 -9907 15399 -9873
rect 15333 -10015 15349 -9981
rect 15383 -10015 15399 -9981
rect 15215 -10101 15220 -10065
rect 15254 -10101 15260 -10065
rect 15215 -10135 15260 -10101
rect 15215 -10171 15220 -10135
rect 15254 -10171 15260 -10135
rect 15215 -10205 15260 -10171
rect 15215 -10241 15220 -10205
rect 15254 -10241 15260 -10205
rect 15075 -10325 15091 -10291
rect 15125 -10325 15141 -10291
rect 15075 -10433 15091 -10399
rect 15125 -10433 15141 -10399
rect 14955 -10519 14962 -10483
rect 14996 -10519 15000 -10483
rect 14955 -10553 15000 -10519
rect 14955 -10589 14962 -10553
rect 14996 -10589 15000 -10553
rect 14955 -10624 15000 -10589
rect 14955 -10660 14962 -10624
rect 14996 -10660 15000 -10624
rect 14817 -10743 14833 -10709
rect 14867 -10743 14883 -10709
rect 14817 -10851 14833 -10817
rect 14867 -10851 14883 -10817
rect 14698 -10937 14704 -10901
rect 14738 -10937 14743 -10901
rect 14698 -10971 14743 -10937
rect 14698 -11007 14704 -10971
rect 14738 -11007 14743 -10971
rect 14698 -11041 14743 -11007
rect 14698 -11077 14704 -11041
rect 14738 -11077 14743 -11041
rect 14559 -11161 14575 -11127
rect 14609 -11161 14625 -11127
rect 14559 -11269 14575 -11235
rect 14609 -11269 14625 -11235
rect 14440 -11355 14446 -11319
rect 14480 -11355 14485 -11319
rect 14440 -11389 14485 -11355
rect 14440 -11425 14446 -11389
rect 14480 -11425 14485 -11389
rect 14440 -11459 14485 -11425
rect 14440 -11495 14446 -11459
rect 14480 -11495 14485 -11459
rect 14440 -11737 14485 -11495
rect 14698 -11319 14743 -11077
rect 14955 -10901 15000 -10660
rect 15215 -10483 15260 -10241
rect 15473 -10065 15518 -9823
rect 15730 -9647 15775 -9603
rect 15730 -9683 15736 -9647
rect 15770 -9683 15775 -9647
rect 15730 -9717 15775 -9683
rect 15730 -9753 15736 -9717
rect 15770 -9753 15775 -9717
rect 15730 -9787 15775 -9753
rect 15730 -9823 15736 -9787
rect 15770 -9823 15775 -9787
rect 15591 -9907 15607 -9873
rect 15641 -9907 15657 -9873
rect 15591 -10015 15607 -9981
rect 15641 -10015 15657 -9981
rect 15473 -10101 15478 -10065
rect 15512 -10101 15518 -10065
rect 15473 -10135 15518 -10101
rect 15473 -10171 15478 -10135
rect 15512 -10171 15518 -10135
rect 15473 -10205 15518 -10171
rect 15473 -10241 15478 -10205
rect 15512 -10241 15518 -10205
rect 15333 -10325 15349 -10291
rect 15383 -10325 15399 -10291
rect 15333 -10433 15349 -10399
rect 15383 -10433 15399 -10399
rect 15215 -10519 15220 -10483
rect 15254 -10519 15260 -10483
rect 15215 -10553 15260 -10519
rect 15215 -10589 15220 -10553
rect 15254 -10589 15260 -10553
rect 15215 -10623 15260 -10589
rect 15215 -10659 15220 -10623
rect 15254 -10659 15260 -10623
rect 15075 -10743 15091 -10709
rect 15125 -10743 15141 -10709
rect 15075 -10851 15091 -10817
rect 15125 -10851 15141 -10817
rect 14955 -10937 14962 -10901
rect 14996 -10937 15000 -10901
rect 14955 -10971 15000 -10937
rect 14955 -11007 14962 -10971
rect 14996 -11007 15000 -10971
rect 14955 -11042 15000 -11007
rect 14955 -11078 14962 -11042
rect 14996 -11078 15000 -11042
rect 14817 -11161 14833 -11127
rect 14867 -11161 14883 -11127
rect 14817 -11269 14833 -11235
rect 14867 -11269 14883 -11235
rect 14698 -11355 14704 -11319
rect 14738 -11355 14743 -11319
rect 14698 -11389 14743 -11355
rect 14698 -11425 14704 -11389
rect 14738 -11425 14743 -11389
rect 14698 -11459 14743 -11425
rect 14698 -11495 14704 -11459
rect 14738 -11495 14743 -11459
rect 14559 -11579 14575 -11545
rect 14609 -11579 14625 -11545
rect 14559 -11687 14575 -11653
rect 14609 -11687 14625 -11653
rect 14440 -11773 14446 -11737
rect 14480 -11773 14485 -11737
rect 14440 -11807 14485 -11773
rect 14440 -11843 14446 -11807
rect 14480 -11843 14485 -11807
rect 14440 -11877 14485 -11843
rect 14440 -11913 14446 -11877
rect 14480 -11913 14485 -11877
rect 14440 -12155 14485 -11913
rect 14698 -11737 14743 -11495
rect 14955 -11319 15000 -11078
rect 15215 -10901 15260 -10659
rect 15473 -10483 15518 -10241
rect 15730 -10065 15775 -9823
rect 15987 -9647 16032 -9603
rect 15987 -9683 15994 -9647
rect 16028 -9683 16032 -9647
rect 15987 -9717 16032 -9683
rect 15987 -9753 15994 -9717
rect 16028 -9753 16032 -9717
rect 15987 -9787 16032 -9753
rect 15987 -9823 15994 -9787
rect 16028 -9823 16032 -9787
rect 15849 -9907 15865 -9873
rect 15899 -9907 15915 -9873
rect 15849 -10015 15865 -9981
rect 15899 -10015 15915 -9981
rect 15730 -10101 15736 -10065
rect 15770 -10101 15775 -10065
rect 15730 -10135 15775 -10101
rect 15730 -10171 15736 -10135
rect 15770 -10171 15775 -10135
rect 15730 -10205 15775 -10171
rect 15730 -10241 15736 -10205
rect 15770 -10241 15775 -10205
rect 15591 -10325 15607 -10291
rect 15641 -10325 15657 -10291
rect 15591 -10433 15607 -10399
rect 15641 -10433 15657 -10399
rect 15473 -10519 15478 -10483
rect 15512 -10519 15518 -10483
rect 15473 -10553 15518 -10519
rect 15473 -10589 15478 -10553
rect 15512 -10589 15518 -10553
rect 15473 -10623 15518 -10589
rect 15473 -10659 15478 -10623
rect 15512 -10659 15518 -10623
rect 15333 -10743 15349 -10709
rect 15383 -10743 15399 -10709
rect 15333 -10851 15349 -10817
rect 15383 -10851 15399 -10817
rect 15215 -10937 15220 -10901
rect 15254 -10937 15260 -10901
rect 15215 -10971 15260 -10937
rect 15215 -11007 15220 -10971
rect 15254 -11007 15260 -10971
rect 15215 -11041 15260 -11007
rect 15215 -11077 15220 -11041
rect 15254 -11077 15260 -11041
rect 15075 -11161 15091 -11127
rect 15125 -11161 15141 -11127
rect 15075 -11269 15091 -11235
rect 15125 -11269 15141 -11235
rect 14955 -11355 14962 -11319
rect 14996 -11355 15000 -11319
rect 14955 -11389 15000 -11355
rect 14955 -11425 14962 -11389
rect 14996 -11425 15000 -11389
rect 14955 -11460 15000 -11425
rect 14955 -11496 14962 -11460
rect 14996 -11496 15000 -11460
rect 14817 -11579 14833 -11545
rect 14867 -11579 14883 -11545
rect 14817 -11687 14833 -11653
rect 14867 -11687 14883 -11653
rect 14698 -11773 14704 -11737
rect 14738 -11773 14743 -11737
rect 14698 -11807 14743 -11773
rect 14698 -11843 14704 -11807
rect 14738 -11843 14743 -11807
rect 14698 -11877 14743 -11843
rect 14698 -11913 14704 -11877
rect 14738 -11913 14743 -11877
rect 14559 -11997 14575 -11963
rect 14609 -11997 14625 -11963
rect 14559 -12105 14575 -12071
rect 14609 -12105 14625 -12071
rect 14440 -12191 14446 -12155
rect 14480 -12191 14485 -12155
rect 14440 -12225 14485 -12191
rect 14440 -12261 14446 -12225
rect 14480 -12261 14485 -12225
rect 14440 -12295 14485 -12261
rect 14440 -12331 14446 -12295
rect 14480 -12331 14485 -12295
rect 14440 -12573 14485 -12331
rect 14698 -12155 14743 -11913
rect 14955 -11737 15000 -11496
rect 15215 -11319 15260 -11077
rect 15473 -10901 15518 -10659
rect 15730 -10483 15775 -10241
rect 15987 -10065 16032 -9823
rect 16246 -9647 16291 -9603
rect 16246 -9683 16252 -9647
rect 16286 -9683 16291 -9647
rect 16246 -9717 16291 -9683
rect 16246 -9753 16252 -9717
rect 16286 -9753 16291 -9717
rect 16246 -9787 16291 -9753
rect 16246 -9823 16252 -9787
rect 16286 -9823 16291 -9787
rect 16107 -9907 16123 -9873
rect 16157 -9907 16173 -9873
rect 16107 -10015 16123 -9981
rect 16157 -10015 16173 -9981
rect 15987 -10101 15994 -10065
rect 16028 -10101 16032 -10065
rect 15987 -10135 16032 -10101
rect 15987 -10171 15994 -10135
rect 16028 -10171 16032 -10135
rect 15987 -10205 16032 -10171
rect 15987 -10241 15994 -10205
rect 16028 -10241 16032 -10205
rect 15849 -10325 15865 -10291
rect 15899 -10325 15915 -10291
rect 15849 -10433 15865 -10399
rect 15899 -10433 15915 -10399
rect 15730 -10519 15736 -10483
rect 15770 -10519 15775 -10483
rect 15730 -10553 15775 -10519
rect 15730 -10589 15736 -10553
rect 15770 -10589 15775 -10553
rect 15730 -10623 15775 -10589
rect 15730 -10659 15736 -10623
rect 15770 -10659 15775 -10623
rect 15591 -10743 15607 -10709
rect 15641 -10743 15657 -10709
rect 15591 -10851 15607 -10817
rect 15641 -10851 15657 -10817
rect 15473 -10937 15478 -10901
rect 15512 -10937 15518 -10901
rect 15473 -10971 15518 -10937
rect 15473 -11007 15478 -10971
rect 15512 -11007 15518 -10971
rect 15473 -11041 15518 -11007
rect 15473 -11077 15478 -11041
rect 15512 -11077 15518 -11041
rect 15333 -11161 15349 -11127
rect 15383 -11161 15399 -11127
rect 15333 -11269 15349 -11235
rect 15383 -11269 15399 -11235
rect 15215 -11355 15220 -11319
rect 15254 -11355 15260 -11319
rect 15215 -11389 15260 -11355
rect 15215 -11425 15220 -11389
rect 15254 -11425 15260 -11389
rect 15215 -11459 15260 -11425
rect 15215 -11495 15220 -11459
rect 15254 -11495 15260 -11459
rect 15075 -11579 15091 -11545
rect 15125 -11579 15141 -11545
rect 15075 -11687 15091 -11653
rect 15125 -11687 15141 -11653
rect 14955 -11773 14962 -11737
rect 14996 -11773 15000 -11737
rect 14955 -11807 15000 -11773
rect 14955 -11843 14962 -11807
rect 14996 -11843 15000 -11807
rect 14955 -11878 15000 -11843
rect 14955 -11914 14962 -11878
rect 14996 -11914 15000 -11878
rect 14817 -11997 14833 -11963
rect 14867 -11997 14883 -11963
rect 14817 -12105 14833 -12071
rect 14867 -12105 14883 -12071
rect 14698 -12191 14704 -12155
rect 14738 -12191 14743 -12155
rect 14698 -12225 14743 -12191
rect 14698 -12261 14704 -12225
rect 14738 -12261 14743 -12225
rect 14698 -12295 14743 -12261
rect 14698 -12331 14704 -12295
rect 14738 -12331 14743 -12295
rect 14559 -12415 14575 -12381
rect 14609 -12415 14625 -12381
rect 14698 -12449 14743 -12331
rect 14955 -12155 15000 -11914
rect 15215 -11737 15260 -11495
rect 15473 -11319 15518 -11077
rect 15730 -10901 15775 -10659
rect 15987 -10483 16032 -10241
rect 16246 -10065 16291 -9823
rect 16504 -9647 16549 -9463
rect 16986 -9489 17138 -9123
rect 16504 -9683 16510 -9647
rect 16544 -9683 16549 -9647
rect 16504 -9717 16549 -9683
rect 16504 -9753 16510 -9717
rect 16544 -9753 16549 -9717
rect 16504 -9787 16549 -9753
rect 16504 -9823 16510 -9787
rect 16544 -9823 16549 -9787
rect 16365 -9907 16381 -9873
rect 16415 -9907 16431 -9873
rect 16365 -10015 16381 -9981
rect 16415 -10015 16431 -9981
rect 16246 -10101 16252 -10065
rect 16286 -10101 16291 -10065
rect 16246 -10135 16291 -10101
rect 16246 -10171 16252 -10135
rect 16286 -10171 16291 -10135
rect 16246 -10205 16291 -10171
rect 16246 -10241 16252 -10205
rect 16286 -10241 16291 -10205
rect 16107 -10325 16123 -10291
rect 16157 -10325 16173 -10291
rect 16107 -10433 16123 -10399
rect 16157 -10433 16173 -10399
rect 15987 -10519 15994 -10483
rect 16028 -10519 16032 -10483
rect 15987 -10553 16032 -10519
rect 15987 -10589 15994 -10553
rect 16028 -10589 16032 -10553
rect 15987 -10623 16032 -10589
rect 15987 -10659 15994 -10623
rect 16028 -10659 16032 -10623
rect 15849 -10743 15865 -10709
rect 15899 -10743 15915 -10709
rect 15849 -10851 15865 -10817
rect 15899 -10851 15915 -10817
rect 15730 -10937 15736 -10901
rect 15770 -10937 15775 -10901
rect 15730 -10971 15775 -10937
rect 15730 -11007 15736 -10971
rect 15770 -11007 15775 -10971
rect 15730 -11041 15775 -11007
rect 15730 -11077 15736 -11041
rect 15770 -11077 15775 -11041
rect 15591 -11161 15607 -11127
rect 15641 -11161 15657 -11127
rect 15591 -11269 15607 -11235
rect 15641 -11269 15657 -11235
rect 15473 -11355 15478 -11319
rect 15512 -11355 15518 -11319
rect 15473 -11389 15518 -11355
rect 15473 -11425 15478 -11389
rect 15512 -11425 15518 -11389
rect 15473 -11459 15518 -11425
rect 15473 -11495 15478 -11459
rect 15512 -11495 15518 -11459
rect 15333 -11579 15349 -11545
rect 15383 -11579 15399 -11545
rect 15333 -11687 15349 -11653
rect 15383 -11687 15399 -11653
rect 15215 -11773 15220 -11737
rect 15254 -11773 15260 -11737
rect 15215 -11807 15260 -11773
rect 15215 -11843 15220 -11807
rect 15254 -11843 15260 -11807
rect 15215 -11877 15260 -11843
rect 15215 -11913 15220 -11877
rect 15254 -11913 15260 -11877
rect 15075 -11997 15091 -11963
rect 15125 -11997 15141 -11963
rect 15075 -12105 15091 -12071
rect 15125 -12105 15141 -12071
rect 14955 -12191 14962 -12155
rect 14996 -12191 15000 -12155
rect 14955 -12225 15000 -12191
rect 14955 -12261 14962 -12225
rect 14996 -12261 15000 -12225
rect 14955 -12296 15000 -12261
rect 14955 -12332 14962 -12296
rect 14996 -12332 15000 -12296
rect 14817 -12415 14833 -12381
rect 14867 -12415 14883 -12381
rect 14955 -12449 15000 -12332
rect 15215 -12155 15260 -11913
rect 15473 -11737 15518 -11495
rect 15730 -11319 15775 -11077
rect 15987 -10901 16032 -10659
rect 16246 -10483 16291 -10241
rect 16504 -10065 16549 -9823
rect 16504 -10101 16510 -10065
rect 16544 -10101 16549 -10065
rect 16504 -10135 16549 -10101
rect 16504 -10171 16510 -10135
rect 16544 -10171 16549 -10135
rect 16504 -10205 16549 -10171
rect 16504 -10241 16510 -10205
rect 16544 -10241 16549 -10205
rect 16365 -10325 16381 -10291
rect 16415 -10325 16431 -10291
rect 16365 -10433 16381 -10399
rect 16415 -10433 16431 -10399
rect 16246 -10519 16252 -10483
rect 16286 -10519 16291 -10483
rect 16246 -10553 16291 -10519
rect 16246 -10589 16252 -10553
rect 16286 -10589 16291 -10553
rect 16246 -10623 16291 -10589
rect 16246 -10659 16252 -10623
rect 16286 -10659 16291 -10623
rect 16107 -10743 16123 -10709
rect 16157 -10743 16173 -10709
rect 16107 -10851 16123 -10817
rect 16157 -10851 16173 -10817
rect 15987 -10937 15994 -10901
rect 16028 -10937 16032 -10901
rect 15987 -10971 16032 -10937
rect 15987 -11007 15994 -10971
rect 16028 -11007 16032 -10971
rect 15987 -11041 16032 -11007
rect 15987 -11077 15994 -11041
rect 16028 -11077 16032 -11041
rect 15849 -11161 15865 -11127
rect 15899 -11161 15915 -11127
rect 15849 -11269 15865 -11235
rect 15899 -11269 15915 -11235
rect 15730 -11355 15736 -11319
rect 15770 -11355 15775 -11319
rect 15730 -11389 15775 -11355
rect 15730 -11425 15736 -11389
rect 15770 -11425 15775 -11389
rect 15730 -11459 15775 -11425
rect 15730 -11495 15736 -11459
rect 15770 -11495 15775 -11459
rect 15591 -11579 15607 -11545
rect 15641 -11579 15657 -11545
rect 15591 -11687 15607 -11653
rect 15641 -11687 15657 -11653
rect 15473 -11773 15478 -11737
rect 15512 -11773 15518 -11737
rect 15473 -11807 15518 -11773
rect 15473 -11843 15478 -11807
rect 15512 -11843 15518 -11807
rect 15473 -11877 15518 -11843
rect 15473 -11913 15478 -11877
rect 15512 -11913 15518 -11877
rect 15333 -11997 15349 -11963
rect 15383 -11997 15399 -11963
rect 15333 -12105 15349 -12071
rect 15383 -12105 15399 -12071
rect 15215 -12191 15220 -12155
rect 15254 -12191 15260 -12155
rect 15215 -12225 15260 -12191
rect 15215 -12261 15220 -12225
rect 15254 -12261 15260 -12225
rect 15215 -12295 15260 -12261
rect 15215 -12331 15220 -12295
rect 15254 -12331 15260 -12295
rect 15075 -12415 15091 -12381
rect 15125 -12415 15141 -12381
rect 15215 -12449 15260 -12331
rect 15473 -12155 15518 -11913
rect 15730 -11737 15775 -11495
rect 15987 -11319 16032 -11077
rect 16246 -10901 16291 -10659
rect 16504 -10483 16549 -10241
rect 16504 -10519 16510 -10483
rect 16544 -10519 16549 -10483
rect 16504 -10553 16549 -10519
rect 16504 -10589 16510 -10553
rect 16544 -10589 16549 -10553
rect 16504 -10623 16549 -10589
rect 16504 -10659 16510 -10623
rect 16544 -10659 16549 -10623
rect 16365 -10743 16381 -10709
rect 16415 -10743 16431 -10709
rect 16365 -10851 16381 -10817
rect 16415 -10851 16431 -10817
rect 16246 -10937 16252 -10901
rect 16286 -10937 16291 -10901
rect 16246 -10971 16291 -10937
rect 16246 -11007 16252 -10971
rect 16286 -11007 16291 -10971
rect 16246 -11041 16291 -11007
rect 16246 -11077 16252 -11041
rect 16286 -11077 16291 -11041
rect 16107 -11161 16123 -11127
rect 16157 -11161 16173 -11127
rect 16107 -11269 16123 -11235
rect 16157 -11269 16173 -11235
rect 15987 -11355 15994 -11319
rect 16028 -11355 16032 -11319
rect 15987 -11389 16032 -11355
rect 15987 -11425 15994 -11389
rect 16028 -11425 16032 -11389
rect 15987 -11459 16032 -11425
rect 15987 -11495 15994 -11459
rect 16028 -11495 16032 -11459
rect 15849 -11579 15865 -11545
rect 15899 -11579 15915 -11545
rect 15849 -11687 15865 -11653
rect 15899 -11687 15915 -11653
rect 15730 -11773 15736 -11737
rect 15770 -11773 15775 -11737
rect 15730 -11807 15775 -11773
rect 15730 -11843 15736 -11807
rect 15770 -11843 15775 -11807
rect 15730 -11877 15775 -11843
rect 15730 -11913 15736 -11877
rect 15770 -11913 15775 -11877
rect 15591 -11997 15607 -11963
rect 15641 -11997 15657 -11963
rect 15591 -12105 15607 -12071
rect 15641 -12105 15657 -12071
rect 15473 -12191 15478 -12155
rect 15512 -12191 15518 -12155
rect 15473 -12225 15518 -12191
rect 15473 -12261 15478 -12225
rect 15512 -12261 15518 -12225
rect 15473 -12295 15518 -12261
rect 15473 -12331 15478 -12295
rect 15512 -12331 15518 -12295
rect 15333 -12415 15349 -12381
rect 15383 -12415 15399 -12381
rect 15473 -12449 15518 -12331
rect 15730 -12155 15775 -11913
rect 15987 -11737 16032 -11495
rect 16246 -11319 16291 -11077
rect 16504 -10901 16549 -10659
rect 16504 -10937 16510 -10901
rect 16544 -10937 16549 -10901
rect 16504 -10971 16549 -10937
rect 16504 -11007 16510 -10971
rect 16544 -11007 16549 -10971
rect 16504 -11041 16549 -11007
rect 16504 -11077 16510 -11041
rect 16544 -11077 16549 -11041
rect 16365 -11161 16381 -11127
rect 16415 -11161 16431 -11127
rect 16365 -11269 16381 -11235
rect 16415 -11269 16431 -11235
rect 16246 -11355 16252 -11319
rect 16286 -11355 16291 -11319
rect 16246 -11389 16291 -11355
rect 16246 -11425 16252 -11389
rect 16286 -11425 16291 -11389
rect 16246 -11459 16291 -11425
rect 16246 -11495 16252 -11459
rect 16286 -11495 16291 -11459
rect 16107 -11579 16123 -11545
rect 16157 -11579 16173 -11545
rect 16107 -11687 16123 -11653
rect 16157 -11687 16173 -11653
rect 15987 -11773 15994 -11737
rect 16028 -11773 16032 -11737
rect 15987 -11807 16032 -11773
rect 15987 -11843 15994 -11807
rect 16028 -11843 16032 -11807
rect 15987 -11877 16032 -11843
rect 15987 -11913 15994 -11877
rect 16028 -11913 16032 -11877
rect 15849 -11997 15865 -11963
rect 15899 -11997 15915 -11963
rect 15849 -12105 15865 -12071
rect 15899 -12105 15915 -12071
rect 15730 -12191 15736 -12155
rect 15770 -12191 15775 -12155
rect 15730 -12225 15775 -12191
rect 15730 -12261 15736 -12225
rect 15770 -12261 15775 -12225
rect 15730 -12295 15775 -12261
rect 15730 -12331 15736 -12295
rect 15770 -12331 15775 -12295
rect 15591 -12415 15607 -12381
rect 15641 -12415 15657 -12381
rect 15730 -12449 15775 -12331
rect 15987 -12155 16032 -11913
rect 16246 -11737 16291 -11495
rect 16504 -11319 16549 -11077
rect 16504 -11355 16510 -11319
rect 16544 -11355 16549 -11319
rect 16504 -11389 16549 -11355
rect 16504 -11425 16510 -11389
rect 16544 -11425 16549 -11389
rect 16504 -11459 16549 -11425
rect 16504 -11495 16510 -11459
rect 16544 -11495 16549 -11459
rect 16365 -11579 16381 -11545
rect 16415 -11579 16431 -11545
rect 16365 -11687 16381 -11653
rect 16415 -11687 16431 -11653
rect 16246 -11773 16252 -11737
rect 16286 -11773 16291 -11737
rect 16246 -11807 16291 -11773
rect 16246 -11843 16252 -11807
rect 16286 -11843 16291 -11807
rect 16246 -11877 16291 -11843
rect 16246 -11913 16252 -11877
rect 16286 -11913 16291 -11877
rect 16107 -11997 16123 -11963
rect 16157 -11997 16173 -11963
rect 16107 -12105 16123 -12071
rect 16157 -12105 16173 -12071
rect 15987 -12191 15994 -12155
rect 16028 -12191 16032 -12155
rect 15987 -12225 16032 -12191
rect 15987 -12261 15994 -12225
rect 16028 -12261 16032 -12225
rect 15987 -12295 16032 -12261
rect 15987 -12331 15994 -12295
rect 16028 -12331 16032 -12295
rect 15849 -12415 15865 -12381
rect 15899 -12415 15915 -12381
rect 15987 -12449 16032 -12331
rect 16246 -12155 16291 -11913
rect 16504 -11737 16549 -11495
rect 16504 -11773 16510 -11737
rect 16544 -11773 16549 -11737
rect 16504 -11807 16549 -11773
rect 16504 -11843 16510 -11807
rect 16544 -11843 16549 -11807
rect 16504 -11877 16549 -11843
rect 16504 -11913 16510 -11877
rect 16544 -11913 16549 -11877
rect 16365 -11997 16381 -11963
rect 16415 -11997 16431 -11963
rect 16365 -12105 16381 -12071
rect 16415 -12105 16431 -12071
rect 16246 -12191 16252 -12155
rect 16286 -12191 16291 -12155
rect 16246 -12225 16291 -12191
rect 16246 -12261 16252 -12225
rect 16286 -12261 16291 -12225
rect 16246 -12295 16291 -12261
rect 16246 -12331 16252 -12295
rect 16286 -12331 16291 -12295
rect 16107 -12415 16123 -12381
rect 16157 -12415 16173 -12381
rect 16246 -12449 16291 -12331
rect 16504 -12155 16549 -11913
rect 16504 -12191 16510 -12155
rect 16544 -12191 16549 -12155
rect 16504 -12225 16549 -12191
rect 16504 -12261 16510 -12225
rect 16544 -12261 16549 -12225
rect 16504 -12295 16549 -12261
rect 16504 -12331 16510 -12295
rect 16544 -12331 16549 -12295
rect 16365 -12415 16381 -12381
rect 16415 -12415 16431 -12381
rect 16504 -12449 16549 -12331
rect 9107 -12669 10333 -12574
rect 11777 -12669 13003 -12574
rect 14440 -12668 15666 -12573
rect 9106 -12758 9122 -12724
rect 9156 -12758 9172 -12724
rect 9646 -12758 9662 -12724
rect 9696 -12758 9712 -12724
rect 10126 -12758 10137 -12724
rect 10187 -12758 10192 -12724
rect 8967 -12810 9029 -12788
rect 8967 -12844 8993 -12810
rect 9027 -12844 9029 -12810
rect 8967 -12878 9029 -12844
rect 8967 -12914 8993 -12878
rect 9027 -12914 9029 -12878
rect 8967 -12948 9029 -12914
rect 8967 -12982 8993 -12948
rect 9027 -12982 9029 -12948
rect 8967 -13024 9029 -12982
rect 9245 -12810 9313 -12790
rect 9245 -12844 9251 -12810
rect 9285 -12844 9313 -12810
rect 9245 -12878 9313 -12844
rect 9245 -12914 9251 -12878
rect 9285 -12914 9313 -12878
rect 9245 -12948 9313 -12914
rect 9245 -12982 9251 -12948
rect 9285 -12982 9313 -12948
rect 9245 -13026 9313 -12982
rect 9507 -12810 9569 -12788
rect 9507 -12844 9533 -12810
rect 9567 -12844 9569 -12810
rect 9507 -12878 9569 -12844
rect 9507 -12914 9533 -12878
rect 9567 -12914 9569 -12878
rect 9507 -12948 9569 -12914
rect 9507 -12982 9533 -12948
rect 9567 -12982 9569 -12948
rect 9507 -13024 9569 -12982
rect 9785 -12810 9853 -12790
rect 9785 -12844 9791 -12810
rect 9825 -12844 9853 -12810
rect 9785 -12878 9853 -12844
rect 9785 -12914 9791 -12878
rect 9825 -12914 9853 -12878
rect 9785 -12948 9853 -12914
rect 9785 -12982 9791 -12948
rect 9825 -12982 9853 -12948
rect 9785 -13026 9853 -12982
rect 9987 -12810 10049 -12788
rect 9987 -12844 10013 -12810
rect 10047 -12844 10049 -12810
rect 9987 -12878 10049 -12844
rect 9987 -12914 10013 -12878
rect 10047 -12914 10049 -12878
rect 9987 -12948 10049 -12914
rect 9987 -12982 10013 -12948
rect 10047 -12982 10049 -12948
rect 9106 -13068 9122 -13034
rect 9156 -13068 9172 -13034
rect 9646 -13068 9662 -13034
rect 9696 -13068 9712 -13034
rect 9987 -13153 10049 -12982
rect 10265 -12810 10333 -12669
rect 10629 -12756 10645 -12722
rect 10679 -12756 10695 -12722
rect 11139 -12746 11155 -12712
rect 11189 -12746 11205 -12712
rect 11776 -12758 11792 -12724
rect 11826 -12758 11842 -12724
rect 12316 -12758 12332 -12724
rect 12366 -12758 12382 -12724
rect 12796 -12758 12807 -12724
rect 12857 -12758 12862 -12724
rect 10265 -12844 10271 -12810
rect 10305 -12844 10333 -12810
rect 10265 -12878 10333 -12844
rect 10265 -12914 10271 -12878
rect 10305 -12914 10333 -12878
rect 10265 -12948 10333 -12914
rect 10265 -12982 10271 -12948
rect 10305 -12982 10333 -12948
rect 10265 -13026 10333 -12982
rect 10490 -12808 10552 -12786
rect 10490 -12842 10516 -12808
rect 10550 -12842 10552 -12808
rect 10490 -12876 10552 -12842
rect 10490 -12912 10516 -12876
rect 10550 -12912 10552 -12876
rect 10490 -12946 10552 -12912
rect 10490 -12980 10516 -12946
rect 10550 -12980 10552 -12946
rect 10490 -13022 10552 -12980
rect 10768 -12808 10836 -12788
rect 10768 -12842 10774 -12808
rect 10808 -12842 10836 -12808
rect 10768 -12876 10836 -12842
rect 10768 -12912 10774 -12876
rect 10808 -12912 10836 -12876
rect 10768 -12946 10836 -12912
rect 10768 -12980 10774 -12946
rect 10808 -12980 10836 -12946
rect 10768 -13024 10836 -12980
rect 11000 -12798 11062 -12776
rect 11000 -12832 11026 -12798
rect 11060 -12832 11062 -12798
rect 11000 -12866 11062 -12832
rect 11000 -12902 11026 -12866
rect 11060 -12902 11062 -12866
rect 11000 -12936 11062 -12902
rect 11000 -12970 11026 -12936
rect 11060 -12970 11062 -12936
rect 11000 -13012 11062 -12970
rect 11278 -12798 11346 -12778
rect 11278 -12832 11284 -12798
rect 11318 -12832 11346 -12798
rect 11278 -12866 11346 -12832
rect 11278 -12902 11284 -12866
rect 11318 -12902 11346 -12866
rect 11278 -12936 11346 -12902
rect 11278 -12970 11284 -12936
rect 11318 -12970 11346 -12936
rect 11278 -13014 11346 -12970
rect 11637 -12810 11699 -12788
rect 11637 -12844 11663 -12810
rect 11697 -12844 11699 -12810
rect 11637 -12878 11699 -12844
rect 11637 -12914 11663 -12878
rect 11697 -12914 11699 -12878
rect 11637 -12948 11699 -12914
rect 11637 -12982 11663 -12948
rect 11697 -12982 11699 -12948
rect 10126 -13068 10140 -13034
rect 10178 -13068 10192 -13034
rect 10629 -13066 10645 -13032
rect 10679 -13066 10695 -13032
rect 11139 -13056 11155 -13022
rect 11189 -13056 11205 -13022
rect 11637 -13024 11699 -12982
rect 11915 -12810 11983 -12790
rect 11915 -12844 11921 -12810
rect 11955 -12844 11983 -12810
rect 11915 -12878 11983 -12844
rect 11915 -12914 11921 -12878
rect 11955 -12914 11983 -12878
rect 11915 -12948 11983 -12914
rect 11915 -12982 11921 -12948
rect 11955 -12982 11983 -12948
rect 11915 -13026 11983 -12982
rect 12177 -12810 12239 -12788
rect 12177 -12844 12203 -12810
rect 12237 -12844 12239 -12810
rect 12177 -12878 12239 -12844
rect 12177 -12914 12203 -12878
rect 12237 -12914 12239 -12878
rect 12177 -12948 12239 -12914
rect 12177 -12982 12203 -12948
rect 12237 -12982 12239 -12948
rect 12177 -13024 12239 -12982
rect 12455 -12810 12523 -12790
rect 12455 -12844 12461 -12810
rect 12495 -12844 12523 -12810
rect 12455 -12878 12523 -12844
rect 12455 -12914 12461 -12878
rect 12495 -12914 12523 -12878
rect 12455 -12948 12523 -12914
rect 12455 -12982 12461 -12948
rect 12495 -12982 12523 -12948
rect 12455 -13026 12523 -12982
rect 12657 -12810 12719 -12788
rect 12657 -12844 12683 -12810
rect 12717 -12844 12719 -12810
rect 12657 -12878 12719 -12844
rect 12657 -12914 12683 -12878
rect 12717 -12914 12719 -12878
rect 12657 -12948 12719 -12914
rect 12657 -12982 12683 -12948
rect 12717 -12982 12719 -12948
rect 11776 -13068 11792 -13034
rect 11826 -13068 11842 -13034
rect 12316 -13068 12332 -13034
rect 12366 -13068 12382 -13034
rect 12657 -13094 12719 -12982
rect 12935 -12810 13003 -12669
rect 13299 -12756 13315 -12722
rect 13349 -12756 13365 -12722
rect 13809 -12746 13825 -12712
rect 13859 -12746 13875 -12712
rect 14439 -12757 14455 -12723
rect 14489 -12757 14505 -12723
rect 14979 -12757 14995 -12723
rect 15029 -12757 15045 -12723
rect 15459 -12757 15470 -12723
rect 15520 -12757 15525 -12723
rect 12935 -12844 12941 -12810
rect 12975 -12844 13003 -12810
rect 12935 -12878 13003 -12844
rect 12935 -12914 12941 -12878
rect 12975 -12914 13003 -12878
rect 12935 -12948 13003 -12914
rect 12935 -12982 12941 -12948
rect 12975 -12982 13003 -12948
rect 12935 -13026 13003 -12982
rect 13160 -12808 13222 -12786
rect 13160 -12842 13186 -12808
rect 13220 -12842 13222 -12808
rect 13160 -12876 13222 -12842
rect 13160 -12912 13186 -12876
rect 13220 -12912 13222 -12876
rect 13160 -12946 13222 -12912
rect 13160 -12980 13186 -12946
rect 13220 -12980 13222 -12946
rect 13160 -13022 13222 -12980
rect 13438 -12808 13506 -12788
rect 13438 -12842 13444 -12808
rect 13478 -12842 13506 -12808
rect 13438 -12876 13506 -12842
rect 13438 -12912 13444 -12876
rect 13478 -12912 13506 -12876
rect 13438 -12946 13506 -12912
rect 13438 -12980 13444 -12946
rect 13478 -12980 13506 -12946
rect 13438 -13024 13506 -12980
rect 13670 -12798 13732 -12776
rect 13670 -12832 13696 -12798
rect 13730 -12832 13732 -12798
rect 13670 -12866 13732 -12832
rect 13670 -12902 13696 -12866
rect 13730 -12902 13732 -12866
rect 13670 -12936 13732 -12902
rect 13670 -12970 13696 -12936
rect 13730 -12970 13732 -12936
rect 13670 -13012 13732 -12970
rect 13948 -12798 14016 -12778
rect 13948 -12832 13954 -12798
rect 13988 -12832 14016 -12798
rect 13948 -12866 14016 -12832
rect 13948 -12902 13954 -12866
rect 13988 -12902 14016 -12866
rect 13948 -12936 14016 -12902
rect 13948 -12970 13954 -12936
rect 13988 -12970 14016 -12936
rect 13948 -13014 14016 -12970
rect 14300 -12809 14362 -12787
rect 14300 -12843 14326 -12809
rect 14360 -12843 14362 -12809
rect 14300 -12877 14362 -12843
rect 14300 -12913 14326 -12877
rect 14360 -12913 14362 -12877
rect 14300 -12947 14362 -12913
rect 14300 -12981 14326 -12947
rect 14360 -12981 14362 -12947
rect 12796 -13068 12810 -13034
rect 12848 -13068 12862 -13034
rect 13299 -13066 13315 -13032
rect 13349 -13066 13365 -13032
rect 13809 -13056 13825 -13022
rect 13859 -13056 13875 -13022
rect 14300 -13023 14362 -12981
rect 14578 -12809 14646 -12789
rect 14578 -12843 14584 -12809
rect 14618 -12843 14646 -12809
rect 14578 -12877 14646 -12843
rect 14578 -12913 14584 -12877
rect 14618 -12913 14646 -12877
rect 14578 -12947 14646 -12913
rect 14578 -12981 14584 -12947
rect 14618 -12981 14646 -12947
rect 14578 -13025 14646 -12981
rect 14840 -12809 14902 -12787
rect 14840 -12843 14866 -12809
rect 14900 -12843 14902 -12809
rect 14840 -12877 14902 -12843
rect 14840 -12913 14866 -12877
rect 14900 -12913 14902 -12877
rect 14840 -12947 14902 -12913
rect 14840 -12981 14866 -12947
rect 14900 -12981 14902 -12947
rect 14840 -13023 14902 -12981
rect 15118 -12809 15186 -12789
rect 15118 -12843 15124 -12809
rect 15158 -12843 15186 -12809
rect 15118 -12877 15186 -12843
rect 15118 -12913 15124 -12877
rect 15158 -12913 15186 -12877
rect 15118 -12947 15186 -12913
rect 15118 -12981 15124 -12947
rect 15158 -12981 15186 -12947
rect 15118 -13025 15186 -12981
rect 15320 -12809 15382 -12787
rect 15320 -12843 15346 -12809
rect 15380 -12843 15382 -12809
rect 15320 -12877 15382 -12843
rect 15320 -12913 15346 -12877
rect 15380 -12913 15382 -12877
rect 15320 -12947 15382 -12913
rect 15320 -12981 15346 -12947
rect 15380 -12981 15382 -12947
rect 14439 -13067 14455 -13033
rect 14489 -13067 14505 -13033
rect 14979 -13067 14995 -13033
rect 15029 -13067 15045 -13033
rect 12656 -13153 12719 -13094
rect 15320 -13153 15382 -12981
rect 15598 -12809 15666 -12668
rect 15962 -12755 15978 -12721
rect 16012 -12755 16028 -12721
rect 16472 -12745 16488 -12711
rect 16522 -12745 16538 -12711
rect 15598 -12843 15604 -12809
rect 15638 -12843 15666 -12809
rect 15598 -12877 15666 -12843
rect 15598 -12913 15604 -12877
rect 15638 -12913 15666 -12877
rect 15598 -12947 15666 -12913
rect 15598 -12981 15604 -12947
rect 15638 -12981 15666 -12947
rect 15598 -13025 15666 -12981
rect 15823 -12807 15885 -12785
rect 15823 -12841 15849 -12807
rect 15883 -12841 15885 -12807
rect 15823 -12875 15885 -12841
rect 15823 -12911 15849 -12875
rect 15883 -12911 15885 -12875
rect 15823 -12945 15885 -12911
rect 15823 -12979 15849 -12945
rect 15883 -12979 15885 -12945
rect 15823 -13021 15885 -12979
rect 16101 -12807 16169 -12787
rect 16101 -12841 16107 -12807
rect 16141 -12841 16169 -12807
rect 16101 -12875 16169 -12841
rect 16101 -12911 16107 -12875
rect 16141 -12911 16169 -12875
rect 16101 -12945 16169 -12911
rect 16101 -12979 16107 -12945
rect 16141 -12979 16169 -12945
rect 16101 -13023 16169 -12979
rect 16333 -12797 16395 -12775
rect 16333 -12831 16359 -12797
rect 16393 -12831 16395 -12797
rect 16333 -12865 16395 -12831
rect 16333 -12901 16359 -12865
rect 16393 -12901 16395 -12865
rect 16333 -12935 16395 -12901
rect 16333 -12969 16359 -12935
rect 16393 -12969 16395 -12935
rect 16333 -13011 16395 -12969
rect 16611 -12797 16679 -12777
rect 16611 -12831 16617 -12797
rect 16651 -12831 16679 -12797
rect 16611 -12865 16679 -12831
rect 16611 -12901 16617 -12865
rect 16651 -12901 16679 -12865
rect 16611 -12935 16679 -12901
rect 16611 -12969 16617 -12935
rect 16651 -12969 16679 -12935
rect 16611 -13013 16679 -12969
rect 15459 -13067 15472 -13033
rect 15510 -13067 15525 -13033
rect 15962 -13065 15978 -13031
rect 16012 -13065 16028 -13031
rect 16472 -13055 16488 -13021
rect 16522 -13055 16538 -13021
rect 8805 -13161 16813 -13153
rect 8805 -13267 9970 -13161
rect 10076 -13267 12634 -13161
rect 12740 -13267 15296 -13161
rect 15402 -13267 16813 -13161
rect 8805 -13273 16813 -13267
rect 8484 -13374 16813 -13373
rect 16987 -13374 17137 -9489
rect 8484 -13493 17137 -13374
rect 8484 -13799 8634 -13493
rect 8484 -14133 8636 -13799
rect 8484 -19151 8634 -14133
rect 9312 -14243 9584 -14213
rect 9312 -14281 9408 -14243
rect 9474 -14281 9584 -14243
rect 9312 -14367 9584 -14281
rect 9312 -14369 9516 -14367
rect 9312 -14405 9330 -14369
rect 9368 -14403 9516 -14369
rect 9554 -14403 9584 -14367
rect 9368 -14405 9584 -14403
rect 9312 -14441 9584 -14405
rect 9664 -14285 9728 -13493
rect 10698 -14244 10970 -14214
rect 10036 -14284 10052 -14250
rect 10206 -14284 10222 -14250
rect 10698 -14282 10794 -14244
rect 10860 -14282 10970 -14244
rect 9664 -14369 9720 -14285
rect 10544 -14316 10608 -14315
rect 9664 -14403 9683 -14369
rect 9717 -14403 9720 -14369
rect 9664 -14441 9720 -14403
rect 10539 -14369 10608 -14316
rect 10539 -14403 10541 -14369
rect 10575 -14403 10608 -14369
rect 10539 -14435 10608 -14403
rect 10036 -14522 10052 -14488
rect 10206 -14522 10222 -14488
rect 10536 -14969 10608 -14435
rect 10698 -14368 10970 -14282
rect 10698 -14370 10902 -14368
rect 10698 -14406 10716 -14370
rect 10754 -14404 10902 -14370
rect 10940 -14404 10970 -14368
rect 10754 -14406 10970 -14404
rect 10698 -14442 10970 -14406
rect 11068 -14244 11340 -14214
rect 11068 -14282 11164 -14244
rect 11230 -14282 11340 -14244
rect 11068 -14368 11340 -14282
rect 11068 -14370 11272 -14368
rect 11068 -14406 11086 -14370
rect 11124 -14404 11272 -14370
rect 11310 -14404 11340 -14368
rect 11124 -14406 11340 -14404
rect 11068 -14442 11340 -14406
rect 11490 -14244 11762 -14214
rect 11490 -14282 11586 -14244
rect 11652 -14282 11762 -14244
rect 11490 -14368 11762 -14282
rect 11490 -14370 11694 -14368
rect 11490 -14406 11508 -14370
rect 11546 -14404 11694 -14370
rect 11732 -14404 11762 -14368
rect 11546 -14406 11762 -14404
rect 11490 -14442 11762 -14406
rect 11912 -14244 12184 -14214
rect 11912 -14282 12008 -14244
rect 12074 -14282 12184 -14244
rect 11912 -14368 12184 -14282
rect 11912 -14370 12116 -14368
rect 11912 -14406 11930 -14370
rect 11968 -14404 12116 -14370
rect 12154 -14404 12184 -14368
rect 11968 -14406 12184 -14404
rect 11912 -14442 12184 -14406
rect 12334 -14299 12398 -13493
rect 13412 -14240 13684 -14212
rect 12713 -14284 12729 -14250
rect 12883 -14284 12899 -14250
rect 13412 -14278 13508 -14240
rect 13574 -14278 13684 -14240
rect 12334 -14369 12396 -14299
rect 12334 -14403 12360 -14369
rect 12394 -14403 12396 -14369
rect 12334 -14445 12396 -14403
rect 13216 -14369 13289 -14301
rect 13216 -14403 13218 -14369
rect 13252 -14403 13289 -14369
rect 13216 -14447 13289 -14403
rect 13412 -14364 13684 -14278
rect 13412 -14366 13616 -14364
rect 13412 -14402 13430 -14366
rect 13468 -14400 13616 -14366
rect 13654 -14400 13684 -14364
rect 13468 -14402 13684 -14400
rect 13412 -14438 13684 -14402
rect 13782 -14240 14054 -14212
rect 13782 -14278 13878 -14240
rect 13944 -14278 14054 -14240
rect 13782 -14364 14054 -14278
rect 13782 -14366 13986 -14364
rect 13782 -14402 13800 -14366
rect 13838 -14400 13986 -14366
rect 14024 -14400 14054 -14364
rect 13838 -14402 14054 -14400
rect 13782 -14438 14054 -14402
rect 14204 -14240 14476 -14212
rect 14204 -14278 14300 -14240
rect 14366 -14278 14476 -14240
rect 14204 -14364 14476 -14278
rect 14204 -14366 14408 -14364
rect 14204 -14402 14222 -14366
rect 14260 -14400 14408 -14366
rect 14446 -14400 14476 -14364
rect 14260 -14402 14476 -14400
rect 14204 -14438 14476 -14402
rect 14626 -14240 14898 -14212
rect 14626 -14278 14722 -14240
rect 14788 -14278 14898 -14240
rect 14626 -14364 14898 -14278
rect 14996 -14347 15060 -13493
rect 16540 -13494 17137 -13493
rect 16987 -13783 17137 -13494
rect 16986 -14165 17138 -13783
rect 16010 -14243 16282 -14213
rect 15377 -14283 15393 -14249
rect 15547 -14283 15563 -14249
rect 16010 -14281 16106 -14243
rect 16172 -14281 16282 -14243
rect 14626 -14366 14830 -14364
rect 14626 -14402 14644 -14366
rect 14682 -14400 14830 -14366
rect 14868 -14400 14898 -14364
rect 14682 -14402 14898 -14400
rect 14626 -14438 14898 -14402
rect 14997 -14368 15060 -14347
rect 14997 -14402 15024 -14368
rect 15058 -14402 15060 -14368
rect 14997 -14425 15060 -14402
rect 15880 -14368 15934 -14297
rect 15880 -14402 15882 -14368
rect 15916 -14402 15934 -14368
rect 12713 -14522 12729 -14488
rect 12883 -14522 12899 -14488
rect 8830 -15005 11218 -14969
rect 8824 -15007 11218 -15005
rect 8824 -15088 8856 -15007
rect 8823 -15171 8856 -15088
rect 9014 -15171 11218 -15007
rect 13216 -15027 13288 -14447
rect 15880 -14461 15934 -14402
rect 16010 -14367 16282 -14281
rect 16010 -14369 16214 -14367
rect 16010 -14405 16028 -14369
rect 16066 -14403 16214 -14369
rect 16252 -14403 16282 -14367
rect 16066 -14405 16282 -14403
rect 16010 -14441 16282 -14405
rect 16407 -14248 16581 -14227
rect 15377 -14521 15393 -14487
rect 15547 -14521 15563 -14487
rect 15879 -14529 15934 -14461
rect 16407 -14510 16428 -14248
rect 16565 -14510 16581 -14248
rect 16407 -14526 16581 -14510
rect 13216 -15033 13888 -15027
rect 15878 -15033 15934 -14529
rect 8823 -15179 11218 -15171
rect 8824 -15187 11218 -15179
rect 8830 -15189 11218 -15187
rect 9038 -15201 11218 -15189
rect 11528 -15057 13888 -15033
rect 11528 -15191 11562 -15057
rect 11680 -15191 13888 -15057
rect 9226 -15315 9242 -15281
rect 9276 -15315 9292 -15281
rect 9484 -15315 9500 -15281
rect 9534 -15315 9550 -15281
rect 9742 -15315 9758 -15281
rect 9792 -15315 9808 -15281
rect 10000 -15315 10016 -15281
rect 10050 -15315 10066 -15281
rect 10258 -15315 10274 -15281
rect 10308 -15315 10324 -15281
rect 10516 -15315 10532 -15281
rect 10566 -15315 10582 -15281
rect 10774 -15315 10790 -15281
rect 10824 -15315 10840 -15281
rect 11032 -15315 11048 -15281
rect 11082 -15315 11098 -15281
rect 9107 -15365 9152 -15347
rect 9107 -15401 9113 -15365
rect 9147 -15401 9152 -15365
rect 9107 -15435 9152 -15401
rect 9107 -15471 9113 -15435
rect 9147 -15471 9152 -15435
rect 9107 -15505 9152 -15471
rect 9107 -15541 9113 -15505
rect 9147 -15541 9152 -15505
rect 9107 -15783 9152 -15541
rect 9365 -15365 9410 -15321
rect 9365 -15401 9371 -15365
rect 9405 -15401 9410 -15365
rect 9365 -15435 9410 -15401
rect 9365 -15471 9371 -15435
rect 9405 -15471 9410 -15435
rect 9365 -15505 9410 -15471
rect 9365 -15541 9371 -15505
rect 9405 -15541 9410 -15505
rect 9226 -15625 9242 -15591
rect 9276 -15625 9292 -15591
rect 9226 -15733 9242 -15699
rect 9276 -15733 9292 -15699
rect 9107 -15819 9113 -15783
rect 9147 -15819 9152 -15783
rect 9107 -15853 9152 -15819
rect 9107 -15889 9113 -15853
rect 9147 -15889 9152 -15853
rect 9107 -15923 9152 -15889
rect 9107 -15959 9113 -15923
rect 9147 -15959 9152 -15923
rect 9107 -16201 9152 -15959
rect 9365 -15783 9410 -15541
rect 9622 -15365 9667 -15321
rect 9622 -15401 9629 -15365
rect 9663 -15401 9667 -15365
rect 9622 -15435 9667 -15401
rect 9622 -15471 9629 -15435
rect 9663 -15471 9667 -15435
rect 9622 -15506 9667 -15471
rect 9622 -15542 9629 -15506
rect 9663 -15542 9667 -15506
rect 9484 -15625 9500 -15591
rect 9534 -15625 9550 -15591
rect 9484 -15733 9500 -15699
rect 9534 -15733 9550 -15699
rect 9365 -15819 9371 -15783
rect 9405 -15819 9410 -15783
rect 9365 -15853 9410 -15819
rect 9365 -15889 9371 -15853
rect 9405 -15889 9410 -15853
rect 9365 -15923 9410 -15889
rect 9365 -15959 9371 -15923
rect 9405 -15959 9410 -15923
rect 9226 -16043 9242 -16009
rect 9276 -16043 9292 -16009
rect 9226 -16151 9242 -16117
rect 9276 -16151 9292 -16117
rect 9107 -16237 9113 -16201
rect 9147 -16237 9152 -16201
rect 9107 -16271 9152 -16237
rect 9107 -16307 9113 -16271
rect 9147 -16307 9152 -16271
rect 9107 -16341 9152 -16307
rect 9107 -16377 9113 -16341
rect 9147 -16377 9152 -16341
rect 9107 -16619 9152 -16377
rect 9365 -16201 9410 -15959
rect 9622 -15783 9667 -15542
rect 9882 -15365 9927 -15321
rect 9882 -15401 9887 -15365
rect 9921 -15401 9927 -15365
rect 9882 -15435 9927 -15401
rect 9882 -15471 9887 -15435
rect 9921 -15471 9927 -15435
rect 9882 -15505 9927 -15471
rect 9882 -15541 9887 -15505
rect 9921 -15541 9927 -15505
rect 9742 -15625 9758 -15591
rect 9792 -15625 9808 -15591
rect 9742 -15733 9758 -15699
rect 9792 -15733 9808 -15699
rect 9622 -15819 9629 -15783
rect 9663 -15819 9667 -15783
rect 9622 -15853 9667 -15819
rect 9622 -15889 9629 -15853
rect 9663 -15889 9667 -15853
rect 9622 -15924 9667 -15889
rect 9622 -15960 9629 -15924
rect 9663 -15960 9667 -15924
rect 9484 -16043 9500 -16009
rect 9534 -16043 9550 -16009
rect 9484 -16151 9500 -16117
rect 9534 -16151 9550 -16117
rect 9365 -16237 9371 -16201
rect 9405 -16237 9410 -16201
rect 9365 -16271 9410 -16237
rect 9365 -16307 9371 -16271
rect 9405 -16307 9410 -16271
rect 9365 -16341 9410 -16307
rect 9365 -16377 9371 -16341
rect 9405 -16377 9410 -16341
rect 9226 -16461 9242 -16427
rect 9276 -16461 9292 -16427
rect 9226 -16569 9242 -16535
rect 9276 -16569 9292 -16535
rect 9107 -16655 9113 -16619
rect 9147 -16655 9152 -16619
rect 9107 -16689 9152 -16655
rect 9107 -16725 9113 -16689
rect 9147 -16725 9152 -16689
rect 9107 -16759 9152 -16725
rect 9107 -16795 9113 -16759
rect 9147 -16795 9152 -16759
rect 9107 -17037 9152 -16795
rect 9365 -16619 9410 -16377
rect 9622 -16201 9667 -15960
rect 9882 -15783 9927 -15541
rect 10140 -15365 10185 -15321
rect 10140 -15401 10145 -15365
rect 10179 -15401 10185 -15365
rect 10140 -15435 10185 -15401
rect 10140 -15471 10145 -15435
rect 10179 -15471 10185 -15435
rect 10140 -15505 10185 -15471
rect 10140 -15541 10145 -15505
rect 10179 -15541 10185 -15505
rect 10000 -15625 10016 -15591
rect 10050 -15625 10066 -15591
rect 10000 -15733 10016 -15699
rect 10050 -15733 10066 -15699
rect 9882 -15819 9887 -15783
rect 9921 -15819 9927 -15783
rect 9882 -15853 9927 -15819
rect 9882 -15889 9887 -15853
rect 9921 -15889 9927 -15853
rect 9882 -15923 9927 -15889
rect 9882 -15959 9887 -15923
rect 9921 -15959 9927 -15923
rect 9742 -16043 9758 -16009
rect 9792 -16043 9808 -16009
rect 9742 -16151 9758 -16117
rect 9792 -16151 9808 -16117
rect 9622 -16237 9629 -16201
rect 9663 -16237 9667 -16201
rect 9622 -16271 9667 -16237
rect 9622 -16307 9629 -16271
rect 9663 -16307 9667 -16271
rect 9622 -16342 9667 -16307
rect 9622 -16378 9629 -16342
rect 9663 -16378 9667 -16342
rect 9484 -16461 9500 -16427
rect 9534 -16461 9550 -16427
rect 9484 -16569 9500 -16535
rect 9534 -16569 9550 -16535
rect 9365 -16655 9371 -16619
rect 9405 -16655 9410 -16619
rect 9365 -16689 9410 -16655
rect 9365 -16725 9371 -16689
rect 9405 -16725 9410 -16689
rect 9365 -16759 9410 -16725
rect 9365 -16795 9371 -16759
rect 9405 -16795 9410 -16759
rect 9226 -16879 9242 -16845
rect 9276 -16879 9292 -16845
rect 9226 -16987 9242 -16953
rect 9276 -16987 9292 -16953
rect 9107 -17073 9113 -17037
rect 9147 -17073 9152 -17037
rect 9107 -17107 9152 -17073
rect 9107 -17143 9113 -17107
rect 9147 -17143 9152 -17107
rect 9107 -17177 9152 -17143
rect 9107 -17213 9113 -17177
rect 9147 -17213 9152 -17177
rect 9107 -17455 9152 -17213
rect 9365 -17037 9410 -16795
rect 9622 -16619 9667 -16378
rect 9882 -16201 9927 -15959
rect 10140 -15783 10185 -15541
rect 10397 -15365 10442 -15321
rect 10397 -15401 10403 -15365
rect 10437 -15401 10442 -15365
rect 10397 -15435 10442 -15401
rect 10397 -15471 10403 -15435
rect 10437 -15471 10442 -15435
rect 10397 -15505 10442 -15471
rect 10397 -15541 10403 -15505
rect 10437 -15541 10442 -15505
rect 10258 -15625 10274 -15591
rect 10308 -15625 10324 -15591
rect 10258 -15733 10274 -15699
rect 10308 -15733 10324 -15699
rect 10140 -15819 10145 -15783
rect 10179 -15819 10185 -15783
rect 10140 -15853 10185 -15819
rect 10140 -15889 10145 -15853
rect 10179 -15889 10185 -15853
rect 10140 -15923 10185 -15889
rect 10140 -15959 10145 -15923
rect 10179 -15959 10185 -15923
rect 10000 -16043 10016 -16009
rect 10050 -16043 10066 -16009
rect 10000 -16151 10016 -16117
rect 10050 -16151 10066 -16117
rect 9882 -16237 9887 -16201
rect 9921 -16237 9927 -16201
rect 9882 -16271 9927 -16237
rect 9882 -16307 9887 -16271
rect 9921 -16307 9927 -16271
rect 9882 -16341 9927 -16307
rect 9882 -16377 9887 -16341
rect 9921 -16377 9927 -16341
rect 9742 -16461 9758 -16427
rect 9792 -16461 9808 -16427
rect 9742 -16569 9758 -16535
rect 9792 -16569 9808 -16535
rect 9622 -16655 9629 -16619
rect 9663 -16655 9667 -16619
rect 9622 -16689 9667 -16655
rect 9622 -16725 9629 -16689
rect 9663 -16725 9667 -16689
rect 9622 -16760 9667 -16725
rect 9622 -16796 9629 -16760
rect 9663 -16796 9667 -16760
rect 9484 -16879 9500 -16845
rect 9534 -16879 9550 -16845
rect 9484 -16987 9500 -16953
rect 9534 -16987 9550 -16953
rect 9365 -17073 9371 -17037
rect 9405 -17073 9410 -17037
rect 9365 -17107 9410 -17073
rect 9365 -17143 9371 -17107
rect 9405 -17143 9410 -17107
rect 9365 -17177 9410 -17143
rect 9365 -17213 9371 -17177
rect 9405 -17213 9410 -17177
rect 9226 -17297 9242 -17263
rect 9276 -17297 9292 -17263
rect 9226 -17405 9242 -17371
rect 9276 -17405 9292 -17371
rect 9107 -17491 9113 -17455
rect 9147 -17491 9152 -17455
rect 9107 -17525 9152 -17491
rect 9107 -17561 9113 -17525
rect 9147 -17561 9152 -17525
rect 9107 -17595 9152 -17561
rect 9107 -17631 9113 -17595
rect 9147 -17631 9152 -17595
rect 9107 -17873 9152 -17631
rect 9365 -17455 9410 -17213
rect 9622 -17037 9667 -16796
rect 9882 -16619 9927 -16377
rect 10140 -16201 10185 -15959
rect 10397 -15783 10442 -15541
rect 10654 -15365 10699 -15321
rect 10654 -15401 10661 -15365
rect 10695 -15401 10699 -15365
rect 10654 -15435 10699 -15401
rect 10654 -15471 10661 -15435
rect 10695 -15471 10699 -15435
rect 10654 -15505 10699 -15471
rect 10654 -15541 10661 -15505
rect 10695 -15541 10699 -15505
rect 10516 -15625 10532 -15591
rect 10566 -15625 10582 -15591
rect 10516 -15733 10532 -15699
rect 10566 -15733 10582 -15699
rect 10397 -15819 10403 -15783
rect 10437 -15819 10442 -15783
rect 10397 -15853 10442 -15819
rect 10397 -15889 10403 -15853
rect 10437 -15889 10442 -15853
rect 10397 -15923 10442 -15889
rect 10397 -15959 10403 -15923
rect 10437 -15959 10442 -15923
rect 10258 -16043 10274 -16009
rect 10308 -16043 10324 -16009
rect 10258 -16151 10274 -16117
rect 10308 -16151 10324 -16117
rect 10140 -16237 10145 -16201
rect 10179 -16237 10185 -16201
rect 10140 -16271 10185 -16237
rect 10140 -16307 10145 -16271
rect 10179 -16307 10185 -16271
rect 10140 -16341 10185 -16307
rect 10140 -16377 10145 -16341
rect 10179 -16377 10185 -16341
rect 10000 -16461 10016 -16427
rect 10050 -16461 10066 -16427
rect 10000 -16569 10016 -16535
rect 10050 -16569 10066 -16535
rect 9882 -16655 9887 -16619
rect 9921 -16655 9927 -16619
rect 9882 -16689 9927 -16655
rect 9882 -16725 9887 -16689
rect 9921 -16725 9927 -16689
rect 9882 -16759 9927 -16725
rect 9882 -16795 9887 -16759
rect 9921 -16795 9927 -16759
rect 9742 -16879 9758 -16845
rect 9792 -16879 9808 -16845
rect 9742 -16987 9758 -16953
rect 9792 -16987 9808 -16953
rect 9622 -17073 9629 -17037
rect 9663 -17073 9667 -17037
rect 9622 -17107 9667 -17073
rect 9622 -17143 9629 -17107
rect 9663 -17143 9667 -17107
rect 9622 -17178 9667 -17143
rect 9622 -17214 9629 -17178
rect 9663 -17214 9667 -17178
rect 9484 -17297 9500 -17263
rect 9534 -17297 9550 -17263
rect 9484 -17405 9500 -17371
rect 9534 -17405 9550 -17371
rect 9365 -17491 9371 -17455
rect 9405 -17491 9410 -17455
rect 9365 -17525 9410 -17491
rect 9365 -17561 9371 -17525
rect 9405 -17561 9410 -17525
rect 9365 -17595 9410 -17561
rect 9365 -17631 9371 -17595
rect 9405 -17631 9410 -17595
rect 9226 -17715 9242 -17681
rect 9276 -17715 9292 -17681
rect 9226 -17823 9242 -17789
rect 9276 -17823 9292 -17789
rect 9107 -17909 9113 -17873
rect 9147 -17909 9152 -17873
rect 9107 -17943 9152 -17909
rect 9107 -17979 9113 -17943
rect 9147 -17979 9152 -17943
rect 9107 -18013 9152 -17979
rect 9107 -18049 9113 -18013
rect 9147 -18049 9152 -18013
rect 9107 -18073 9152 -18049
rect 9106 -18275 9152 -18073
rect 9365 -17873 9410 -17631
rect 9622 -17455 9667 -17214
rect 9882 -17037 9927 -16795
rect 10140 -16619 10185 -16377
rect 10397 -16201 10442 -15959
rect 10654 -15783 10699 -15541
rect 10913 -15365 10958 -15321
rect 11170 -15357 11216 -15201
rect 11528 -15223 13888 -15191
rect 14134 -15067 16668 -15033
rect 14134 -15191 14168 -15067
rect 14280 -15191 16668 -15067
rect 14134 -15213 16668 -15191
rect 15878 -15219 16552 -15213
rect 11528 -15225 13886 -15223
rect 11896 -15315 11912 -15281
rect 11946 -15315 11962 -15281
rect 12154 -15315 12170 -15281
rect 12204 -15315 12220 -15281
rect 12412 -15315 12428 -15281
rect 12462 -15315 12478 -15281
rect 12670 -15315 12686 -15281
rect 12720 -15315 12736 -15281
rect 12928 -15315 12944 -15281
rect 12978 -15315 12994 -15281
rect 13186 -15315 13202 -15281
rect 13236 -15315 13252 -15281
rect 13444 -15315 13460 -15281
rect 13494 -15315 13510 -15281
rect 13702 -15315 13718 -15281
rect 13752 -15315 13768 -15281
rect 10913 -15401 10919 -15365
rect 10953 -15401 10958 -15365
rect 10913 -15435 10958 -15401
rect 10913 -15471 10919 -15435
rect 10953 -15471 10958 -15435
rect 10913 -15505 10958 -15471
rect 10913 -15541 10919 -15505
rect 10953 -15541 10958 -15505
rect 10774 -15625 10790 -15591
rect 10824 -15625 10840 -15591
rect 10774 -15733 10790 -15699
rect 10824 -15733 10840 -15699
rect 10654 -15819 10661 -15783
rect 10695 -15819 10699 -15783
rect 10654 -15853 10699 -15819
rect 10654 -15889 10661 -15853
rect 10695 -15889 10699 -15853
rect 10654 -15923 10699 -15889
rect 10654 -15959 10661 -15923
rect 10695 -15959 10699 -15923
rect 10516 -16043 10532 -16009
rect 10566 -16043 10582 -16009
rect 10516 -16151 10532 -16117
rect 10566 -16151 10582 -16117
rect 10397 -16237 10403 -16201
rect 10437 -16237 10442 -16201
rect 10397 -16271 10442 -16237
rect 10397 -16307 10403 -16271
rect 10437 -16307 10442 -16271
rect 10397 -16341 10442 -16307
rect 10397 -16377 10403 -16341
rect 10437 -16377 10442 -16341
rect 10258 -16461 10274 -16427
rect 10308 -16461 10324 -16427
rect 10258 -16569 10274 -16535
rect 10308 -16569 10324 -16535
rect 10140 -16655 10145 -16619
rect 10179 -16655 10185 -16619
rect 10140 -16689 10185 -16655
rect 10140 -16725 10145 -16689
rect 10179 -16725 10185 -16689
rect 10140 -16759 10185 -16725
rect 10140 -16795 10145 -16759
rect 10179 -16795 10185 -16759
rect 10000 -16879 10016 -16845
rect 10050 -16879 10066 -16845
rect 10000 -16987 10016 -16953
rect 10050 -16987 10066 -16953
rect 9882 -17073 9887 -17037
rect 9921 -17073 9927 -17037
rect 9882 -17107 9927 -17073
rect 9882 -17143 9887 -17107
rect 9921 -17143 9927 -17107
rect 9882 -17177 9927 -17143
rect 9882 -17213 9887 -17177
rect 9921 -17213 9927 -17177
rect 9742 -17297 9758 -17263
rect 9792 -17297 9808 -17263
rect 9742 -17405 9758 -17371
rect 9792 -17405 9808 -17371
rect 9622 -17491 9629 -17455
rect 9663 -17491 9667 -17455
rect 9622 -17525 9667 -17491
rect 9622 -17561 9629 -17525
rect 9663 -17561 9667 -17525
rect 9622 -17596 9667 -17561
rect 9622 -17632 9629 -17596
rect 9663 -17632 9667 -17596
rect 9484 -17715 9500 -17681
rect 9534 -17715 9550 -17681
rect 9484 -17823 9500 -17789
rect 9534 -17823 9550 -17789
rect 9365 -17909 9371 -17873
rect 9405 -17909 9410 -17873
rect 9365 -17943 9410 -17909
rect 9365 -17979 9371 -17943
rect 9405 -17979 9410 -17943
rect 9365 -18013 9410 -17979
rect 9365 -18049 9371 -18013
rect 9405 -18049 9410 -18013
rect 9226 -18133 9242 -18099
rect 9276 -18133 9292 -18099
rect 9365 -18167 9410 -18049
rect 9622 -17873 9667 -17632
rect 9882 -17455 9927 -17213
rect 10140 -17037 10185 -16795
rect 10397 -16619 10442 -16377
rect 10654 -16201 10699 -15959
rect 10913 -15783 10958 -15541
rect 11171 -15365 11216 -15357
rect 11171 -15401 11177 -15365
rect 11211 -15401 11216 -15365
rect 11171 -15435 11216 -15401
rect 11171 -15471 11177 -15435
rect 11211 -15471 11216 -15435
rect 11171 -15505 11216 -15471
rect 11171 -15541 11177 -15505
rect 11211 -15541 11216 -15505
rect 11032 -15625 11048 -15591
rect 11082 -15625 11098 -15591
rect 11032 -15733 11048 -15699
rect 11082 -15733 11098 -15699
rect 10913 -15819 10919 -15783
rect 10953 -15819 10958 -15783
rect 10913 -15853 10958 -15819
rect 10913 -15889 10919 -15853
rect 10953 -15889 10958 -15853
rect 10913 -15923 10958 -15889
rect 10913 -15959 10919 -15923
rect 10953 -15959 10958 -15923
rect 10774 -16043 10790 -16009
rect 10824 -16043 10840 -16009
rect 10774 -16151 10790 -16117
rect 10824 -16151 10840 -16117
rect 10654 -16237 10661 -16201
rect 10695 -16237 10699 -16201
rect 10654 -16271 10699 -16237
rect 10654 -16307 10661 -16271
rect 10695 -16307 10699 -16271
rect 10654 -16341 10699 -16307
rect 10654 -16377 10661 -16341
rect 10695 -16377 10699 -16341
rect 10516 -16461 10532 -16427
rect 10566 -16461 10582 -16427
rect 10516 -16569 10532 -16535
rect 10566 -16569 10582 -16535
rect 10397 -16655 10403 -16619
rect 10437 -16655 10442 -16619
rect 10397 -16689 10442 -16655
rect 10397 -16725 10403 -16689
rect 10437 -16725 10442 -16689
rect 10397 -16759 10442 -16725
rect 10397 -16795 10403 -16759
rect 10437 -16795 10442 -16759
rect 10258 -16879 10274 -16845
rect 10308 -16879 10324 -16845
rect 10258 -16987 10274 -16953
rect 10308 -16987 10324 -16953
rect 10140 -17073 10145 -17037
rect 10179 -17073 10185 -17037
rect 10140 -17107 10185 -17073
rect 10140 -17143 10145 -17107
rect 10179 -17143 10185 -17107
rect 10140 -17177 10185 -17143
rect 10140 -17213 10145 -17177
rect 10179 -17213 10185 -17177
rect 10000 -17297 10016 -17263
rect 10050 -17297 10066 -17263
rect 10000 -17405 10016 -17371
rect 10050 -17405 10066 -17371
rect 9882 -17491 9887 -17455
rect 9921 -17491 9927 -17455
rect 9882 -17525 9927 -17491
rect 9882 -17561 9887 -17525
rect 9921 -17561 9927 -17525
rect 9882 -17595 9927 -17561
rect 9882 -17631 9887 -17595
rect 9921 -17631 9927 -17595
rect 9742 -17715 9758 -17681
rect 9792 -17715 9808 -17681
rect 9742 -17823 9758 -17789
rect 9792 -17823 9808 -17789
rect 9622 -17909 9629 -17873
rect 9663 -17909 9667 -17873
rect 9622 -17943 9667 -17909
rect 9622 -17979 9629 -17943
rect 9663 -17979 9667 -17943
rect 9622 -18014 9667 -17979
rect 9622 -18050 9629 -18014
rect 9663 -18050 9667 -18014
rect 9484 -18133 9500 -18099
rect 9534 -18133 9550 -18099
rect 9622 -18167 9667 -18050
rect 9882 -17873 9927 -17631
rect 10140 -17455 10185 -17213
rect 10397 -17037 10442 -16795
rect 10654 -16619 10699 -16377
rect 10913 -16201 10958 -15959
rect 11171 -15783 11216 -15541
rect 11171 -15819 11177 -15783
rect 11211 -15819 11216 -15783
rect 11171 -15853 11216 -15819
rect 11171 -15889 11177 -15853
rect 11211 -15889 11216 -15853
rect 11171 -15923 11216 -15889
rect 11171 -15959 11177 -15923
rect 11211 -15959 11216 -15923
rect 11032 -16043 11048 -16009
rect 11082 -16043 11098 -16009
rect 11032 -16151 11048 -16117
rect 11082 -16151 11098 -16117
rect 10913 -16237 10919 -16201
rect 10953 -16237 10958 -16201
rect 10913 -16271 10958 -16237
rect 10913 -16307 10919 -16271
rect 10953 -16307 10958 -16271
rect 10913 -16341 10958 -16307
rect 10913 -16377 10919 -16341
rect 10953 -16377 10958 -16341
rect 10774 -16461 10790 -16427
rect 10824 -16461 10840 -16427
rect 10774 -16569 10790 -16535
rect 10824 -16569 10840 -16535
rect 10654 -16655 10661 -16619
rect 10695 -16655 10699 -16619
rect 10654 -16689 10699 -16655
rect 10654 -16725 10661 -16689
rect 10695 -16725 10699 -16689
rect 10654 -16759 10699 -16725
rect 10654 -16795 10661 -16759
rect 10695 -16795 10699 -16759
rect 10516 -16879 10532 -16845
rect 10566 -16879 10582 -16845
rect 10516 -16987 10532 -16953
rect 10566 -16987 10582 -16953
rect 10397 -17073 10403 -17037
rect 10437 -17073 10442 -17037
rect 10397 -17107 10442 -17073
rect 10397 -17143 10403 -17107
rect 10437 -17143 10442 -17107
rect 10397 -17177 10442 -17143
rect 10397 -17213 10403 -17177
rect 10437 -17213 10442 -17177
rect 10258 -17297 10274 -17263
rect 10308 -17297 10324 -17263
rect 10258 -17405 10274 -17371
rect 10308 -17405 10324 -17371
rect 10140 -17491 10145 -17455
rect 10179 -17491 10185 -17455
rect 10140 -17525 10185 -17491
rect 10140 -17561 10145 -17525
rect 10179 -17561 10185 -17525
rect 10140 -17595 10185 -17561
rect 10140 -17631 10145 -17595
rect 10179 -17631 10185 -17595
rect 10000 -17715 10016 -17681
rect 10050 -17715 10066 -17681
rect 10000 -17823 10016 -17789
rect 10050 -17823 10066 -17789
rect 9882 -17909 9887 -17873
rect 9921 -17909 9927 -17873
rect 9882 -17943 9927 -17909
rect 9882 -17979 9887 -17943
rect 9921 -17979 9927 -17943
rect 9882 -18013 9927 -17979
rect 9882 -18049 9887 -18013
rect 9921 -18049 9927 -18013
rect 9742 -18133 9758 -18099
rect 9792 -18133 9808 -18099
rect 9882 -18167 9927 -18049
rect 10140 -17873 10185 -17631
rect 10397 -17455 10442 -17213
rect 10654 -17037 10699 -16795
rect 10913 -16619 10958 -16377
rect 11171 -16201 11216 -15959
rect 11171 -16237 11177 -16201
rect 11211 -16237 11216 -16201
rect 11171 -16271 11216 -16237
rect 11171 -16307 11177 -16271
rect 11211 -16307 11216 -16271
rect 11171 -16341 11216 -16307
rect 11171 -16377 11177 -16341
rect 11211 -16377 11216 -16341
rect 11032 -16461 11048 -16427
rect 11082 -16461 11098 -16427
rect 11032 -16569 11048 -16535
rect 11082 -16569 11098 -16535
rect 10913 -16655 10919 -16619
rect 10953 -16655 10958 -16619
rect 10913 -16689 10958 -16655
rect 10913 -16725 10919 -16689
rect 10953 -16725 10958 -16689
rect 10913 -16759 10958 -16725
rect 10913 -16795 10919 -16759
rect 10953 -16795 10958 -16759
rect 10774 -16879 10790 -16845
rect 10824 -16879 10840 -16845
rect 10774 -16987 10790 -16953
rect 10824 -16987 10840 -16953
rect 10654 -17073 10661 -17037
rect 10695 -17073 10699 -17037
rect 10654 -17107 10699 -17073
rect 10654 -17143 10661 -17107
rect 10695 -17143 10699 -17107
rect 10654 -17177 10699 -17143
rect 10654 -17213 10661 -17177
rect 10695 -17213 10699 -17177
rect 10516 -17297 10532 -17263
rect 10566 -17297 10582 -17263
rect 10516 -17405 10532 -17371
rect 10566 -17405 10582 -17371
rect 10397 -17491 10403 -17455
rect 10437 -17491 10442 -17455
rect 10397 -17525 10442 -17491
rect 10397 -17561 10403 -17525
rect 10437 -17561 10442 -17525
rect 10397 -17595 10442 -17561
rect 10397 -17631 10403 -17595
rect 10437 -17631 10442 -17595
rect 10258 -17715 10274 -17681
rect 10308 -17715 10324 -17681
rect 10258 -17823 10274 -17789
rect 10308 -17823 10324 -17789
rect 10140 -17909 10145 -17873
rect 10179 -17909 10185 -17873
rect 10140 -17943 10185 -17909
rect 10140 -17979 10145 -17943
rect 10179 -17979 10185 -17943
rect 10140 -18013 10185 -17979
rect 10140 -18049 10145 -18013
rect 10179 -18049 10185 -18013
rect 10000 -18133 10016 -18099
rect 10050 -18133 10066 -18099
rect 10140 -18167 10185 -18049
rect 10397 -17873 10442 -17631
rect 10654 -17455 10699 -17213
rect 10913 -17037 10958 -16795
rect 11171 -16619 11216 -16377
rect 11171 -16655 11177 -16619
rect 11211 -16655 11216 -16619
rect 11171 -16689 11216 -16655
rect 11171 -16725 11177 -16689
rect 11211 -16725 11216 -16689
rect 11171 -16759 11216 -16725
rect 11171 -16795 11177 -16759
rect 11211 -16795 11216 -16759
rect 11032 -16879 11048 -16845
rect 11082 -16879 11098 -16845
rect 11032 -16987 11048 -16953
rect 11082 -16987 11098 -16953
rect 10913 -17073 10919 -17037
rect 10953 -17073 10958 -17037
rect 10913 -17107 10958 -17073
rect 10913 -17143 10919 -17107
rect 10953 -17143 10958 -17107
rect 10913 -17177 10958 -17143
rect 10913 -17213 10919 -17177
rect 10953 -17213 10958 -17177
rect 10774 -17297 10790 -17263
rect 10824 -17297 10840 -17263
rect 10774 -17405 10790 -17371
rect 10824 -17405 10840 -17371
rect 10654 -17491 10661 -17455
rect 10695 -17491 10699 -17455
rect 10654 -17525 10699 -17491
rect 10654 -17561 10661 -17525
rect 10695 -17561 10699 -17525
rect 10654 -17595 10699 -17561
rect 10654 -17631 10661 -17595
rect 10695 -17631 10699 -17595
rect 10516 -17715 10532 -17681
rect 10566 -17715 10582 -17681
rect 10516 -17823 10532 -17789
rect 10566 -17823 10582 -17789
rect 10397 -17909 10403 -17873
rect 10437 -17909 10442 -17873
rect 10397 -17943 10442 -17909
rect 10397 -17979 10403 -17943
rect 10437 -17979 10442 -17943
rect 10397 -18013 10442 -17979
rect 10397 -18049 10403 -18013
rect 10437 -18049 10442 -18013
rect 10258 -18133 10274 -18099
rect 10308 -18133 10324 -18099
rect 10397 -18167 10442 -18049
rect 10654 -17873 10699 -17631
rect 10913 -17455 10958 -17213
rect 11171 -17037 11216 -16795
rect 11171 -17073 11177 -17037
rect 11211 -17073 11216 -17037
rect 11171 -17107 11216 -17073
rect 11171 -17143 11177 -17107
rect 11211 -17143 11216 -17107
rect 11171 -17177 11216 -17143
rect 11171 -17213 11177 -17177
rect 11211 -17213 11216 -17177
rect 11032 -17297 11048 -17263
rect 11082 -17297 11098 -17263
rect 11032 -17405 11048 -17371
rect 11082 -17405 11098 -17371
rect 10913 -17491 10919 -17455
rect 10953 -17491 10958 -17455
rect 10913 -17525 10958 -17491
rect 10913 -17561 10919 -17525
rect 10953 -17561 10958 -17525
rect 10913 -17595 10958 -17561
rect 10913 -17631 10919 -17595
rect 10953 -17631 10958 -17595
rect 10774 -17715 10790 -17681
rect 10824 -17715 10840 -17681
rect 10774 -17823 10790 -17789
rect 10824 -17823 10840 -17789
rect 10654 -17909 10661 -17873
rect 10695 -17909 10699 -17873
rect 10654 -17943 10699 -17909
rect 10654 -17979 10661 -17943
rect 10695 -17979 10699 -17943
rect 10654 -18013 10699 -17979
rect 10654 -18049 10661 -18013
rect 10695 -18049 10699 -18013
rect 10516 -18133 10532 -18099
rect 10566 -18133 10582 -18099
rect 10654 -18167 10699 -18049
rect 10913 -17873 10958 -17631
rect 11171 -17455 11216 -17213
rect 11171 -17491 11177 -17455
rect 11211 -17491 11216 -17455
rect 11171 -17525 11216 -17491
rect 11171 -17561 11177 -17525
rect 11211 -17561 11216 -17525
rect 11171 -17595 11216 -17561
rect 11171 -17631 11177 -17595
rect 11211 -17631 11216 -17595
rect 11032 -17715 11048 -17681
rect 11082 -17715 11098 -17681
rect 11032 -17823 11048 -17789
rect 11082 -17823 11098 -17789
rect 10913 -17909 10919 -17873
rect 10953 -17909 10958 -17873
rect 10913 -17943 10958 -17909
rect 10913 -17979 10919 -17943
rect 10953 -17979 10958 -17943
rect 10913 -18013 10958 -17979
rect 10913 -18049 10919 -18013
rect 10953 -18049 10958 -18013
rect 10774 -18133 10790 -18099
rect 10824 -18133 10840 -18099
rect 10913 -18167 10958 -18049
rect 11171 -17873 11216 -17631
rect 11171 -17909 11177 -17873
rect 11211 -17909 11216 -17873
rect 11171 -17943 11216 -17909
rect 11171 -17979 11177 -17943
rect 11211 -17979 11216 -17943
rect 11171 -18013 11216 -17979
rect 11171 -18049 11177 -18013
rect 11211 -18049 11216 -18013
rect 11171 -18097 11216 -18049
rect 11777 -15365 11822 -15347
rect 11777 -15401 11783 -15365
rect 11817 -15401 11822 -15365
rect 11777 -15435 11822 -15401
rect 11777 -15471 11783 -15435
rect 11817 -15471 11822 -15435
rect 11777 -15505 11822 -15471
rect 11777 -15541 11783 -15505
rect 11817 -15541 11822 -15505
rect 11777 -15783 11822 -15541
rect 12035 -15365 12080 -15321
rect 12035 -15401 12041 -15365
rect 12075 -15401 12080 -15365
rect 12035 -15435 12080 -15401
rect 12035 -15471 12041 -15435
rect 12075 -15471 12080 -15435
rect 12035 -15505 12080 -15471
rect 12035 -15541 12041 -15505
rect 12075 -15541 12080 -15505
rect 11896 -15625 11912 -15591
rect 11946 -15625 11962 -15591
rect 11896 -15733 11912 -15699
rect 11946 -15733 11962 -15699
rect 11777 -15819 11783 -15783
rect 11817 -15819 11822 -15783
rect 11777 -15853 11822 -15819
rect 11777 -15889 11783 -15853
rect 11817 -15889 11822 -15853
rect 11777 -15923 11822 -15889
rect 11777 -15959 11783 -15923
rect 11817 -15959 11822 -15923
rect 11777 -16201 11822 -15959
rect 12035 -15783 12080 -15541
rect 12292 -15365 12337 -15321
rect 12292 -15401 12299 -15365
rect 12333 -15401 12337 -15365
rect 12292 -15435 12337 -15401
rect 12292 -15471 12299 -15435
rect 12333 -15471 12337 -15435
rect 12292 -15506 12337 -15471
rect 12292 -15542 12299 -15506
rect 12333 -15542 12337 -15506
rect 12154 -15625 12170 -15591
rect 12204 -15625 12220 -15591
rect 12154 -15733 12170 -15699
rect 12204 -15733 12220 -15699
rect 12035 -15819 12041 -15783
rect 12075 -15819 12080 -15783
rect 12035 -15853 12080 -15819
rect 12035 -15889 12041 -15853
rect 12075 -15889 12080 -15853
rect 12035 -15923 12080 -15889
rect 12035 -15959 12041 -15923
rect 12075 -15959 12080 -15923
rect 11896 -16043 11912 -16009
rect 11946 -16043 11962 -16009
rect 11896 -16151 11912 -16117
rect 11946 -16151 11962 -16117
rect 11777 -16237 11783 -16201
rect 11817 -16237 11822 -16201
rect 11777 -16271 11822 -16237
rect 11777 -16307 11783 -16271
rect 11817 -16307 11822 -16271
rect 11777 -16341 11822 -16307
rect 11777 -16377 11783 -16341
rect 11817 -16377 11822 -16341
rect 11777 -16619 11822 -16377
rect 12035 -16201 12080 -15959
rect 12292 -15783 12337 -15542
rect 12552 -15365 12597 -15321
rect 12552 -15401 12557 -15365
rect 12591 -15401 12597 -15365
rect 12552 -15435 12597 -15401
rect 12552 -15471 12557 -15435
rect 12591 -15471 12597 -15435
rect 12552 -15505 12597 -15471
rect 12552 -15541 12557 -15505
rect 12591 -15541 12597 -15505
rect 12412 -15625 12428 -15591
rect 12462 -15625 12478 -15591
rect 12412 -15733 12428 -15699
rect 12462 -15733 12478 -15699
rect 12292 -15819 12299 -15783
rect 12333 -15819 12337 -15783
rect 12292 -15853 12337 -15819
rect 12292 -15889 12299 -15853
rect 12333 -15889 12337 -15853
rect 12292 -15924 12337 -15889
rect 12292 -15960 12299 -15924
rect 12333 -15960 12337 -15924
rect 12154 -16043 12170 -16009
rect 12204 -16043 12220 -16009
rect 12154 -16151 12170 -16117
rect 12204 -16151 12220 -16117
rect 12035 -16237 12041 -16201
rect 12075 -16237 12080 -16201
rect 12035 -16271 12080 -16237
rect 12035 -16307 12041 -16271
rect 12075 -16307 12080 -16271
rect 12035 -16341 12080 -16307
rect 12035 -16377 12041 -16341
rect 12075 -16377 12080 -16341
rect 11896 -16461 11912 -16427
rect 11946 -16461 11962 -16427
rect 11896 -16569 11912 -16535
rect 11946 -16569 11962 -16535
rect 11777 -16655 11783 -16619
rect 11817 -16655 11822 -16619
rect 11777 -16689 11822 -16655
rect 11777 -16725 11783 -16689
rect 11817 -16725 11822 -16689
rect 11777 -16759 11822 -16725
rect 11777 -16795 11783 -16759
rect 11817 -16795 11822 -16759
rect 11777 -17037 11822 -16795
rect 12035 -16619 12080 -16377
rect 12292 -16201 12337 -15960
rect 12552 -15783 12597 -15541
rect 12810 -15365 12855 -15321
rect 12810 -15401 12815 -15365
rect 12849 -15401 12855 -15365
rect 12810 -15435 12855 -15401
rect 12810 -15471 12815 -15435
rect 12849 -15471 12855 -15435
rect 12810 -15505 12855 -15471
rect 12810 -15541 12815 -15505
rect 12849 -15541 12855 -15505
rect 12670 -15625 12686 -15591
rect 12720 -15625 12736 -15591
rect 12670 -15733 12686 -15699
rect 12720 -15733 12736 -15699
rect 12552 -15819 12557 -15783
rect 12591 -15819 12597 -15783
rect 12552 -15853 12597 -15819
rect 12552 -15889 12557 -15853
rect 12591 -15889 12597 -15853
rect 12552 -15923 12597 -15889
rect 12552 -15959 12557 -15923
rect 12591 -15959 12597 -15923
rect 12412 -16043 12428 -16009
rect 12462 -16043 12478 -16009
rect 12412 -16151 12428 -16117
rect 12462 -16151 12478 -16117
rect 12292 -16237 12299 -16201
rect 12333 -16237 12337 -16201
rect 12292 -16271 12337 -16237
rect 12292 -16307 12299 -16271
rect 12333 -16307 12337 -16271
rect 12292 -16342 12337 -16307
rect 12292 -16378 12299 -16342
rect 12333 -16378 12337 -16342
rect 12154 -16461 12170 -16427
rect 12204 -16461 12220 -16427
rect 12154 -16569 12170 -16535
rect 12204 -16569 12220 -16535
rect 12035 -16655 12041 -16619
rect 12075 -16655 12080 -16619
rect 12035 -16689 12080 -16655
rect 12035 -16725 12041 -16689
rect 12075 -16725 12080 -16689
rect 12035 -16759 12080 -16725
rect 12035 -16795 12041 -16759
rect 12075 -16795 12080 -16759
rect 11896 -16879 11912 -16845
rect 11946 -16879 11962 -16845
rect 11896 -16987 11912 -16953
rect 11946 -16987 11962 -16953
rect 11777 -17073 11783 -17037
rect 11817 -17073 11822 -17037
rect 11777 -17107 11822 -17073
rect 11777 -17143 11783 -17107
rect 11817 -17143 11822 -17107
rect 11777 -17177 11822 -17143
rect 11777 -17213 11783 -17177
rect 11817 -17213 11822 -17177
rect 11777 -17455 11822 -17213
rect 12035 -17037 12080 -16795
rect 12292 -16619 12337 -16378
rect 12552 -16201 12597 -15959
rect 12810 -15783 12855 -15541
rect 13067 -15365 13112 -15321
rect 13067 -15401 13073 -15365
rect 13107 -15401 13112 -15365
rect 13067 -15435 13112 -15401
rect 13067 -15471 13073 -15435
rect 13107 -15471 13112 -15435
rect 13067 -15505 13112 -15471
rect 13067 -15541 13073 -15505
rect 13107 -15541 13112 -15505
rect 12928 -15625 12944 -15591
rect 12978 -15625 12994 -15591
rect 12928 -15733 12944 -15699
rect 12978 -15733 12994 -15699
rect 12810 -15819 12815 -15783
rect 12849 -15819 12855 -15783
rect 12810 -15853 12855 -15819
rect 12810 -15889 12815 -15853
rect 12849 -15889 12855 -15853
rect 12810 -15923 12855 -15889
rect 12810 -15959 12815 -15923
rect 12849 -15959 12855 -15923
rect 12670 -16043 12686 -16009
rect 12720 -16043 12736 -16009
rect 12670 -16151 12686 -16117
rect 12720 -16151 12736 -16117
rect 12552 -16237 12557 -16201
rect 12591 -16237 12597 -16201
rect 12552 -16271 12597 -16237
rect 12552 -16307 12557 -16271
rect 12591 -16307 12597 -16271
rect 12552 -16341 12597 -16307
rect 12552 -16377 12557 -16341
rect 12591 -16377 12597 -16341
rect 12412 -16461 12428 -16427
rect 12462 -16461 12478 -16427
rect 12412 -16569 12428 -16535
rect 12462 -16569 12478 -16535
rect 12292 -16655 12299 -16619
rect 12333 -16655 12337 -16619
rect 12292 -16689 12337 -16655
rect 12292 -16725 12299 -16689
rect 12333 -16725 12337 -16689
rect 12292 -16760 12337 -16725
rect 12292 -16796 12299 -16760
rect 12333 -16796 12337 -16760
rect 12154 -16879 12170 -16845
rect 12204 -16879 12220 -16845
rect 12154 -16987 12170 -16953
rect 12204 -16987 12220 -16953
rect 12035 -17073 12041 -17037
rect 12075 -17073 12080 -17037
rect 12035 -17107 12080 -17073
rect 12035 -17143 12041 -17107
rect 12075 -17143 12080 -17107
rect 12035 -17177 12080 -17143
rect 12035 -17213 12041 -17177
rect 12075 -17213 12080 -17177
rect 11896 -17297 11912 -17263
rect 11946 -17297 11962 -17263
rect 11896 -17405 11912 -17371
rect 11946 -17405 11962 -17371
rect 11777 -17491 11783 -17455
rect 11817 -17491 11822 -17455
rect 11777 -17525 11822 -17491
rect 11777 -17561 11783 -17525
rect 11817 -17561 11822 -17525
rect 11777 -17595 11822 -17561
rect 11777 -17631 11783 -17595
rect 11817 -17631 11822 -17595
rect 11777 -17873 11822 -17631
rect 12035 -17455 12080 -17213
rect 12292 -17037 12337 -16796
rect 12552 -16619 12597 -16377
rect 12810 -16201 12855 -15959
rect 13067 -15783 13112 -15541
rect 13324 -15365 13369 -15321
rect 13324 -15401 13331 -15365
rect 13365 -15401 13369 -15365
rect 13324 -15435 13369 -15401
rect 13324 -15471 13331 -15435
rect 13365 -15471 13369 -15435
rect 13324 -15505 13369 -15471
rect 13324 -15541 13331 -15505
rect 13365 -15541 13369 -15505
rect 13186 -15625 13202 -15591
rect 13236 -15625 13252 -15591
rect 13186 -15733 13202 -15699
rect 13236 -15733 13252 -15699
rect 13067 -15819 13073 -15783
rect 13107 -15819 13112 -15783
rect 13067 -15853 13112 -15819
rect 13067 -15889 13073 -15853
rect 13107 -15889 13112 -15853
rect 13067 -15923 13112 -15889
rect 13067 -15959 13073 -15923
rect 13107 -15959 13112 -15923
rect 12928 -16043 12944 -16009
rect 12978 -16043 12994 -16009
rect 12928 -16151 12944 -16117
rect 12978 -16151 12994 -16117
rect 12810 -16237 12815 -16201
rect 12849 -16237 12855 -16201
rect 12810 -16271 12855 -16237
rect 12810 -16307 12815 -16271
rect 12849 -16307 12855 -16271
rect 12810 -16341 12855 -16307
rect 12810 -16377 12815 -16341
rect 12849 -16377 12855 -16341
rect 12670 -16461 12686 -16427
rect 12720 -16461 12736 -16427
rect 12670 -16569 12686 -16535
rect 12720 -16569 12736 -16535
rect 12552 -16655 12557 -16619
rect 12591 -16655 12597 -16619
rect 12552 -16689 12597 -16655
rect 12552 -16725 12557 -16689
rect 12591 -16725 12597 -16689
rect 12552 -16759 12597 -16725
rect 12552 -16795 12557 -16759
rect 12591 -16795 12597 -16759
rect 12412 -16879 12428 -16845
rect 12462 -16879 12478 -16845
rect 12412 -16987 12428 -16953
rect 12462 -16987 12478 -16953
rect 12292 -17073 12299 -17037
rect 12333 -17073 12337 -17037
rect 12292 -17107 12337 -17073
rect 12292 -17143 12299 -17107
rect 12333 -17143 12337 -17107
rect 12292 -17178 12337 -17143
rect 12292 -17214 12299 -17178
rect 12333 -17214 12337 -17178
rect 12154 -17297 12170 -17263
rect 12204 -17297 12220 -17263
rect 12154 -17405 12170 -17371
rect 12204 -17405 12220 -17371
rect 12035 -17491 12041 -17455
rect 12075 -17491 12080 -17455
rect 12035 -17525 12080 -17491
rect 12035 -17561 12041 -17525
rect 12075 -17561 12080 -17525
rect 12035 -17595 12080 -17561
rect 12035 -17631 12041 -17595
rect 12075 -17631 12080 -17595
rect 11896 -17715 11912 -17681
rect 11946 -17715 11962 -17681
rect 11896 -17823 11912 -17789
rect 11946 -17823 11962 -17789
rect 11777 -17909 11783 -17873
rect 11817 -17909 11822 -17873
rect 11777 -17943 11822 -17909
rect 11777 -17979 11783 -17943
rect 11817 -17979 11822 -17943
rect 11777 -18013 11822 -17979
rect 11777 -18049 11783 -18013
rect 11817 -18049 11822 -18013
rect 11032 -18133 11048 -18099
rect 11082 -18133 11098 -18099
rect 11777 -18117 11822 -18049
rect 12035 -17873 12080 -17631
rect 12292 -17455 12337 -17214
rect 12552 -17037 12597 -16795
rect 12810 -16619 12855 -16377
rect 13067 -16201 13112 -15959
rect 13324 -15783 13369 -15541
rect 13583 -15365 13628 -15321
rect 13842 -15345 13886 -15225
rect 14559 -15314 14575 -15280
rect 14609 -15314 14625 -15280
rect 14817 -15314 14833 -15280
rect 14867 -15314 14883 -15280
rect 15075 -15314 15091 -15280
rect 15125 -15314 15141 -15280
rect 15333 -15314 15349 -15280
rect 15383 -15314 15399 -15280
rect 15591 -15314 15607 -15280
rect 15641 -15314 15657 -15280
rect 15849 -15314 15865 -15280
rect 15899 -15314 15915 -15280
rect 16107 -15314 16123 -15280
rect 16157 -15314 16173 -15280
rect 16365 -15314 16381 -15280
rect 16415 -15314 16431 -15280
rect 13583 -15401 13589 -15365
rect 13623 -15401 13628 -15365
rect 13583 -15435 13628 -15401
rect 13583 -15471 13589 -15435
rect 13623 -15471 13628 -15435
rect 13583 -15505 13628 -15471
rect 13583 -15541 13589 -15505
rect 13623 -15541 13628 -15505
rect 13444 -15625 13460 -15591
rect 13494 -15625 13510 -15591
rect 13444 -15733 13460 -15699
rect 13494 -15733 13510 -15699
rect 13324 -15819 13331 -15783
rect 13365 -15819 13369 -15783
rect 13324 -15853 13369 -15819
rect 13324 -15889 13331 -15853
rect 13365 -15889 13369 -15853
rect 13324 -15923 13369 -15889
rect 13324 -15959 13331 -15923
rect 13365 -15959 13369 -15923
rect 13186 -16043 13202 -16009
rect 13236 -16043 13252 -16009
rect 13186 -16151 13202 -16117
rect 13236 -16151 13252 -16117
rect 13067 -16237 13073 -16201
rect 13107 -16237 13112 -16201
rect 13067 -16271 13112 -16237
rect 13067 -16307 13073 -16271
rect 13107 -16307 13112 -16271
rect 13067 -16341 13112 -16307
rect 13067 -16377 13073 -16341
rect 13107 -16377 13112 -16341
rect 12928 -16461 12944 -16427
rect 12978 -16461 12994 -16427
rect 12928 -16569 12944 -16535
rect 12978 -16569 12994 -16535
rect 12810 -16655 12815 -16619
rect 12849 -16655 12855 -16619
rect 12810 -16689 12855 -16655
rect 12810 -16725 12815 -16689
rect 12849 -16725 12855 -16689
rect 12810 -16759 12855 -16725
rect 12810 -16795 12815 -16759
rect 12849 -16795 12855 -16759
rect 12670 -16879 12686 -16845
rect 12720 -16879 12736 -16845
rect 12670 -16987 12686 -16953
rect 12720 -16987 12736 -16953
rect 12552 -17073 12557 -17037
rect 12591 -17073 12597 -17037
rect 12552 -17107 12597 -17073
rect 12552 -17143 12557 -17107
rect 12591 -17143 12597 -17107
rect 12552 -17177 12597 -17143
rect 12552 -17213 12557 -17177
rect 12591 -17213 12597 -17177
rect 12412 -17297 12428 -17263
rect 12462 -17297 12478 -17263
rect 12412 -17405 12428 -17371
rect 12462 -17405 12478 -17371
rect 12292 -17491 12299 -17455
rect 12333 -17491 12337 -17455
rect 12292 -17525 12337 -17491
rect 12292 -17561 12299 -17525
rect 12333 -17561 12337 -17525
rect 12292 -17596 12337 -17561
rect 12292 -17632 12299 -17596
rect 12333 -17632 12337 -17596
rect 12154 -17715 12170 -17681
rect 12204 -17715 12220 -17681
rect 12154 -17823 12170 -17789
rect 12204 -17823 12220 -17789
rect 12035 -17909 12041 -17873
rect 12075 -17909 12080 -17873
rect 12035 -17943 12080 -17909
rect 12035 -17979 12041 -17943
rect 12075 -17979 12080 -17943
rect 12035 -18013 12080 -17979
rect 12035 -18049 12041 -18013
rect 12075 -18049 12080 -18013
rect 9106 -18357 10336 -18275
rect 11774 -18299 11822 -18117
rect 11896 -18133 11912 -18099
rect 11946 -18133 11962 -18099
rect 12035 -18167 12080 -18049
rect 12292 -17873 12337 -17632
rect 12552 -17455 12597 -17213
rect 12810 -17037 12855 -16795
rect 13067 -16619 13112 -16377
rect 13324 -16201 13369 -15959
rect 13583 -15783 13628 -15541
rect 13841 -15365 13886 -15345
rect 13841 -15401 13847 -15365
rect 13881 -15401 13886 -15365
rect 13841 -15435 13886 -15401
rect 13841 -15471 13847 -15435
rect 13881 -15471 13886 -15435
rect 13841 -15505 13886 -15471
rect 13841 -15541 13847 -15505
rect 13881 -15541 13886 -15505
rect 13702 -15625 13718 -15591
rect 13752 -15625 13768 -15591
rect 13702 -15733 13718 -15699
rect 13752 -15733 13768 -15699
rect 13583 -15819 13589 -15783
rect 13623 -15819 13628 -15783
rect 13583 -15853 13628 -15819
rect 13583 -15889 13589 -15853
rect 13623 -15889 13628 -15853
rect 13583 -15923 13628 -15889
rect 13583 -15959 13589 -15923
rect 13623 -15959 13628 -15923
rect 13444 -16043 13460 -16009
rect 13494 -16043 13510 -16009
rect 13444 -16151 13460 -16117
rect 13494 -16151 13510 -16117
rect 13324 -16237 13331 -16201
rect 13365 -16237 13369 -16201
rect 13324 -16271 13369 -16237
rect 13324 -16307 13331 -16271
rect 13365 -16307 13369 -16271
rect 13324 -16341 13369 -16307
rect 13324 -16377 13331 -16341
rect 13365 -16377 13369 -16341
rect 13186 -16461 13202 -16427
rect 13236 -16461 13252 -16427
rect 13186 -16569 13202 -16535
rect 13236 -16569 13252 -16535
rect 13067 -16655 13073 -16619
rect 13107 -16655 13112 -16619
rect 13067 -16689 13112 -16655
rect 13067 -16725 13073 -16689
rect 13107 -16725 13112 -16689
rect 13067 -16759 13112 -16725
rect 13067 -16795 13073 -16759
rect 13107 -16795 13112 -16759
rect 12928 -16879 12944 -16845
rect 12978 -16879 12994 -16845
rect 12928 -16987 12944 -16953
rect 12978 -16987 12994 -16953
rect 12810 -17073 12815 -17037
rect 12849 -17073 12855 -17037
rect 12810 -17107 12855 -17073
rect 12810 -17143 12815 -17107
rect 12849 -17143 12855 -17107
rect 12810 -17177 12855 -17143
rect 12810 -17213 12815 -17177
rect 12849 -17213 12855 -17177
rect 12670 -17297 12686 -17263
rect 12720 -17297 12736 -17263
rect 12670 -17405 12686 -17371
rect 12720 -17405 12736 -17371
rect 12552 -17491 12557 -17455
rect 12591 -17491 12597 -17455
rect 12552 -17525 12597 -17491
rect 12552 -17561 12557 -17525
rect 12591 -17561 12597 -17525
rect 12552 -17595 12597 -17561
rect 12552 -17631 12557 -17595
rect 12591 -17631 12597 -17595
rect 12412 -17715 12428 -17681
rect 12462 -17715 12478 -17681
rect 12412 -17823 12428 -17789
rect 12462 -17823 12478 -17789
rect 12292 -17909 12299 -17873
rect 12333 -17909 12337 -17873
rect 12292 -17943 12337 -17909
rect 12292 -17979 12299 -17943
rect 12333 -17979 12337 -17943
rect 12292 -18014 12337 -17979
rect 12292 -18050 12299 -18014
rect 12333 -18050 12337 -18014
rect 12154 -18133 12170 -18099
rect 12204 -18133 12220 -18099
rect 12292 -18167 12337 -18050
rect 12552 -17873 12597 -17631
rect 12810 -17455 12855 -17213
rect 13067 -17037 13112 -16795
rect 13324 -16619 13369 -16377
rect 13583 -16201 13628 -15959
rect 13841 -15783 13886 -15541
rect 13841 -15819 13847 -15783
rect 13881 -15819 13886 -15783
rect 13841 -15853 13886 -15819
rect 13841 -15889 13847 -15853
rect 13881 -15889 13886 -15853
rect 13841 -15923 13886 -15889
rect 13841 -15959 13847 -15923
rect 13881 -15959 13886 -15923
rect 13702 -16043 13718 -16009
rect 13752 -16043 13768 -16009
rect 13702 -16151 13718 -16117
rect 13752 -16151 13768 -16117
rect 13583 -16237 13589 -16201
rect 13623 -16237 13628 -16201
rect 13583 -16271 13628 -16237
rect 13583 -16307 13589 -16271
rect 13623 -16307 13628 -16271
rect 13583 -16341 13628 -16307
rect 13583 -16377 13589 -16341
rect 13623 -16377 13628 -16341
rect 13444 -16461 13460 -16427
rect 13494 -16461 13510 -16427
rect 13444 -16569 13460 -16535
rect 13494 -16569 13510 -16535
rect 13324 -16655 13331 -16619
rect 13365 -16655 13369 -16619
rect 13324 -16689 13369 -16655
rect 13324 -16725 13331 -16689
rect 13365 -16725 13369 -16689
rect 13324 -16759 13369 -16725
rect 13324 -16795 13331 -16759
rect 13365 -16795 13369 -16759
rect 13186 -16879 13202 -16845
rect 13236 -16879 13252 -16845
rect 13186 -16987 13202 -16953
rect 13236 -16987 13252 -16953
rect 13067 -17073 13073 -17037
rect 13107 -17073 13112 -17037
rect 13067 -17107 13112 -17073
rect 13067 -17143 13073 -17107
rect 13107 -17143 13112 -17107
rect 13067 -17177 13112 -17143
rect 13067 -17213 13073 -17177
rect 13107 -17213 13112 -17177
rect 12928 -17297 12944 -17263
rect 12978 -17297 12994 -17263
rect 12928 -17405 12944 -17371
rect 12978 -17405 12994 -17371
rect 12810 -17491 12815 -17455
rect 12849 -17491 12855 -17455
rect 12810 -17525 12855 -17491
rect 12810 -17561 12815 -17525
rect 12849 -17561 12855 -17525
rect 12810 -17595 12855 -17561
rect 12810 -17631 12815 -17595
rect 12849 -17631 12855 -17595
rect 12670 -17715 12686 -17681
rect 12720 -17715 12736 -17681
rect 12670 -17823 12686 -17789
rect 12720 -17823 12736 -17789
rect 12552 -17909 12557 -17873
rect 12591 -17909 12597 -17873
rect 12552 -17943 12597 -17909
rect 12552 -17979 12557 -17943
rect 12591 -17979 12597 -17943
rect 12552 -18013 12597 -17979
rect 12552 -18049 12557 -18013
rect 12591 -18049 12597 -18013
rect 12412 -18133 12428 -18099
rect 12462 -18133 12478 -18099
rect 12552 -18167 12597 -18049
rect 12810 -17873 12855 -17631
rect 13067 -17455 13112 -17213
rect 13324 -17037 13369 -16795
rect 13583 -16619 13628 -16377
rect 13841 -16201 13886 -15959
rect 13841 -16237 13847 -16201
rect 13881 -16237 13886 -16201
rect 13841 -16271 13886 -16237
rect 13841 -16307 13847 -16271
rect 13881 -16307 13886 -16271
rect 13841 -16341 13886 -16307
rect 13841 -16377 13847 -16341
rect 13881 -16377 13886 -16341
rect 13702 -16461 13718 -16427
rect 13752 -16461 13768 -16427
rect 13702 -16569 13718 -16535
rect 13752 -16569 13768 -16535
rect 13583 -16655 13589 -16619
rect 13623 -16655 13628 -16619
rect 13583 -16689 13628 -16655
rect 13583 -16725 13589 -16689
rect 13623 -16725 13628 -16689
rect 13583 -16759 13628 -16725
rect 13583 -16795 13589 -16759
rect 13623 -16795 13628 -16759
rect 13444 -16879 13460 -16845
rect 13494 -16879 13510 -16845
rect 13444 -16987 13460 -16953
rect 13494 -16987 13510 -16953
rect 13324 -17073 13331 -17037
rect 13365 -17073 13369 -17037
rect 13324 -17107 13369 -17073
rect 13324 -17143 13331 -17107
rect 13365 -17143 13369 -17107
rect 13324 -17177 13369 -17143
rect 13324 -17213 13331 -17177
rect 13365 -17213 13369 -17177
rect 13186 -17297 13202 -17263
rect 13236 -17297 13252 -17263
rect 13186 -17405 13202 -17371
rect 13236 -17405 13252 -17371
rect 13067 -17491 13073 -17455
rect 13107 -17491 13112 -17455
rect 13067 -17525 13112 -17491
rect 13067 -17561 13073 -17525
rect 13107 -17561 13112 -17525
rect 13067 -17595 13112 -17561
rect 13067 -17631 13073 -17595
rect 13107 -17631 13112 -17595
rect 12928 -17715 12944 -17681
rect 12978 -17715 12994 -17681
rect 12928 -17823 12944 -17789
rect 12978 -17823 12994 -17789
rect 12810 -17909 12815 -17873
rect 12849 -17909 12855 -17873
rect 12810 -17943 12855 -17909
rect 12810 -17979 12815 -17943
rect 12849 -17979 12855 -17943
rect 12810 -18013 12855 -17979
rect 12810 -18049 12815 -18013
rect 12849 -18049 12855 -18013
rect 12670 -18133 12686 -18099
rect 12720 -18133 12736 -18099
rect 12810 -18167 12855 -18049
rect 13067 -17873 13112 -17631
rect 13324 -17455 13369 -17213
rect 13583 -17037 13628 -16795
rect 13841 -16619 13886 -16377
rect 13841 -16655 13847 -16619
rect 13881 -16655 13886 -16619
rect 13841 -16689 13886 -16655
rect 13841 -16725 13847 -16689
rect 13881 -16725 13886 -16689
rect 13841 -16759 13886 -16725
rect 13841 -16795 13847 -16759
rect 13881 -16795 13886 -16759
rect 13702 -16879 13718 -16845
rect 13752 -16879 13768 -16845
rect 13702 -16987 13718 -16953
rect 13752 -16987 13768 -16953
rect 13583 -17073 13589 -17037
rect 13623 -17073 13628 -17037
rect 13583 -17107 13628 -17073
rect 13583 -17143 13589 -17107
rect 13623 -17143 13628 -17107
rect 13583 -17177 13628 -17143
rect 13583 -17213 13589 -17177
rect 13623 -17213 13628 -17177
rect 13444 -17297 13460 -17263
rect 13494 -17297 13510 -17263
rect 13444 -17405 13460 -17371
rect 13494 -17405 13510 -17371
rect 13324 -17491 13331 -17455
rect 13365 -17491 13369 -17455
rect 13324 -17525 13369 -17491
rect 13324 -17561 13331 -17525
rect 13365 -17561 13369 -17525
rect 13324 -17595 13369 -17561
rect 13324 -17631 13331 -17595
rect 13365 -17631 13369 -17595
rect 13186 -17715 13202 -17681
rect 13236 -17715 13252 -17681
rect 13186 -17823 13202 -17789
rect 13236 -17823 13252 -17789
rect 13067 -17909 13073 -17873
rect 13107 -17909 13112 -17873
rect 13067 -17943 13112 -17909
rect 13067 -17979 13073 -17943
rect 13107 -17979 13112 -17943
rect 13067 -18013 13112 -17979
rect 13067 -18049 13073 -18013
rect 13107 -18049 13112 -18013
rect 12928 -18133 12944 -18099
rect 12978 -18133 12994 -18099
rect 13067 -18167 13112 -18049
rect 13324 -17873 13369 -17631
rect 13583 -17455 13628 -17213
rect 13841 -17037 13886 -16795
rect 13841 -17073 13847 -17037
rect 13881 -17073 13886 -17037
rect 13841 -17107 13886 -17073
rect 13841 -17143 13847 -17107
rect 13881 -17143 13886 -17107
rect 13841 -17177 13886 -17143
rect 13841 -17213 13847 -17177
rect 13881 -17213 13886 -17177
rect 13702 -17297 13718 -17263
rect 13752 -17297 13768 -17263
rect 13702 -17405 13718 -17371
rect 13752 -17405 13768 -17371
rect 13583 -17491 13589 -17455
rect 13623 -17491 13628 -17455
rect 13583 -17525 13628 -17491
rect 13583 -17561 13589 -17525
rect 13623 -17561 13628 -17525
rect 13583 -17595 13628 -17561
rect 13583 -17631 13589 -17595
rect 13623 -17631 13628 -17595
rect 13444 -17715 13460 -17681
rect 13494 -17715 13510 -17681
rect 13444 -17823 13460 -17789
rect 13494 -17823 13510 -17789
rect 13324 -17909 13331 -17873
rect 13365 -17909 13369 -17873
rect 13324 -17943 13369 -17909
rect 13324 -17979 13331 -17943
rect 13365 -17979 13369 -17943
rect 13324 -18013 13369 -17979
rect 13324 -18049 13331 -18013
rect 13365 -18049 13369 -18013
rect 13186 -18133 13202 -18099
rect 13236 -18133 13252 -18099
rect 13324 -18167 13369 -18049
rect 13583 -17873 13628 -17631
rect 13841 -17455 13886 -17213
rect 13841 -17491 13847 -17455
rect 13881 -17491 13886 -17455
rect 13841 -17525 13886 -17491
rect 13841 -17561 13847 -17525
rect 13881 -17561 13886 -17525
rect 13841 -17595 13886 -17561
rect 13841 -17631 13847 -17595
rect 13881 -17631 13886 -17595
rect 13702 -17715 13718 -17681
rect 13752 -17715 13768 -17681
rect 13702 -17823 13718 -17789
rect 13752 -17823 13768 -17789
rect 13583 -17909 13589 -17873
rect 13623 -17909 13628 -17873
rect 13583 -17943 13628 -17909
rect 13583 -17979 13589 -17943
rect 13623 -17979 13628 -17943
rect 13583 -18013 13628 -17979
rect 13583 -18049 13589 -18013
rect 13623 -18049 13628 -18013
rect 13444 -18133 13460 -18099
rect 13494 -18133 13510 -18099
rect 13583 -18167 13628 -18049
rect 13841 -17873 13886 -17631
rect 13841 -17909 13847 -17873
rect 13881 -17909 13886 -17873
rect 13841 -17943 13886 -17909
rect 13841 -17979 13847 -17943
rect 13881 -17979 13886 -17943
rect 13841 -18013 13886 -17979
rect 13841 -18049 13847 -18013
rect 13881 -18049 13886 -18013
rect 13841 -18079 13886 -18049
rect 14440 -15364 14485 -15347
rect 14440 -15400 14446 -15364
rect 14480 -15400 14485 -15364
rect 14440 -15434 14485 -15400
rect 14440 -15470 14446 -15434
rect 14480 -15470 14485 -15434
rect 14440 -15504 14485 -15470
rect 14440 -15540 14446 -15504
rect 14480 -15540 14485 -15504
rect 14440 -15782 14485 -15540
rect 14698 -15364 14743 -15320
rect 14698 -15400 14704 -15364
rect 14738 -15400 14743 -15364
rect 14698 -15434 14743 -15400
rect 14698 -15470 14704 -15434
rect 14738 -15470 14743 -15434
rect 14698 -15504 14743 -15470
rect 14698 -15540 14704 -15504
rect 14738 -15540 14743 -15504
rect 14559 -15624 14575 -15590
rect 14609 -15624 14625 -15590
rect 14559 -15732 14575 -15698
rect 14609 -15732 14625 -15698
rect 14440 -15818 14446 -15782
rect 14480 -15818 14485 -15782
rect 14440 -15852 14485 -15818
rect 14440 -15888 14446 -15852
rect 14480 -15888 14485 -15852
rect 14440 -15922 14485 -15888
rect 14440 -15958 14446 -15922
rect 14480 -15958 14485 -15922
rect 14440 -16200 14485 -15958
rect 14698 -15782 14743 -15540
rect 14955 -15364 15000 -15320
rect 14955 -15400 14962 -15364
rect 14996 -15400 15000 -15364
rect 14955 -15434 15000 -15400
rect 14955 -15470 14962 -15434
rect 14996 -15470 15000 -15434
rect 14955 -15505 15000 -15470
rect 14955 -15541 14962 -15505
rect 14996 -15541 15000 -15505
rect 14817 -15624 14833 -15590
rect 14867 -15624 14883 -15590
rect 14817 -15732 14833 -15698
rect 14867 -15732 14883 -15698
rect 14698 -15818 14704 -15782
rect 14738 -15818 14743 -15782
rect 14698 -15852 14743 -15818
rect 14698 -15888 14704 -15852
rect 14738 -15888 14743 -15852
rect 14698 -15922 14743 -15888
rect 14698 -15958 14704 -15922
rect 14738 -15958 14743 -15922
rect 14559 -16042 14575 -16008
rect 14609 -16042 14625 -16008
rect 14559 -16150 14575 -16116
rect 14609 -16150 14625 -16116
rect 14440 -16236 14446 -16200
rect 14480 -16236 14485 -16200
rect 14440 -16270 14485 -16236
rect 14440 -16306 14446 -16270
rect 14480 -16306 14485 -16270
rect 14440 -16340 14485 -16306
rect 14440 -16376 14446 -16340
rect 14480 -16376 14485 -16340
rect 14440 -16618 14485 -16376
rect 14698 -16200 14743 -15958
rect 14955 -15782 15000 -15541
rect 15215 -15364 15260 -15320
rect 15215 -15400 15220 -15364
rect 15254 -15400 15260 -15364
rect 15215 -15434 15260 -15400
rect 15215 -15470 15220 -15434
rect 15254 -15470 15260 -15434
rect 15215 -15504 15260 -15470
rect 15215 -15540 15220 -15504
rect 15254 -15540 15260 -15504
rect 15075 -15624 15091 -15590
rect 15125 -15624 15141 -15590
rect 15075 -15732 15091 -15698
rect 15125 -15732 15141 -15698
rect 14955 -15818 14962 -15782
rect 14996 -15818 15000 -15782
rect 14955 -15852 15000 -15818
rect 14955 -15888 14962 -15852
rect 14996 -15888 15000 -15852
rect 14955 -15923 15000 -15888
rect 14955 -15959 14962 -15923
rect 14996 -15959 15000 -15923
rect 14817 -16042 14833 -16008
rect 14867 -16042 14883 -16008
rect 14817 -16150 14833 -16116
rect 14867 -16150 14883 -16116
rect 14698 -16236 14704 -16200
rect 14738 -16236 14743 -16200
rect 14698 -16270 14743 -16236
rect 14698 -16306 14704 -16270
rect 14738 -16306 14743 -16270
rect 14698 -16340 14743 -16306
rect 14698 -16376 14704 -16340
rect 14738 -16376 14743 -16340
rect 14559 -16460 14575 -16426
rect 14609 -16460 14625 -16426
rect 14559 -16568 14575 -16534
rect 14609 -16568 14625 -16534
rect 14440 -16654 14446 -16618
rect 14480 -16654 14485 -16618
rect 14440 -16688 14485 -16654
rect 14440 -16724 14446 -16688
rect 14480 -16724 14485 -16688
rect 14440 -16758 14485 -16724
rect 14440 -16794 14446 -16758
rect 14480 -16794 14485 -16758
rect 14440 -17036 14485 -16794
rect 14698 -16618 14743 -16376
rect 14955 -16200 15000 -15959
rect 15215 -15782 15260 -15540
rect 15473 -15364 15518 -15320
rect 15473 -15400 15478 -15364
rect 15512 -15400 15518 -15364
rect 15473 -15434 15518 -15400
rect 15473 -15470 15478 -15434
rect 15512 -15470 15518 -15434
rect 15473 -15504 15518 -15470
rect 15473 -15540 15478 -15504
rect 15512 -15540 15518 -15504
rect 15333 -15624 15349 -15590
rect 15383 -15624 15399 -15590
rect 15333 -15732 15349 -15698
rect 15383 -15732 15399 -15698
rect 15215 -15818 15220 -15782
rect 15254 -15818 15260 -15782
rect 15215 -15852 15260 -15818
rect 15215 -15888 15220 -15852
rect 15254 -15888 15260 -15852
rect 15215 -15922 15260 -15888
rect 15215 -15958 15220 -15922
rect 15254 -15958 15260 -15922
rect 15075 -16042 15091 -16008
rect 15125 -16042 15141 -16008
rect 15075 -16150 15091 -16116
rect 15125 -16150 15141 -16116
rect 14955 -16236 14962 -16200
rect 14996 -16236 15000 -16200
rect 14955 -16270 15000 -16236
rect 14955 -16306 14962 -16270
rect 14996 -16306 15000 -16270
rect 14955 -16341 15000 -16306
rect 14955 -16377 14962 -16341
rect 14996 -16377 15000 -16341
rect 14817 -16460 14833 -16426
rect 14867 -16460 14883 -16426
rect 14817 -16568 14833 -16534
rect 14867 -16568 14883 -16534
rect 14698 -16654 14704 -16618
rect 14738 -16654 14743 -16618
rect 14698 -16688 14743 -16654
rect 14698 -16724 14704 -16688
rect 14738 -16724 14743 -16688
rect 14698 -16758 14743 -16724
rect 14698 -16794 14704 -16758
rect 14738 -16794 14743 -16758
rect 14559 -16878 14575 -16844
rect 14609 -16878 14625 -16844
rect 14559 -16986 14575 -16952
rect 14609 -16986 14625 -16952
rect 14440 -17072 14446 -17036
rect 14480 -17072 14485 -17036
rect 14440 -17106 14485 -17072
rect 14440 -17142 14446 -17106
rect 14480 -17142 14485 -17106
rect 14440 -17176 14485 -17142
rect 14440 -17212 14446 -17176
rect 14480 -17212 14485 -17176
rect 14440 -17454 14485 -17212
rect 14698 -17036 14743 -16794
rect 14955 -16618 15000 -16377
rect 15215 -16200 15260 -15958
rect 15473 -15782 15518 -15540
rect 15730 -15364 15775 -15320
rect 15730 -15400 15736 -15364
rect 15770 -15400 15775 -15364
rect 15730 -15434 15775 -15400
rect 15730 -15470 15736 -15434
rect 15770 -15470 15775 -15434
rect 15730 -15504 15775 -15470
rect 15730 -15540 15736 -15504
rect 15770 -15540 15775 -15504
rect 15591 -15624 15607 -15590
rect 15641 -15624 15657 -15590
rect 15591 -15732 15607 -15698
rect 15641 -15732 15657 -15698
rect 15473 -15818 15478 -15782
rect 15512 -15818 15518 -15782
rect 15473 -15852 15518 -15818
rect 15473 -15888 15478 -15852
rect 15512 -15888 15518 -15852
rect 15473 -15922 15518 -15888
rect 15473 -15958 15478 -15922
rect 15512 -15958 15518 -15922
rect 15333 -16042 15349 -16008
rect 15383 -16042 15399 -16008
rect 15333 -16150 15349 -16116
rect 15383 -16150 15399 -16116
rect 15215 -16236 15220 -16200
rect 15254 -16236 15260 -16200
rect 15215 -16270 15260 -16236
rect 15215 -16306 15220 -16270
rect 15254 -16306 15260 -16270
rect 15215 -16340 15260 -16306
rect 15215 -16376 15220 -16340
rect 15254 -16376 15260 -16340
rect 15075 -16460 15091 -16426
rect 15125 -16460 15141 -16426
rect 15075 -16568 15091 -16534
rect 15125 -16568 15141 -16534
rect 14955 -16654 14962 -16618
rect 14996 -16654 15000 -16618
rect 14955 -16688 15000 -16654
rect 14955 -16724 14962 -16688
rect 14996 -16724 15000 -16688
rect 14955 -16759 15000 -16724
rect 14955 -16795 14962 -16759
rect 14996 -16795 15000 -16759
rect 14817 -16878 14833 -16844
rect 14867 -16878 14883 -16844
rect 14817 -16986 14833 -16952
rect 14867 -16986 14883 -16952
rect 14698 -17072 14704 -17036
rect 14738 -17072 14743 -17036
rect 14698 -17106 14743 -17072
rect 14698 -17142 14704 -17106
rect 14738 -17142 14743 -17106
rect 14698 -17176 14743 -17142
rect 14698 -17212 14704 -17176
rect 14738 -17212 14743 -17176
rect 14559 -17296 14575 -17262
rect 14609 -17296 14625 -17262
rect 14559 -17404 14575 -17370
rect 14609 -17404 14625 -17370
rect 14440 -17490 14446 -17454
rect 14480 -17490 14485 -17454
rect 14440 -17524 14485 -17490
rect 14440 -17560 14446 -17524
rect 14480 -17560 14485 -17524
rect 14440 -17594 14485 -17560
rect 14440 -17630 14446 -17594
rect 14480 -17630 14485 -17594
rect 14440 -17872 14485 -17630
rect 14698 -17454 14743 -17212
rect 14955 -17036 15000 -16795
rect 15215 -16618 15260 -16376
rect 15473 -16200 15518 -15958
rect 15730 -15782 15775 -15540
rect 15987 -15364 16032 -15320
rect 15987 -15400 15994 -15364
rect 16028 -15400 16032 -15364
rect 15987 -15434 16032 -15400
rect 15987 -15470 15994 -15434
rect 16028 -15470 16032 -15434
rect 15987 -15504 16032 -15470
rect 15987 -15540 15994 -15504
rect 16028 -15540 16032 -15504
rect 15849 -15624 15865 -15590
rect 15899 -15624 15915 -15590
rect 15849 -15732 15865 -15698
rect 15899 -15732 15915 -15698
rect 15730 -15818 15736 -15782
rect 15770 -15818 15775 -15782
rect 15730 -15852 15775 -15818
rect 15730 -15888 15736 -15852
rect 15770 -15888 15775 -15852
rect 15730 -15922 15775 -15888
rect 15730 -15958 15736 -15922
rect 15770 -15958 15775 -15922
rect 15591 -16042 15607 -16008
rect 15641 -16042 15657 -16008
rect 15591 -16150 15607 -16116
rect 15641 -16150 15657 -16116
rect 15473 -16236 15478 -16200
rect 15512 -16236 15518 -16200
rect 15473 -16270 15518 -16236
rect 15473 -16306 15478 -16270
rect 15512 -16306 15518 -16270
rect 15473 -16340 15518 -16306
rect 15473 -16376 15478 -16340
rect 15512 -16376 15518 -16340
rect 15333 -16460 15349 -16426
rect 15383 -16460 15399 -16426
rect 15333 -16568 15349 -16534
rect 15383 -16568 15399 -16534
rect 15215 -16654 15220 -16618
rect 15254 -16654 15260 -16618
rect 15215 -16688 15260 -16654
rect 15215 -16724 15220 -16688
rect 15254 -16724 15260 -16688
rect 15215 -16758 15260 -16724
rect 15215 -16794 15220 -16758
rect 15254 -16794 15260 -16758
rect 15075 -16878 15091 -16844
rect 15125 -16878 15141 -16844
rect 15075 -16986 15091 -16952
rect 15125 -16986 15141 -16952
rect 14955 -17072 14962 -17036
rect 14996 -17072 15000 -17036
rect 14955 -17106 15000 -17072
rect 14955 -17142 14962 -17106
rect 14996 -17142 15000 -17106
rect 14955 -17177 15000 -17142
rect 14955 -17213 14962 -17177
rect 14996 -17213 15000 -17177
rect 14817 -17296 14833 -17262
rect 14867 -17296 14883 -17262
rect 14817 -17404 14833 -17370
rect 14867 -17404 14883 -17370
rect 14698 -17490 14704 -17454
rect 14738 -17490 14743 -17454
rect 14698 -17524 14743 -17490
rect 14698 -17560 14704 -17524
rect 14738 -17560 14743 -17524
rect 14698 -17594 14743 -17560
rect 14698 -17630 14704 -17594
rect 14738 -17630 14743 -17594
rect 14559 -17714 14575 -17680
rect 14609 -17714 14625 -17680
rect 14559 -17822 14575 -17788
rect 14609 -17822 14625 -17788
rect 14440 -17908 14446 -17872
rect 14480 -17908 14485 -17872
rect 14440 -17942 14485 -17908
rect 14440 -17978 14446 -17942
rect 14480 -17978 14485 -17942
rect 14440 -18012 14485 -17978
rect 14440 -18048 14446 -18012
rect 14480 -18048 14485 -18012
rect 13702 -18133 13718 -18099
rect 13752 -18133 13768 -18099
rect 14440 -18205 14485 -18048
rect 14698 -17872 14743 -17630
rect 14955 -17454 15000 -17213
rect 15215 -17036 15260 -16794
rect 15473 -16618 15518 -16376
rect 15730 -16200 15775 -15958
rect 15987 -15782 16032 -15540
rect 16246 -15364 16291 -15320
rect 16246 -15400 16252 -15364
rect 16286 -15400 16291 -15364
rect 16246 -15434 16291 -15400
rect 16246 -15470 16252 -15434
rect 16286 -15470 16291 -15434
rect 16246 -15504 16291 -15470
rect 16246 -15540 16252 -15504
rect 16286 -15540 16291 -15504
rect 16107 -15624 16123 -15590
rect 16157 -15624 16173 -15590
rect 16107 -15732 16123 -15698
rect 16157 -15732 16173 -15698
rect 15987 -15818 15994 -15782
rect 16028 -15818 16032 -15782
rect 15987 -15852 16032 -15818
rect 15987 -15888 15994 -15852
rect 16028 -15888 16032 -15852
rect 15987 -15922 16032 -15888
rect 15987 -15958 15994 -15922
rect 16028 -15958 16032 -15922
rect 15849 -16042 15865 -16008
rect 15899 -16042 15915 -16008
rect 15849 -16150 15865 -16116
rect 15899 -16150 15915 -16116
rect 15730 -16236 15736 -16200
rect 15770 -16236 15775 -16200
rect 15730 -16270 15775 -16236
rect 15730 -16306 15736 -16270
rect 15770 -16306 15775 -16270
rect 15730 -16340 15775 -16306
rect 15730 -16376 15736 -16340
rect 15770 -16376 15775 -16340
rect 15591 -16460 15607 -16426
rect 15641 -16460 15657 -16426
rect 15591 -16568 15607 -16534
rect 15641 -16568 15657 -16534
rect 15473 -16654 15478 -16618
rect 15512 -16654 15518 -16618
rect 15473 -16688 15518 -16654
rect 15473 -16724 15478 -16688
rect 15512 -16724 15518 -16688
rect 15473 -16758 15518 -16724
rect 15473 -16794 15478 -16758
rect 15512 -16794 15518 -16758
rect 15333 -16878 15349 -16844
rect 15383 -16878 15399 -16844
rect 15333 -16986 15349 -16952
rect 15383 -16986 15399 -16952
rect 15215 -17072 15220 -17036
rect 15254 -17072 15260 -17036
rect 15215 -17106 15260 -17072
rect 15215 -17142 15220 -17106
rect 15254 -17142 15260 -17106
rect 15215 -17176 15260 -17142
rect 15215 -17212 15220 -17176
rect 15254 -17212 15260 -17176
rect 15075 -17296 15091 -17262
rect 15125 -17296 15141 -17262
rect 15075 -17404 15091 -17370
rect 15125 -17404 15141 -17370
rect 14955 -17490 14962 -17454
rect 14996 -17490 15000 -17454
rect 14955 -17524 15000 -17490
rect 14955 -17560 14962 -17524
rect 14996 -17560 15000 -17524
rect 14955 -17595 15000 -17560
rect 14955 -17631 14962 -17595
rect 14996 -17631 15000 -17595
rect 14817 -17714 14833 -17680
rect 14867 -17714 14883 -17680
rect 14817 -17822 14833 -17788
rect 14867 -17822 14883 -17788
rect 14698 -17908 14704 -17872
rect 14738 -17908 14743 -17872
rect 14698 -17942 14743 -17908
rect 14698 -17978 14704 -17942
rect 14738 -17978 14743 -17942
rect 14698 -18012 14743 -17978
rect 14698 -18048 14704 -18012
rect 14738 -18048 14743 -18012
rect 14559 -18132 14575 -18098
rect 14609 -18132 14625 -18098
rect 14698 -18166 14743 -18048
rect 14955 -17872 15000 -17631
rect 15215 -17454 15260 -17212
rect 15473 -17036 15518 -16794
rect 15730 -16618 15775 -16376
rect 15987 -16200 16032 -15958
rect 16246 -15782 16291 -15540
rect 16504 -15349 16550 -15219
rect 16504 -15364 16549 -15349
rect 16504 -15400 16510 -15364
rect 16544 -15400 16549 -15364
rect 16504 -15434 16549 -15400
rect 16504 -15470 16510 -15434
rect 16544 -15470 16549 -15434
rect 16504 -15504 16549 -15470
rect 16504 -15540 16510 -15504
rect 16544 -15540 16549 -15504
rect 16365 -15624 16381 -15590
rect 16415 -15624 16431 -15590
rect 16365 -15732 16381 -15698
rect 16415 -15732 16431 -15698
rect 16246 -15818 16252 -15782
rect 16286 -15818 16291 -15782
rect 16246 -15852 16291 -15818
rect 16246 -15888 16252 -15852
rect 16286 -15888 16291 -15852
rect 16246 -15922 16291 -15888
rect 16246 -15958 16252 -15922
rect 16286 -15958 16291 -15922
rect 16107 -16042 16123 -16008
rect 16157 -16042 16173 -16008
rect 16107 -16150 16123 -16116
rect 16157 -16150 16173 -16116
rect 15987 -16236 15994 -16200
rect 16028 -16236 16032 -16200
rect 15987 -16270 16032 -16236
rect 15987 -16306 15994 -16270
rect 16028 -16306 16032 -16270
rect 15987 -16340 16032 -16306
rect 15987 -16376 15994 -16340
rect 16028 -16376 16032 -16340
rect 15849 -16460 15865 -16426
rect 15899 -16460 15915 -16426
rect 15849 -16568 15865 -16534
rect 15899 -16568 15915 -16534
rect 15730 -16654 15736 -16618
rect 15770 -16654 15775 -16618
rect 15730 -16688 15775 -16654
rect 15730 -16724 15736 -16688
rect 15770 -16724 15775 -16688
rect 15730 -16758 15775 -16724
rect 15730 -16794 15736 -16758
rect 15770 -16794 15775 -16758
rect 15591 -16878 15607 -16844
rect 15641 -16878 15657 -16844
rect 15591 -16986 15607 -16952
rect 15641 -16986 15657 -16952
rect 15473 -17072 15478 -17036
rect 15512 -17072 15518 -17036
rect 15473 -17106 15518 -17072
rect 15473 -17142 15478 -17106
rect 15512 -17142 15518 -17106
rect 15473 -17176 15518 -17142
rect 15473 -17212 15478 -17176
rect 15512 -17212 15518 -17176
rect 15333 -17296 15349 -17262
rect 15383 -17296 15399 -17262
rect 15333 -17404 15349 -17370
rect 15383 -17404 15399 -17370
rect 15215 -17490 15220 -17454
rect 15254 -17490 15260 -17454
rect 15215 -17524 15260 -17490
rect 15215 -17560 15220 -17524
rect 15254 -17560 15260 -17524
rect 15215 -17594 15260 -17560
rect 15215 -17630 15220 -17594
rect 15254 -17630 15260 -17594
rect 15075 -17714 15091 -17680
rect 15125 -17714 15141 -17680
rect 15075 -17822 15091 -17788
rect 15125 -17822 15141 -17788
rect 14955 -17908 14962 -17872
rect 14996 -17908 15000 -17872
rect 14955 -17942 15000 -17908
rect 14955 -17978 14962 -17942
rect 14996 -17978 15000 -17942
rect 14955 -18013 15000 -17978
rect 14955 -18049 14962 -18013
rect 14996 -18049 15000 -18013
rect 14817 -18132 14833 -18098
rect 14867 -18132 14883 -18098
rect 14955 -18166 15000 -18049
rect 15215 -17872 15260 -17630
rect 15473 -17454 15518 -17212
rect 15730 -17036 15775 -16794
rect 15987 -16618 16032 -16376
rect 16246 -16200 16291 -15958
rect 16504 -15782 16549 -15540
rect 16504 -15818 16510 -15782
rect 16544 -15818 16549 -15782
rect 16504 -15852 16549 -15818
rect 16504 -15888 16510 -15852
rect 16544 -15888 16549 -15852
rect 16504 -15922 16549 -15888
rect 16504 -15958 16510 -15922
rect 16544 -15958 16549 -15922
rect 16365 -16042 16381 -16008
rect 16415 -16042 16431 -16008
rect 16365 -16150 16381 -16116
rect 16415 -16150 16431 -16116
rect 16246 -16236 16252 -16200
rect 16286 -16236 16291 -16200
rect 16246 -16270 16291 -16236
rect 16246 -16306 16252 -16270
rect 16286 -16306 16291 -16270
rect 16246 -16340 16291 -16306
rect 16246 -16376 16252 -16340
rect 16286 -16376 16291 -16340
rect 16107 -16460 16123 -16426
rect 16157 -16460 16173 -16426
rect 16107 -16568 16123 -16534
rect 16157 -16568 16173 -16534
rect 15987 -16654 15994 -16618
rect 16028 -16654 16032 -16618
rect 15987 -16688 16032 -16654
rect 15987 -16724 15994 -16688
rect 16028 -16724 16032 -16688
rect 15987 -16758 16032 -16724
rect 15987 -16794 15994 -16758
rect 16028 -16794 16032 -16758
rect 15849 -16878 15865 -16844
rect 15899 -16878 15915 -16844
rect 15849 -16986 15865 -16952
rect 15899 -16986 15915 -16952
rect 15730 -17072 15736 -17036
rect 15770 -17072 15775 -17036
rect 15730 -17106 15775 -17072
rect 15730 -17142 15736 -17106
rect 15770 -17142 15775 -17106
rect 15730 -17176 15775 -17142
rect 15730 -17212 15736 -17176
rect 15770 -17212 15775 -17176
rect 15591 -17296 15607 -17262
rect 15641 -17296 15657 -17262
rect 15591 -17404 15607 -17370
rect 15641 -17404 15657 -17370
rect 15473 -17490 15478 -17454
rect 15512 -17490 15518 -17454
rect 15473 -17524 15518 -17490
rect 15473 -17560 15478 -17524
rect 15512 -17560 15518 -17524
rect 15473 -17594 15518 -17560
rect 15473 -17630 15478 -17594
rect 15512 -17630 15518 -17594
rect 15333 -17714 15349 -17680
rect 15383 -17714 15399 -17680
rect 15333 -17822 15349 -17788
rect 15383 -17822 15399 -17788
rect 15215 -17908 15220 -17872
rect 15254 -17908 15260 -17872
rect 15215 -17942 15260 -17908
rect 15215 -17978 15220 -17942
rect 15254 -17978 15260 -17942
rect 15215 -18012 15260 -17978
rect 15215 -18048 15220 -18012
rect 15254 -18048 15260 -18012
rect 15075 -18132 15091 -18098
rect 15125 -18132 15141 -18098
rect 15215 -18166 15260 -18048
rect 15473 -17872 15518 -17630
rect 15730 -17454 15775 -17212
rect 15987 -17036 16032 -16794
rect 16246 -16618 16291 -16376
rect 16504 -16200 16549 -15958
rect 16504 -16236 16510 -16200
rect 16544 -16236 16549 -16200
rect 16504 -16270 16549 -16236
rect 16504 -16306 16510 -16270
rect 16544 -16306 16549 -16270
rect 16504 -16340 16549 -16306
rect 16504 -16376 16510 -16340
rect 16544 -16376 16549 -16340
rect 16365 -16460 16381 -16426
rect 16415 -16460 16431 -16426
rect 16365 -16568 16381 -16534
rect 16415 -16568 16431 -16534
rect 16246 -16654 16252 -16618
rect 16286 -16654 16291 -16618
rect 16246 -16688 16291 -16654
rect 16246 -16724 16252 -16688
rect 16286 -16724 16291 -16688
rect 16246 -16758 16291 -16724
rect 16246 -16794 16252 -16758
rect 16286 -16794 16291 -16758
rect 16107 -16878 16123 -16844
rect 16157 -16878 16173 -16844
rect 16107 -16986 16123 -16952
rect 16157 -16986 16173 -16952
rect 15987 -17072 15994 -17036
rect 16028 -17072 16032 -17036
rect 15987 -17106 16032 -17072
rect 15987 -17142 15994 -17106
rect 16028 -17142 16032 -17106
rect 15987 -17176 16032 -17142
rect 15987 -17212 15994 -17176
rect 16028 -17212 16032 -17176
rect 15849 -17296 15865 -17262
rect 15899 -17296 15915 -17262
rect 15849 -17404 15865 -17370
rect 15899 -17404 15915 -17370
rect 15730 -17490 15736 -17454
rect 15770 -17490 15775 -17454
rect 15730 -17524 15775 -17490
rect 15730 -17560 15736 -17524
rect 15770 -17560 15775 -17524
rect 15730 -17594 15775 -17560
rect 15730 -17630 15736 -17594
rect 15770 -17630 15775 -17594
rect 15591 -17714 15607 -17680
rect 15641 -17714 15657 -17680
rect 15591 -17822 15607 -17788
rect 15641 -17822 15657 -17788
rect 15473 -17908 15478 -17872
rect 15512 -17908 15518 -17872
rect 15473 -17942 15518 -17908
rect 15473 -17978 15478 -17942
rect 15512 -17978 15518 -17942
rect 15473 -18012 15518 -17978
rect 15473 -18048 15478 -18012
rect 15512 -18048 15518 -18012
rect 15333 -18132 15349 -18098
rect 15383 -18132 15399 -18098
rect 15473 -18166 15518 -18048
rect 15730 -17872 15775 -17630
rect 15987 -17454 16032 -17212
rect 16246 -17036 16291 -16794
rect 16504 -16618 16549 -16376
rect 16504 -16654 16510 -16618
rect 16544 -16654 16549 -16618
rect 16504 -16688 16549 -16654
rect 16504 -16724 16510 -16688
rect 16544 -16724 16549 -16688
rect 16504 -16758 16549 -16724
rect 16504 -16794 16510 -16758
rect 16544 -16794 16549 -16758
rect 16365 -16878 16381 -16844
rect 16415 -16878 16431 -16844
rect 16365 -16986 16381 -16952
rect 16415 -16986 16431 -16952
rect 16246 -17072 16252 -17036
rect 16286 -17072 16291 -17036
rect 16246 -17106 16291 -17072
rect 16246 -17142 16252 -17106
rect 16286 -17142 16291 -17106
rect 16246 -17176 16291 -17142
rect 16246 -17212 16252 -17176
rect 16286 -17212 16291 -17176
rect 16107 -17296 16123 -17262
rect 16157 -17296 16173 -17262
rect 16107 -17404 16123 -17370
rect 16157 -17404 16173 -17370
rect 15987 -17490 15994 -17454
rect 16028 -17490 16032 -17454
rect 15987 -17524 16032 -17490
rect 15987 -17560 15994 -17524
rect 16028 -17560 16032 -17524
rect 15987 -17594 16032 -17560
rect 15987 -17630 15994 -17594
rect 16028 -17630 16032 -17594
rect 15849 -17714 15865 -17680
rect 15899 -17714 15915 -17680
rect 15849 -17822 15865 -17788
rect 15899 -17822 15915 -17788
rect 15730 -17908 15736 -17872
rect 15770 -17908 15775 -17872
rect 15730 -17942 15775 -17908
rect 15730 -17978 15736 -17942
rect 15770 -17978 15775 -17942
rect 15730 -18012 15775 -17978
rect 15730 -18048 15736 -18012
rect 15770 -18048 15775 -18012
rect 15591 -18132 15607 -18098
rect 15641 -18132 15657 -18098
rect 15730 -18166 15775 -18048
rect 15987 -17872 16032 -17630
rect 16246 -17454 16291 -17212
rect 16504 -17036 16549 -16794
rect 16504 -17072 16510 -17036
rect 16544 -17072 16549 -17036
rect 16504 -17106 16549 -17072
rect 16504 -17142 16510 -17106
rect 16544 -17142 16549 -17106
rect 16504 -17176 16549 -17142
rect 16504 -17212 16510 -17176
rect 16544 -17212 16549 -17176
rect 16365 -17296 16381 -17262
rect 16415 -17296 16431 -17262
rect 16365 -17404 16381 -17370
rect 16415 -17404 16431 -17370
rect 16246 -17490 16252 -17454
rect 16286 -17490 16291 -17454
rect 16246 -17524 16291 -17490
rect 16246 -17560 16252 -17524
rect 16286 -17560 16291 -17524
rect 16246 -17594 16291 -17560
rect 16246 -17630 16252 -17594
rect 16286 -17630 16291 -17594
rect 16107 -17714 16123 -17680
rect 16157 -17714 16173 -17680
rect 16107 -17822 16123 -17788
rect 16157 -17822 16173 -17788
rect 15987 -17908 15994 -17872
rect 16028 -17908 16032 -17872
rect 15987 -17942 16032 -17908
rect 15987 -17978 15994 -17942
rect 16028 -17978 16032 -17942
rect 15987 -18012 16032 -17978
rect 15987 -18048 15994 -18012
rect 16028 -18048 16032 -18012
rect 15849 -18132 15865 -18098
rect 15899 -18132 15915 -18098
rect 15987 -18166 16032 -18048
rect 16246 -17872 16291 -17630
rect 16504 -17454 16549 -17212
rect 16504 -17490 16510 -17454
rect 16544 -17490 16549 -17454
rect 16504 -17524 16549 -17490
rect 16504 -17560 16510 -17524
rect 16544 -17560 16549 -17524
rect 16504 -17594 16549 -17560
rect 16504 -17630 16510 -17594
rect 16544 -17630 16549 -17594
rect 16365 -17714 16381 -17680
rect 16415 -17714 16431 -17680
rect 16365 -17822 16381 -17788
rect 16415 -17822 16431 -17788
rect 16246 -17908 16252 -17872
rect 16286 -17908 16291 -17872
rect 16246 -17942 16291 -17908
rect 16246 -17978 16252 -17942
rect 16286 -17978 16291 -17942
rect 16246 -18012 16291 -17978
rect 16246 -18048 16252 -18012
rect 16286 -18048 16291 -18012
rect 16107 -18132 16123 -18098
rect 16157 -18132 16173 -18098
rect 16246 -18166 16291 -18048
rect 16504 -17872 16549 -17630
rect 16504 -17908 16510 -17872
rect 16544 -17908 16549 -17872
rect 16504 -17942 16549 -17908
rect 16504 -17978 16510 -17942
rect 16544 -17978 16549 -17942
rect 16504 -18012 16549 -17978
rect 16504 -18048 16510 -18012
rect 16544 -18048 16549 -18012
rect 16987 -18029 17137 -14165
rect 16504 -18069 16549 -18048
rect 16365 -18132 16381 -18098
rect 16415 -18132 16431 -18098
rect 14434 -18289 14486 -18205
rect 14434 -18290 15664 -18289
rect 10264 -18417 10334 -18357
rect 11774 -18387 13002 -18299
rect 14434 -18351 15666 -18290
rect 11774 -18395 13003 -18387
rect 9106 -18475 9122 -18441
rect 9156 -18475 9172 -18441
rect 9646 -18475 9662 -18441
rect 9696 -18475 9712 -18441
rect 10126 -18475 10137 -18441
rect 10187 -18475 10192 -18441
rect 8967 -18527 9029 -18505
rect 8967 -18561 8993 -18527
rect 9027 -18561 9029 -18527
rect 8967 -18595 9029 -18561
rect 8967 -18631 8993 -18595
rect 9027 -18631 9029 -18595
rect 8967 -18665 9029 -18631
rect 8967 -18699 8993 -18665
rect 9027 -18699 9029 -18665
rect 8967 -18741 9029 -18699
rect 9245 -18527 9313 -18507
rect 9245 -18561 9251 -18527
rect 9285 -18561 9313 -18527
rect 9245 -18595 9313 -18561
rect 9245 -18631 9251 -18595
rect 9285 -18631 9313 -18595
rect 9245 -18665 9313 -18631
rect 9245 -18699 9251 -18665
rect 9285 -18699 9313 -18665
rect 9245 -18743 9313 -18699
rect 9507 -18527 9569 -18505
rect 9507 -18561 9533 -18527
rect 9567 -18561 9569 -18527
rect 9507 -18595 9569 -18561
rect 9507 -18631 9533 -18595
rect 9567 -18631 9569 -18595
rect 9507 -18665 9569 -18631
rect 9507 -18699 9533 -18665
rect 9567 -18699 9569 -18665
rect 9507 -18741 9569 -18699
rect 9785 -18527 9853 -18507
rect 9785 -18561 9791 -18527
rect 9825 -18561 9853 -18527
rect 9785 -18595 9853 -18561
rect 9785 -18631 9791 -18595
rect 9825 -18631 9853 -18595
rect 9785 -18665 9853 -18631
rect 9785 -18699 9791 -18665
rect 9825 -18699 9853 -18665
rect 9785 -18743 9853 -18699
rect 9987 -18527 10049 -18505
rect 9987 -18561 10013 -18527
rect 10047 -18561 10049 -18527
rect 9987 -18595 10049 -18561
rect 9987 -18631 10013 -18595
rect 10047 -18631 10049 -18595
rect 9987 -18665 10049 -18631
rect 9987 -18699 10013 -18665
rect 10047 -18699 10049 -18665
rect 9106 -18785 9122 -18751
rect 9156 -18785 9172 -18751
rect 9646 -18785 9662 -18751
rect 9696 -18785 9712 -18751
rect 9987 -18870 10049 -18699
rect 10265 -18527 10333 -18417
rect 10629 -18473 10645 -18439
rect 10679 -18473 10695 -18439
rect 11139 -18463 11155 -18429
rect 11189 -18463 11205 -18429
rect 11776 -18475 11792 -18441
rect 11826 -18475 11842 -18441
rect 12316 -18475 12332 -18441
rect 12366 -18475 12382 -18441
rect 12796 -18475 12807 -18441
rect 12857 -18475 12862 -18441
rect 10265 -18561 10271 -18527
rect 10305 -18561 10333 -18527
rect 10265 -18595 10333 -18561
rect 10265 -18631 10271 -18595
rect 10305 -18631 10333 -18595
rect 10265 -18665 10333 -18631
rect 10265 -18699 10271 -18665
rect 10305 -18699 10333 -18665
rect 10265 -18743 10333 -18699
rect 10490 -18525 10552 -18503
rect 10490 -18559 10516 -18525
rect 10550 -18559 10552 -18525
rect 10490 -18593 10552 -18559
rect 10490 -18629 10516 -18593
rect 10550 -18629 10552 -18593
rect 10490 -18663 10552 -18629
rect 10490 -18697 10516 -18663
rect 10550 -18697 10552 -18663
rect 10490 -18739 10552 -18697
rect 10768 -18525 10836 -18505
rect 10768 -18559 10774 -18525
rect 10808 -18559 10836 -18525
rect 10768 -18593 10836 -18559
rect 10768 -18629 10774 -18593
rect 10808 -18629 10836 -18593
rect 10768 -18663 10836 -18629
rect 10768 -18697 10774 -18663
rect 10808 -18697 10836 -18663
rect 10768 -18741 10836 -18697
rect 11000 -18515 11062 -18493
rect 11000 -18549 11026 -18515
rect 11060 -18549 11062 -18515
rect 11000 -18583 11062 -18549
rect 11000 -18619 11026 -18583
rect 11060 -18619 11062 -18583
rect 11000 -18653 11062 -18619
rect 11000 -18687 11026 -18653
rect 11060 -18687 11062 -18653
rect 11000 -18729 11062 -18687
rect 11278 -18515 11346 -18495
rect 11278 -18549 11284 -18515
rect 11318 -18549 11346 -18515
rect 11278 -18583 11346 -18549
rect 11278 -18619 11284 -18583
rect 11318 -18619 11346 -18583
rect 11278 -18653 11346 -18619
rect 11278 -18687 11284 -18653
rect 11318 -18687 11346 -18653
rect 11278 -18731 11346 -18687
rect 11637 -18527 11699 -18505
rect 11637 -18561 11663 -18527
rect 11697 -18561 11699 -18527
rect 11637 -18595 11699 -18561
rect 11637 -18631 11663 -18595
rect 11697 -18631 11699 -18595
rect 11637 -18665 11699 -18631
rect 11637 -18699 11663 -18665
rect 11697 -18699 11699 -18665
rect 10126 -18785 10140 -18751
rect 10180 -18785 10192 -18751
rect 10629 -18783 10645 -18749
rect 10679 -18783 10695 -18749
rect 11139 -18773 11155 -18739
rect 11189 -18773 11205 -18739
rect 11637 -18741 11699 -18699
rect 11915 -18527 11983 -18507
rect 11915 -18561 11921 -18527
rect 11955 -18561 11983 -18527
rect 11915 -18595 11983 -18561
rect 11915 -18631 11921 -18595
rect 11955 -18631 11983 -18595
rect 11915 -18665 11983 -18631
rect 11915 -18699 11921 -18665
rect 11955 -18699 11983 -18665
rect 11915 -18743 11983 -18699
rect 12177 -18527 12239 -18505
rect 12177 -18561 12203 -18527
rect 12237 -18561 12239 -18527
rect 12177 -18595 12239 -18561
rect 12177 -18631 12203 -18595
rect 12237 -18631 12239 -18595
rect 12177 -18665 12239 -18631
rect 12177 -18699 12203 -18665
rect 12237 -18699 12239 -18665
rect 12177 -18741 12239 -18699
rect 12455 -18527 12523 -18507
rect 12455 -18561 12461 -18527
rect 12495 -18561 12523 -18527
rect 12455 -18595 12523 -18561
rect 12455 -18631 12461 -18595
rect 12495 -18631 12523 -18595
rect 12455 -18665 12523 -18631
rect 12455 -18699 12461 -18665
rect 12495 -18699 12523 -18665
rect 12455 -18743 12523 -18699
rect 12657 -18527 12719 -18505
rect 12657 -18561 12683 -18527
rect 12717 -18561 12719 -18527
rect 12657 -18595 12719 -18561
rect 12657 -18631 12683 -18595
rect 12717 -18631 12719 -18595
rect 12657 -18665 12719 -18631
rect 12657 -18699 12683 -18665
rect 12717 -18699 12719 -18665
rect 11776 -18785 11792 -18751
rect 11826 -18785 11842 -18751
rect 12316 -18785 12332 -18751
rect 12366 -18785 12382 -18751
rect 12657 -18811 12719 -18699
rect 12935 -18527 13003 -18395
rect 13299 -18473 13315 -18439
rect 13349 -18473 13365 -18439
rect 13809 -18463 13825 -18429
rect 13859 -18463 13875 -18429
rect 14439 -18474 14455 -18440
rect 14489 -18474 14505 -18440
rect 14979 -18474 14995 -18440
rect 15029 -18474 15045 -18440
rect 15459 -18474 15470 -18440
rect 15520 -18474 15525 -18440
rect 12935 -18561 12941 -18527
rect 12975 -18561 13003 -18527
rect 12935 -18595 13003 -18561
rect 12935 -18631 12941 -18595
rect 12975 -18631 13003 -18595
rect 12935 -18665 13003 -18631
rect 12935 -18699 12941 -18665
rect 12975 -18699 13003 -18665
rect 12935 -18743 13003 -18699
rect 13160 -18525 13222 -18503
rect 13160 -18559 13186 -18525
rect 13220 -18559 13222 -18525
rect 13160 -18593 13222 -18559
rect 13160 -18629 13186 -18593
rect 13220 -18629 13222 -18593
rect 13160 -18663 13222 -18629
rect 13160 -18697 13186 -18663
rect 13220 -18697 13222 -18663
rect 13160 -18739 13222 -18697
rect 13438 -18525 13506 -18505
rect 13438 -18559 13444 -18525
rect 13478 -18559 13506 -18525
rect 13438 -18593 13506 -18559
rect 13438 -18629 13444 -18593
rect 13478 -18629 13506 -18593
rect 13438 -18663 13506 -18629
rect 13438 -18697 13444 -18663
rect 13478 -18697 13506 -18663
rect 13438 -18741 13506 -18697
rect 13670 -18515 13732 -18493
rect 13670 -18549 13696 -18515
rect 13730 -18549 13732 -18515
rect 13670 -18583 13732 -18549
rect 13670 -18619 13696 -18583
rect 13730 -18619 13732 -18583
rect 13670 -18653 13732 -18619
rect 13670 -18687 13696 -18653
rect 13730 -18687 13732 -18653
rect 13670 -18729 13732 -18687
rect 13948 -18515 14016 -18495
rect 13948 -18549 13954 -18515
rect 13988 -18549 14016 -18515
rect 13948 -18583 14016 -18549
rect 13948 -18619 13954 -18583
rect 13988 -18619 14016 -18583
rect 13948 -18653 14016 -18619
rect 13948 -18687 13954 -18653
rect 13988 -18687 14016 -18653
rect 13948 -18731 14016 -18687
rect 14300 -18526 14362 -18504
rect 14300 -18560 14326 -18526
rect 14360 -18560 14362 -18526
rect 14300 -18594 14362 -18560
rect 14300 -18630 14326 -18594
rect 14360 -18630 14362 -18594
rect 14300 -18664 14362 -18630
rect 14300 -18698 14326 -18664
rect 14360 -18698 14362 -18664
rect 12796 -18785 12810 -18751
rect 12850 -18785 12862 -18751
rect 13299 -18783 13315 -18749
rect 13349 -18783 13365 -18749
rect 13809 -18773 13825 -18739
rect 13859 -18773 13875 -18739
rect 14300 -18740 14362 -18698
rect 14578 -18526 14646 -18506
rect 14578 -18560 14584 -18526
rect 14618 -18560 14646 -18526
rect 14578 -18594 14646 -18560
rect 14578 -18630 14584 -18594
rect 14618 -18630 14646 -18594
rect 14578 -18664 14646 -18630
rect 14578 -18698 14584 -18664
rect 14618 -18698 14646 -18664
rect 14578 -18742 14646 -18698
rect 14840 -18526 14902 -18504
rect 14840 -18560 14866 -18526
rect 14900 -18560 14902 -18526
rect 14840 -18594 14902 -18560
rect 14840 -18630 14866 -18594
rect 14900 -18630 14902 -18594
rect 14840 -18664 14902 -18630
rect 14840 -18698 14866 -18664
rect 14900 -18698 14902 -18664
rect 14840 -18740 14902 -18698
rect 15118 -18526 15186 -18506
rect 15118 -18560 15124 -18526
rect 15158 -18560 15186 -18526
rect 15118 -18594 15186 -18560
rect 15118 -18630 15124 -18594
rect 15158 -18630 15186 -18594
rect 15118 -18664 15186 -18630
rect 15118 -18698 15124 -18664
rect 15158 -18698 15186 -18664
rect 15118 -18742 15186 -18698
rect 15320 -18526 15382 -18504
rect 15320 -18560 15346 -18526
rect 15380 -18560 15382 -18526
rect 15320 -18594 15382 -18560
rect 15320 -18630 15346 -18594
rect 15380 -18630 15382 -18594
rect 15320 -18664 15382 -18630
rect 15320 -18698 15346 -18664
rect 15380 -18698 15382 -18664
rect 14439 -18784 14455 -18750
rect 14489 -18784 14505 -18750
rect 14979 -18784 14995 -18750
rect 15029 -18784 15045 -18750
rect 12656 -18870 12719 -18811
rect 15320 -18870 15382 -18698
rect 15598 -18526 15666 -18351
rect 15962 -18472 15978 -18438
rect 16012 -18472 16028 -18438
rect 16472 -18462 16488 -18428
rect 16522 -18462 16538 -18428
rect 15598 -18560 15604 -18526
rect 15638 -18560 15666 -18526
rect 15598 -18594 15666 -18560
rect 15598 -18630 15604 -18594
rect 15638 -18630 15666 -18594
rect 15598 -18664 15666 -18630
rect 15598 -18698 15604 -18664
rect 15638 -18698 15666 -18664
rect 15598 -18742 15666 -18698
rect 15823 -18524 15885 -18502
rect 15823 -18558 15849 -18524
rect 15883 -18558 15885 -18524
rect 15823 -18592 15885 -18558
rect 15823 -18628 15849 -18592
rect 15883 -18628 15885 -18592
rect 15823 -18662 15885 -18628
rect 15823 -18696 15849 -18662
rect 15883 -18696 15885 -18662
rect 15823 -18738 15885 -18696
rect 16101 -18524 16169 -18504
rect 16101 -18558 16107 -18524
rect 16141 -18558 16169 -18524
rect 16101 -18592 16169 -18558
rect 16101 -18628 16107 -18592
rect 16141 -18628 16169 -18592
rect 16101 -18662 16169 -18628
rect 16101 -18696 16107 -18662
rect 16141 -18696 16169 -18662
rect 16101 -18740 16169 -18696
rect 16333 -18514 16395 -18492
rect 16333 -18548 16359 -18514
rect 16393 -18548 16395 -18514
rect 16333 -18582 16395 -18548
rect 16333 -18618 16359 -18582
rect 16393 -18618 16395 -18582
rect 16333 -18652 16395 -18618
rect 16333 -18686 16359 -18652
rect 16393 -18686 16395 -18652
rect 16333 -18728 16395 -18686
rect 16611 -18514 16679 -18494
rect 16611 -18548 16617 -18514
rect 16651 -18548 16679 -18514
rect 16611 -18582 16679 -18548
rect 16611 -18618 16617 -18582
rect 16651 -18618 16679 -18582
rect 16611 -18652 16679 -18618
rect 16611 -18686 16617 -18652
rect 16651 -18686 16679 -18652
rect 16611 -18730 16679 -18686
rect 15459 -18784 15470 -18750
rect 15512 -18784 15525 -18750
rect 15962 -18782 15978 -18748
rect 16012 -18782 16028 -18748
rect 16472 -18772 16488 -18738
rect 16522 -18772 16538 -18738
rect 8823 -18880 16813 -18870
rect 8823 -18986 9964 -18880
rect 10070 -18885 16813 -18880
rect 10070 -18979 12640 -18885
rect 12732 -18979 15306 -18885
rect 15398 -18979 16813 -18885
rect 10070 -18986 16813 -18979
rect 8823 -18990 16813 -18986
rect 12656 -18991 12718 -18990
rect 16986 -19151 17138 -18029
rect 8484 -19275 17138 -19151
rect 8951 -20123 9135 -20104
rect 8951 -20387 8970 -20123
rect 9113 -20387 9135 -20123
rect 9357 -20167 9619 -20137
rect 9664 -20167 9728 -19275
rect 12332 -20131 12396 -19275
rect 9357 -20205 9453 -20167
rect 9519 -20205 9619 -20167
rect 9357 -20291 9619 -20205
rect 9357 -20293 9561 -20291
rect 9357 -20329 9375 -20293
rect 9413 -20327 9561 -20293
rect 9599 -20327 9619 -20291
rect 9413 -20329 9619 -20327
rect 9357 -20365 9619 -20329
rect 9665 -20294 9727 -20167
rect 10698 -20169 10970 -20139
rect 10044 -20209 10060 -20175
rect 10214 -20209 10230 -20175
rect 10698 -20207 10794 -20169
rect 10860 -20207 10970 -20169
rect 9665 -20328 9691 -20294
rect 9725 -20328 9727 -20294
rect 8951 -20420 9135 -20387
rect 9665 -20399 9727 -20328
rect 10549 -20294 10594 -20278
rect 10583 -20328 10594 -20294
rect 10044 -20447 10060 -20413
rect 10214 -20447 10230 -20413
rect 10549 -20535 10594 -20328
rect 10698 -20293 10970 -20207
rect 10698 -20295 10902 -20293
rect 10698 -20331 10716 -20295
rect 10754 -20329 10902 -20295
rect 10940 -20329 10970 -20293
rect 10754 -20331 10970 -20329
rect 10698 -20367 10970 -20331
rect 11068 -20169 11340 -20139
rect 11068 -20207 11164 -20169
rect 11230 -20207 11340 -20169
rect 11068 -20293 11340 -20207
rect 11068 -20295 11272 -20293
rect 11068 -20331 11086 -20295
rect 11124 -20329 11272 -20295
rect 11310 -20329 11340 -20293
rect 11124 -20331 11340 -20329
rect 11068 -20367 11340 -20331
rect 11490 -20169 11762 -20139
rect 11490 -20207 11586 -20169
rect 11652 -20207 11762 -20169
rect 11490 -20293 11762 -20207
rect 11490 -20295 11694 -20293
rect 11490 -20331 11508 -20295
rect 11546 -20329 11694 -20295
rect 11732 -20329 11762 -20293
rect 11546 -20331 11762 -20329
rect 11490 -20367 11762 -20331
rect 11912 -20169 12184 -20139
rect 12332 -20147 12397 -20131
rect 11912 -20207 12008 -20169
rect 12074 -20207 12184 -20169
rect 11912 -20293 12184 -20207
rect 11912 -20295 12116 -20293
rect 11912 -20331 11930 -20295
rect 11968 -20329 12116 -20295
rect 12154 -20329 12184 -20293
rect 11968 -20331 12184 -20329
rect 11912 -20367 12184 -20331
rect 12335 -20294 12397 -20147
rect 13399 -20169 13671 -20139
rect 12714 -20209 12730 -20175
rect 12884 -20209 12900 -20175
rect 13399 -20207 13495 -20169
rect 13561 -20207 13671 -20169
rect 12335 -20328 12361 -20294
rect 12395 -20328 12397 -20294
rect 12335 -20399 12397 -20328
rect 13219 -20294 13264 -20278
rect 13253 -20328 13264 -20294
rect 12714 -20447 12730 -20413
rect 12884 -20447 12900 -20413
rect 13219 -20522 13264 -20328
rect 13399 -20293 13671 -20207
rect 13399 -20295 13603 -20293
rect 13399 -20331 13417 -20295
rect 13455 -20329 13603 -20295
rect 13641 -20329 13671 -20293
rect 13455 -20331 13671 -20329
rect 13399 -20367 13671 -20331
rect 13769 -20169 14041 -20139
rect 13769 -20207 13865 -20169
rect 13931 -20207 14041 -20169
rect 13769 -20293 14041 -20207
rect 13769 -20295 13973 -20293
rect 13769 -20331 13787 -20295
rect 13825 -20329 13973 -20295
rect 14011 -20329 14041 -20293
rect 13825 -20331 14041 -20329
rect 13769 -20367 14041 -20331
rect 14191 -20169 14463 -20139
rect 14191 -20207 14287 -20169
rect 14353 -20207 14463 -20169
rect 14191 -20293 14463 -20207
rect 14191 -20295 14395 -20293
rect 14191 -20331 14209 -20295
rect 14247 -20329 14395 -20295
rect 14433 -20329 14463 -20293
rect 14247 -20331 14463 -20329
rect 14191 -20367 14463 -20331
rect 14613 -20169 14885 -20139
rect 14613 -20207 14709 -20169
rect 14775 -20207 14885 -20169
rect 14613 -20293 14885 -20207
rect 14613 -20295 14817 -20293
rect 14613 -20331 14631 -20295
rect 14669 -20329 14817 -20295
rect 14855 -20329 14885 -20293
rect 14669 -20331 14885 -20329
rect 14613 -20367 14885 -20331
rect 14998 -20179 15062 -19275
rect 16233 -19577 16467 -19563
rect 16682 -19575 16698 -19541
rect 16732 -19575 16748 -19541
rect 17072 -19577 17088 -19543
rect 17122 -19577 17138 -19543
rect 16233 -19892 16247 -19577
rect 16449 -19579 16467 -19577
rect 16450 -19730 16467 -19579
rect 16654 -19634 16688 -19618
rect 16450 -19731 16512 -19730
rect 16450 -19749 16654 -19731
rect 16450 -19811 16510 -19749
rect 16566 -19811 16654 -19749
rect 16450 -19825 16654 -19811
rect 16450 -19827 16598 -19825
rect 16450 -19830 16512 -19827
rect 16233 -19893 16248 -19892
rect 16450 -19893 16467 -19830
rect 16233 -19910 16467 -19893
rect 16642 -19946 16654 -19825
rect 16642 -19962 16688 -19946
rect 16742 -19634 16776 -19618
rect 17044 -19636 17078 -19620
rect 16884 -19747 17044 -19733
rect 16884 -19819 16887 -19747
rect 16958 -19819 17044 -19747
rect 16884 -19827 17044 -19819
rect 16776 -19946 16836 -19827
rect 16884 -19829 16988 -19827
rect 16642 -19963 16676 -19962
rect 16742 -19963 16836 -19946
rect 16682 -20039 16698 -20005
rect 16732 -20039 16748 -20005
rect 16792 -20169 16836 -19963
rect 17032 -19948 17044 -19827
rect 17032 -19964 17078 -19948
rect 17132 -19636 17166 -19620
rect 17166 -19948 17226 -19829
rect 17032 -19965 17066 -19964
rect 17132 -19965 17226 -19948
rect 17072 -20041 17088 -20007
rect 17122 -20041 17138 -20007
rect 17182 -20163 17226 -19965
rect 14998 -20293 15060 -20179
rect 15377 -20208 15393 -20174
rect 15547 -20208 15563 -20174
rect 16792 -20181 16922 -20169
rect 16792 -20219 16848 -20181
rect 16902 -20219 16922 -20181
rect 16792 -20227 16922 -20219
rect 17182 -20183 17298 -20163
rect 17182 -20227 17236 -20183
rect 17284 -20227 17298 -20183
rect 14998 -20327 15024 -20293
rect 15058 -20327 15060 -20293
rect 14998 -20398 15060 -20327
rect 15882 -20293 15927 -20277
rect 15916 -20327 15927 -20293
rect 15377 -20446 15393 -20412
rect 15547 -20446 15563 -20412
rect 10549 -20914 10593 -20535
rect 10548 -20976 10593 -20914
rect 13218 -20939 13264 -20522
rect 15882 -20914 15927 -20327
rect 16686 -20371 16702 -20337
rect 16736 -20371 16752 -20337
rect 16510 -20405 16582 -20399
rect 16792 -20405 16836 -20227
rect 17182 -20243 17298 -20227
rect 17076 -20371 17092 -20337
rect 17126 -20371 17142 -20337
rect 16510 -20415 16694 -20405
rect 16510 -20488 16523 -20415
rect 16579 -20421 16694 -20415
rect 16579 -20481 16658 -20421
rect 16692 -20481 16694 -20421
rect 16579 -20488 16694 -20481
rect 16510 -20497 16694 -20488
rect 16746 -20421 16836 -20405
rect 16780 -20481 16836 -20421
rect 16746 -20497 16836 -20481
rect 16900 -20405 16972 -20399
rect 17182 -20405 17226 -20243
rect 16900 -20415 17084 -20405
rect 16900 -20488 16915 -20415
rect 16961 -20421 17084 -20415
rect 16961 -20481 17048 -20421
rect 17082 -20481 17084 -20421
rect 16961 -20488 17084 -20481
rect 16900 -20497 17084 -20488
rect 17136 -20421 17226 -20405
rect 17170 -20481 17226 -20421
rect 17136 -20497 17226 -20481
rect 16510 -20503 16582 -20497
rect 16900 -20503 16972 -20497
rect 16686 -20565 16702 -20531
rect 16736 -20565 16752 -20531
rect 17076 -20565 17092 -20531
rect 17126 -20565 17142 -20531
rect 13218 -20976 13263 -20939
rect 10548 -20987 12889 -20976
rect 10548 -21066 12755 -20987
rect 12850 -21066 12889 -20987
rect 10548 -21081 12889 -21066
rect 10548 -21083 11219 -21081
rect 12626 -21082 12889 -21081
rect 13218 -20987 15547 -20976
rect 15881 -20977 15927 -20914
rect 16496 -20699 16790 -20697
rect 16496 -20741 16842 -20699
rect 16496 -20977 16542 -20741
rect 13218 -21066 15428 -20987
rect 15523 -21066 15547 -20987
rect 13218 -21081 15547 -21066
rect 15878 -21031 16542 -20977
rect 16792 -21031 16842 -20741
rect 15878 -21067 16842 -21031
rect 13218 -21083 13894 -21081
rect 15299 -21082 15547 -21081
rect 15881 -21081 16842 -21067
rect 15881 -21082 16813 -21081
rect 9226 -21219 9242 -21185
rect 9276 -21219 9292 -21185
rect 9484 -21219 9500 -21185
rect 9534 -21219 9550 -21185
rect 9742 -21219 9758 -21185
rect 9792 -21219 9808 -21185
rect 10000 -21219 10016 -21185
rect 10050 -21219 10066 -21185
rect 10258 -21219 10274 -21185
rect 10308 -21219 10324 -21185
rect 10516 -21219 10532 -21185
rect 10566 -21219 10582 -21185
rect 10774 -21219 10790 -21185
rect 10824 -21219 10840 -21185
rect 11032 -21219 11048 -21185
rect 11082 -21219 11098 -21185
rect 9107 -21269 9152 -21225
rect 9107 -21305 9113 -21269
rect 9147 -21305 9152 -21269
rect 9107 -21339 9152 -21305
rect 9107 -21375 9113 -21339
rect 9147 -21375 9152 -21339
rect 9107 -21409 9152 -21375
rect 9107 -21445 9113 -21409
rect 9147 -21445 9152 -21409
rect 9107 -21687 9152 -21445
rect 9365 -21269 9410 -21225
rect 9365 -21305 9371 -21269
rect 9405 -21305 9410 -21269
rect 9365 -21339 9410 -21305
rect 9365 -21375 9371 -21339
rect 9405 -21375 9410 -21339
rect 9365 -21409 9410 -21375
rect 9365 -21445 9371 -21409
rect 9405 -21445 9410 -21409
rect 9226 -21529 9242 -21495
rect 9276 -21529 9292 -21495
rect 9226 -21637 9242 -21603
rect 9276 -21637 9292 -21603
rect 9107 -21723 9113 -21687
rect 9147 -21723 9152 -21687
rect 9107 -21757 9152 -21723
rect 9107 -21793 9113 -21757
rect 9147 -21793 9152 -21757
rect 9107 -21827 9152 -21793
rect 9107 -21863 9113 -21827
rect 9147 -21863 9152 -21827
rect 9107 -22105 9152 -21863
rect 9365 -21687 9410 -21445
rect 9622 -21269 9667 -21225
rect 9622 -21305 9629 -21269
rect 9663 -21305 9667 -21269
rect 9622 -21339 9667 -21305
rect 9622 -21375 9629 -21339
rect 9663 -21375 9667 -21339
rect 9622 -21410 9667 -21375
rect 9622 -21446 9629 -21410
rect 9663 -21446 9667 -21410
rect 9484 -21529 9500 -21495
rect 9534 -21529 9550 -21495
rect 9484 -21637 9500 -21603
rect 9534 -21637 9550 -21603
rect 9365 -21723 9371 -21687
rect 9405 -21723 9410 -21687
rect 9365 -21757 9410 -21723
rect 9365 -21793 9371 -21757
rect 9405 -21793 9410 -21757
rect 9365 -21827 9410 -21793
rect 9365 -21863 9371 -21827
rect 9405 -21863 9410 -21827
rect 9226 -21947 9242 -21913
rect 9276 -21947 9292 -21913
rect 9226 -22055 9242 -22021
rect 9276 -22055 9292 -22021
rect 9107 -22141 9113 -22105
rect 9147 -22141 9152 -22105
rect 9107 -22175 9152 -22141
rect 9107 -22211 9113 -22175
rect 9147 -22211 9152 -22175
rect 9107 -22245 9152 -22211
rect 9107 -22281 9113 -22245
rect 9147 -22281 9152 -22245
rect 9107 -22523 9152 -22281
rect 9365 -22105 9410 -21863
rect 9622 -21687 9667 -21446
rect 9882 -21269 9927 -21225
rect 9882 -21305 9887 -21269
rect 9921 -21305 9927 -21269
rect 9882 -21339 9927 -21305
rect 9882 -21375 9887 -21339
rect 9921 -21375 9927 -21339
rect 9882 -21409 9927 -21375
rect 9882 -21445 9887 -21409
rect 9921 -21445 9927 -21409
rect 9742 -21529 9758 -21495
rect 9792 -21529 9808 -21495
rect 9742 -21637 9758 -21603
rect 9792 -21637 9808 -21603
rect 9622 -21723 9629 -21687
rect 9663 -21723 9667 -21687
rect 9622 -21757 9667 -21723
rect 9622 -21793 9629 -21757
rect 9663 -21793 9667 -21757
rect 9622 -21828 9667 -21793
rect 9622 -21864 9629 -21828
rect 9663 -21864 9667 -21828
rect 9484 -21947 9500 -21913
rect 9534 -21947 9550 -21913
rect 9484 -22055 9500 -22021
rect 9534 -22055 9550 -22021
rect 9365 -22141 9371 -22105
rect 9405 -22141 9410 -22105
rect 9365 -22175 9410 -22141
rect 9365 -22211 9371 -22175
rect 9405 -22211 9410 -22175
rect 9365 -22245 9410 -22211
rect 9365 -22281 9371 -22245
rect 9405 -22281 9410 -22245
rect 9226 -22365 9242 -22331
rect 9276 -22365 9292 -22331
rect 9226 -22473 9242 -22439
rect 9276 -22473 9292 -22439
rect 9107 -22559 9113 -22523
rect 9147 -22559 9152 -22523
rect 9107 -22593 9152 -22559
rect 9107 -22629 9113 -22593
rect 9147 -22629 9152 -22593
rect 9107 -22663 9152 -22629
rect 9107 -22699 9113 -22663
rect 9147 -22699 9152 -22663
rect 9107 -22941 9152 -22699
rect 9365 -22523 9410 -22281
rect 9622 -22105 9667 -21864
rect 9882 -21687 9927 -21445
rect 10140 -21269 10185 -21225
rect 10140 -21305 10145 -21269
rect 10179 -21305 10185 -21269
rect 10140 -21339 10185 -21305
rect 10140 -21375 10145 -21339
rect 10179 -21375 10185 -21339
rect 10140 -21409 10185 -21375
rect 10140 -21445 10145 -21409
rect 10179 -21445 10185 -21409
rect 10000 -21529 10016 -21495
rect 10050 -21529 10066 -21495
rect 10000 -21637 10016 -21603
rect 10050 -21637 10066 -21603
rect 9882 -21723 9887 -21687
rect 9921 -21723 9927 -21687
rect 9882 -21757 9927 -21723
rect 9882 -21793 9887 -21757
rect 9921 -21793 9927 -21757
rect 9882 -21827 9927 -21793
rect 9882 -21863 9887 -21827
rect 9921 -21863 9927 -21827
rect 9742 -21947 9758 -21913
rect 9792 -21947 9808 -21913
rect 9742 -22055 9758 -22021
rect 9792 -22055 9808 -22021
rect 9622 -22141 9629 -22105
rect 9663 -22141 9667 -22105
rect 9622 -22175 9667 -22141
rect 9622 -22211 9629 -22175
rect 9663 -22211 9667 -22175
rect 9622 -22246 9667 -22211
rect 9622 -22282 9629 -22246
rect 9663 -22282 9667 -22246
rect 9484 -22365 9500 -22331
rect 9534 -22365 9550 -22331
rect 9484 -22473 9500 -22439
rect 9534 -22473 9550 -22439
rect 9365 -22559 9371 -22523
rect 9405 -22559 9410 -22523
rect 9365 -22593 9410 -22559
rect 9365 -22629 9371 -22593
rect 9405 -22629 9410 -22593
rect 9365 -22663 9410 -22629
rect 9365 -22699 9371 -22663
rect 9405 -22699 9410 -22663
rect 9226 -22783 9242 -22749
rect 9276 -22783 9292 -22749
rect 9226 -22891 9242 -22857
rect 9276 -22891 9292 -22857
rect 9107 -22977 9113 -22941
rect 9147 -22977 9152 -22941
rect 9107 -23011 9152 -22977
rect 9107 -23047 9113 -23011
rect 9147 -23047 9152 -23011
rect 9107 -23081 9152 -23047
rect 9107 -23117 9113 -23081
rect 9147 -23117 9152 -23081
rect 9107 -23359 9152 -23117
rect 9365 -22941 9410 -22699
rect 9622 -22523 9667 -22282
rect 9882 -22105 9927 -21863
rect 10140 -21687 10185 -21445
rect 10397 -21269 10442 -21225
rect 10397 -21305 10403 -21269
rect 10437 -21305 10442 -21269
rect 10397 -21339 10442 -21305
rect 10397 -21375 10403 -21339
rect 10437 -21375 10442 -21339
rect 10397 -21409 10442 -21375
rect 10397 -21445 10403 -21409
rect 10437 -21445 10442 -21409
rect 10258 -21529 10274 -21495
rect 10308 -21529 10324 -21495
rect 10258 -21637 10274 -21603
rect 10308 -21637 10324 -21603
rect 10140 -21723 10145 -21687
rect 10179 -21723 10185 -21687
rect 10140 -21757 10185 -21723
rect 10140 -21793 10145 -21757
rect 10179 -21793 10185 -21757
rect 10140 -21827 10185 -21793
rect 10140 -21863 10145 -21827
rect 10179 -21863 10185 -21827
rect 10000 -21947 10016 -21913
rect 10050 -21947 10066 -21913
rect 10000 -22055 10016 -22021
rect 10050 -22055 10066 -22021
rect 9882 -22141 9887 -22105
rect 9921 -22141 9927 -22105
rect 9882 -22175 9927 -22141
rect 9882 -22211 9887 -22175
rect 9921 -22211 9927 -22175
rect 9882 -22245 9927 -22211
rect 9882 -22281 9887 -22245
rect 9921 -22281 9927 -22245
rect 9742 -22365 9758 -22331
rect 9792 -22365 9808 -22331
rect 9742 -22473 9758 -22439
rect 9792 -22473 9808 -22439
rect 9622 -22559 9629 -22523
rect 9663 -22559 9667 -22523
rect 9622 -22593 9667 -22559
rect 9622 -22629 9629 -22593
rect 9663 -22629 9667 -22593
rect 9622 -22664 9667 -22629
rect 9622 -22700 9629 -22664
rect 9663 -22700 9667 -22664
rect 9484 -22783 9500 -22749
rect 9534 -22783 9550 -22749
rect 9484 -22891 9500 -22857
rect 9534 -22891 9550 -22857
rect 9365 -22977 9371 -22941
rect 9405 -22977 9410 -22941
rect 9365 -23011 9410 -22977
rect 9365 -23047 9371 -23011
rect 9405 -23047 9410 -23011
rect 9365 -23081 9410 -23047
rect 9365 -23117 9371 -23081
rect 9405 -23117 9410 -23081
rect 9226 -23201 9242 -23167
rect 9276 -23201 9292 -23167
rect 9226 -23309 9242 -23275
rect 9276 -23309 9292 -23275
rect 9107 -23395 9113 -23359
rect 9147 -23395 9152 -23359
rect 9107 -23429 9152 -23395
rect 9107 -23465 9113 -23429
rect 9147 -23465 9152 -23429
rect 9107 -23499 9152 -23465
rect 9107 -23535 9113 -23499
rect 9147 -23535 9152 -23499
rect 9107 -23777 9152 -23535
rect 9365 -23359 9410 -23117
rect 9622 -22941 9667 -22700
rect 9882 -22523 9927 -22281
rect 10140 -22105 10185 -21863
rect 10397 -21687 10442 -21445
rect 10654 -21269 10699 -21225
rect 10654 -21305 10661 -21269
rect 10695 -21305 10699 -21269
rect 10654 -21339 10699 -21305
rect 10654 -21375 10661 -21339
rect 10695 -21375 10699 -21339
rect 10654 -21409 10699 -21375
rect 10654 -21445 10661 -21409
rect 10695 -21445 10699 -21409
rect 10516 -21529 10532 -21495
rect 10566 -21529 10582 -21495
rect 10516 -21637 10532 -21603
rect 10566 -21637 10582 -21603
rect 10397 -21723 10403 -21687
rect 10437 -21723 10442 -21687
rect 10397 -21757 10442 -21723
rect 10397 -21793 10403 -21757
rect 10437 -21793 10442 -21757
rect 10397 -21827 10442 -21793
rect 10397 -21863 10403 -21827
rect 10437 -21863 10442 -21827
rect 10258 -21947 10274 -21913
rect 10308 -21947 10324 -21913
rect 10258 -22055 10274 -22021
rect 10308 -22055 10324 -22021
rect 10140 -22141 10145 -22105
rect 10179 -22141 10185 -22105
rect 10140 -22175 10185 -22141
rect 10140 -22211 10145 -22175
rect 10179 -22211 10185 -22175
rect 10140 -22245 10185 -22211
rect 10140 -22281 10145 -22245
rect 10179 -22281 10185 -22245
rect 10000 -22365 10016 -22331
rect 10050 -22365 10066 -22331
rect 10000 -22473 10016 -22439
rect 10050 -22473 10066 -22439
rect 9882 -22559 9887 -22523
rect 9921 -22559 9927 -22523
rect 9882 -22593 9927 -22559
rect 9882 -22629 9887 -22593
rect 9921 -22629 9927 -22593
rect 9882 -22663 9927 -22629
rect 9882 -22699 9887 -22663
rect 9921 -22699 9927 -22663
rect 9742 -22783 9758 -22749
rect 9792 -22783 9808 -22749
rect 9742 -22891 9758 -22857
rect 9792 -22891 9808 -22857
rect 9622 -22977 9629 -22941
rect 9663 -22977 9667 -22941
rect 9622 -23011 9667 -22977
rect 9622 -23047 9629 -23011
rect 9663 -23047 9667 -23011
rect 9622 -23082 9667 -23047
rect 9622 -23118 9629 -23082
rect 9663 -23118 9667 -23082
rect 9484 -23201 9500 -23167
rect 9534 -23201 9550 -23167
rect 9484 -23309 9500 -23275
rect 9534 -23309 9550 -23275
rect 9365 -23395 9371 -23359
rect 9405 -23395 9410 -23359
rect 9365 -23429 9410 -23395
rect 9365 -23465 9371 -23429
rect 9405 -23465 9410 -23429
rect 9365 -23499 9410 -23465
rect 9365 -23535 9371 -23499
rect 9405 -23535 9410 -23499
rect 9226 -23619 9242 -23585
rect 9276 -23619 9292 -23585
rect 9226 -23727 9242 -23693
rect 9276 -23727 9292 -23693
rect 9107 -23813 9113 -23777
rect 9147 -23813 9152 -23777
rect 9107 -23847 9152 -23813
rect 9107 -23883 9113 -23847
rect 9147 -23883 9152 -23847
rect 9107 -23917 9152 -23883
rect 9107 -23953 9113 -23917
rect 9147 -23953 9152 -23917
rect 9107 -24195 9152 -23953
rect 9365 -23777 9410 -23535
rect 9622 -23359 9667 -23118
rect 9882 -22941 9927 -22699
rect 10140 -22523 10185 -22281
rect 10397 -22105 10442 -21863
rect 10654 -21687 10699 -21445
rect 10913 -21269 10958 -21225
rect 10913 -21305 10919 -21269
rect 10953 -21305 10958 -21269
rect 10913 -21339 10958 -21305
rect 10913 -21375 10919 -21339
rect 10953 -21375 10958 -21339
rect 10913 -21409 10958 -21375
rect 10913 -21445 10919 -21409
rect 10953 -21445 10958 -21409
rect 10774 -21529 10790 -21495
rect 10824 -21529 10840 -21495
rect 10774 -21637 10790 -21603
rect 10824 -21637 10840 -21603
rect 10654 -21723 10661 -21687
rect 10695 -21723 10699 -21687
rect 10654 -21757 10699 -21723
rect 10654 -21793 10661 -21757
rect 10695 -21793 10699 -21757
rect 10654 -21827 10699 -21793
rect 10654 -21863 10661 -21827
rect 10695 -21863 10699 -21827
rect 10516 -21947 10532 -21913
rect 10566 -21947 10582 -21913
rect 10516 -22055 10532 -22021
rect 10566 -22055 10582 -22021
rect 10397 -22141 10403 -22105
rect 10437 -22141 10442 -22105
rect 10397 -22175 10442 -22141
rect 10397 -22211 10403 -22175
rect 10437 -22211 10442 -22175
rect 10397 -22245 10442 -22211
rect 10397 -22281 10403 -22245
rect 10437 -22281 10442 -22245
rect 10258 -22365 10274 -22331
rect 10308 -22365 10324 -22331
rect 10258 -22473 10274 -22439
rect 10308 -22473 10324 -22439
rect 10140 -22559 10145 -22523
rect 10179 -22559 10185 -22523
rect 10140 -22593 10185 -22559
rect 10140 -22629 10145 -22593
rect 10179 -22629 10185 -22593
rect 10140 -22663 10185 -22629
rect 10140 -22699 10145 -22663
rect 10179 -22699 10185 -22663
rect 10000 -22783 10016 -22749
rect 10050 -22783 10066 -22749
rect 10000 -22891 10016 -22857
rect 10050 -22891 10066 -22857
rect 9882 -22977 9887 -22941
rect 9921 -22977 9927 -22941
rect 9882 -23011 9927 -22977
rect 9882 -23047 9887 -23011
rect 9921 -23047 9927 -23011
rect 9882 -23081 9927 -23047
rect 9882 -23117 9887 -23081
rect 9921 -23117 9927 -23081
rect 9742 -23201 9758 -23167
rect 9792 -23201 9808 -23167
rect 9742 -23309 9758 -23275
rect 9792 -23309 9808 -23275
rect 9622 -23395 9629 -23359
rect 9663 -23395 9667 -23359
rect 9622 -23429 9667 -23395
rect 9622 -23465 9629 -23429
rect 9663 -23465 9667 -23429
rect 9622 -23500 9667 -23465
rect 9622 -23536 9629 -23500
rect 9663 -23536 9667 -23500
rect 9484 -23619 9500 -23585
rect 9534 -23619 9550 -23585
rect 9484 -23727 9500 -23693
rect 9534 -23727 9550 -23693
rect 9365 -23813 9371 -23777
rect 9405 -23813 9410 -23777
rect 9365 -23847 9410 -23813
rect 9365 -23883 9371 -23847
rect 9405 -23883 9410 -23847
rect 9365 -23917 9410 -23883
rect 9365 -23953 9371 -23917
rect 9405 -23953 9410 -23917
rect 9226 -24037 9242 -24003
rect 9276 -24037 9292 -24003
rect 9365 -24071 9410 -23953
rect 9622 -23777 9667 -23536
rect 9882 -23359 9927 -23117
rect 10140 -22941 10185 -22699
rect 10397 -22523 10442 -22281
rect 10654 -22105 10699 -21863
rect 10913 -21687 10958 -21445
rect 11171 -21269 11216 -21083
rect 11896 -21219 11912 -21185
rect 11946 -21219 11962 -21185
rect 12154 -21219 12170 -21185
rect 12204 -21219 12220 -21185
rect 12412 -21219 12428 -21185
rect 12462 -21219 12478 -21185
rect 12670 -21219 12686 -21185
rect 12720 -21219 12736 -21185
rect 12928 -21219 12944 -21185
rect 12978 -21219 12994 -21185
rect 13186 -21219 13202 -21185
rect 13236 -21219 13252 -21185
rect 13444 -21219 13460 -21185
rect 13494 -21219 13510 -21185
rect 13702 -21219 13718 -21185
rect 13752 -21219 13768 -21185
rect 11171 -21305 11177 -21269
rect 11211 -21305 11216 -21269
rect 11171 -21339 11216 -21305
rect 11171 -21375 11177 -21339
rect 11211 -21375 11216 -21339
rect 11171 -21409 11216 -21375
rect 11171 -21445 11177 -21409
rect 11211 -21445 11216 -21409
rect 11032 -21529 11048 -21495
rect 11082 -21529 11098 -21495
rect 11032 -21637 11048 -21603
rect 11082 -21637 11098 -21603
rect 10913 -21723 10919 -21687
rect 10953 -21723 10958 -21687
rect 10913 -21757 10958 -21723
rect 10913 -21793 10919 -21757
rect 10953 -21793 10958 -21757
rect 10913 -21827 10958 -21793
rect 10913 -21863 10919 -21827
rect 10953 -21863 10958 -21827
rect 10774 -21947 10790 -21913
rect 10824 -21947 10840 -21913
rect 10774 -22055 10790 -22021
rect 10824 -22055 10840 -22021
rect 10654 -22141 10661 -22105
rect 10695 -22141 10699 -22105
rect 10654 -22175 10699 -22141
rect 10654 -22211 10661 -22175
rect 10695 -22211 10699 -22175
rect 10654 -22245 10699 -22211
rect 10654 -22281 10661 -22245
rect 10695 -22281 10699 -22245
rect 10516 -22365 10532 -22331
rect 10566 -22365 10582 -22331
rect 10516 -22473 10532 -22439
rect 10566 -22473 10582 -22439
rect 10397 -22559 10403 -22523
rect 10437 -22559 10442 -22523
rect 10397 -22593 10442 -22559
rect 10397 -22629 10403 -22593
rect 10437 -22629 10442 -22593
rect 10397 -22663 10442 -22629
rect 10397 -22699 10403 -22663
rect 10437 -22699 10442 -22663
rect 10258 -22783 10274 -22749
rect 10308 -22783 10324 -22749
rect 10258 -22891 10274 -22857
rect 10308 -22891 10324 -22857
rect 10140 -22977 10145 -22941
rect 10179 -22977 10185 -22941
rect 10140 -23011 10185 -22977
rect 10140 -23047 10145 -23011
rect 10179 -23047 10185 -23011
rect 10140 -23081 10185 -23047
rect 10140 -23117 10145 -23081
rect 10179 -23117 10185 -23081
rect 10000 -23201 10016 -23167
rect 10050 -23201 10066 -23167
rect 10000 -23309 10016 -23275
rect 10050 -23309 10066 -23275
rect 9882 -23395 9887 -23359
rect 9921 -23395 9927 -23359
rect 9882 -23429 9927 -23395
rect 9882 -23465 9887 -23429
rect 9921 -23465 9927 -23429
rect 9882 -23499 9927 -23465
rect 9882 -23535 9887 -23499
rect 9921 -23535 9927 -23499
rect 9742 -23619 9758 -23585
rect 9792 -23619 9808 -23585
rect 9742 -23727 9758 -23693
rect 9792 -23727 9808 -23693
rect 9622 -23813 9629 -23777
rect 9663 -23813 9667 -23777
rect 9622 -23847 9667 -23813
rect 9622 -23883 9629 -23847
rect 9663 -23883 9667 -23847
rect 9622 -23918 9667 -23883
rect 9622 -23954 9629 -23918
rect 9663 -23954 9667 -23918
rect 9484 -24037 9500 -24003
rect 9534 -24037 9550 -24003
rect 9622 -24071 9667 -23954
rect 9882 -23777 9927 -23535
rect 10140 -23359 10185 -23117
rect 10397 -22941 10442 -22699
rect 10654 -22523 10699 -22281
rect 10913 -22105 10958 -21863
rect 11171 -21687 11216 -21445
rect 11171 -21723 11177 -21687
rect 11211 -21723 11216 -21687
rect 11171 -21757 11216 -21723
rect 11171 -21793 11177 -21757
rect 11211 -21793 11216 -21757
rect 11171 -21827 11216 -21793
rect 11171 -21863 11177 -21827
rect 11211 -21863 11216 -21827
rect 11032 -21947 11048 -21913
rect 11082 -21947 11098 -21913
rect 11032 -22055 11048 -22021
rect 11082 -22055 11098 -22021
rect 10913 -22141 10919 -22105
rect 10953 -22141 10958 -22105
rect 10913 -22175 10958 -22141
rect 10913 -22211 10919 -22175
rect 10953 -22211 10958 -22175
rect 10913 -22245 10958 -22211
rect 10913 -22281 10919 -22245
rect 10953 -22281 10958 -22245
rect 10774 -22365 10790 -22331
rect 10824 -22365 10840 -22331
rect 10774 -22473 10790 -22439
rect 10824 -22473 10840 -22439
rect 10654 -22559 10661 -22523
rect 10695 -22559 10699 -22523
rect 10654 -22593 10699 -22559
rect 10654 -22629 10661 -22593
rect 10695 -22629 10699 -22593
rect 10654 -22663 10699 -22629
rect 10654 -22699 10661 -22663
rect 10695 -22699 10699 -22663
rect 10516 -22783 10532 -22749
rect 10566 -22783 10582 -22749
rect 10516 -22891 10532 -22857
rect 10566 -22891 10582 -22857
rect 10397 -22977 10403 -22941
rect 10437 -22977 10442 -22941
rect 10397 -23011 10442 -22977
rect 10397 -23047 10403 -23011
rect 10437 -23047 10442 -23011
rect 10397 -23081 10442 -23047
rect 10397 -23117 10403 -23081
rect 10437 -23117 10442 -23081
rect 10258 -23201 10274 -23167
rect 10308 -23201 10324 -23167
rect 10258 -23309 10274 -23275
rect 10308 -23309 10324 -23275
rect 10140 -23395 10145 -23359
rect 10179 -23395 10185 -23359
rect 10140 -23429 10185 -23395
rect 10140 -23465 10145 -23429
rect 10179 -23465 10185 -23429
rect 10140 -23499 10185 -23465
rect 10140 -23535 10145 -23499
rect 10179 -23535 10185 -23499
rect 10000 -23619 10016 -23585
rect 10050 -23619 10066 -23585
rect 10000 -23727 10016 -23693
rect 10050 -23727 10066 -23693
rect 9882 -23813 9887 -23777
rect 9921 -23813 9927 -23777
rect 9882 -23847 9927 -23813
rect 9882 -23883 9887 -23847
rect 9921 -23883 9927 -23847
rect 9882 -23917 9927 -23883
rect 9882 -23953 9887 -23917
rect 9921 -23953 9927 -23917
rect 9742 -24037 9758 -24003
rect 9792 -24037 9808 -24003
rect 9882 -24071 9927 -23953
rect 10140 -23777 10185 -23535
rect 10397 -23359 10442 -23117
rect 10654 -22941 10699 -22699
rect 10913 -22523 10958 -22281
rect 11171 -22105 11216 -21863
rect 11171 -22141 11177 -22105
rect 11211 -22141 11216 -22105
rect 11171 -22175 11216 -22141
rect 11171 -22211 11177 -22175
rect 11211 -22211 11216 -22175
rect 11171 -22245 11216 -22211
rect 11171 -22281 11177 -22245
rect 11211 -22281 11216 -22245
rect 11032 -22365 11048 -22331
rect 11082 -22365 11098 -22331
rect 11032 -22473 11048 -22439
rect 11082 -22473 11098 -22439
rect 10913 -22559 10919 -22523
rect 10953 -22559 10958 -22523
rect 10913 -22593 10958 -22559
rect 10913 -22629 10919 -22593
rect 10953 -22629 10958 -22593
rect 10913 -22663 10958 -22629
rect 10913 -22699 10919 -22663
rect 10953 -22699 10958 -22663
rect 10774 -22783 10790 -22749
rect 10824 -22783 10840 -22749
rect 10774 -22891 10790 -22857
rect 10824 -22891 10840 -22857
rect 10654 -22977 10661 -22941
rect 10695 -22977 10699 -22941
rect 10654 -23011 10699 -22977
rect 10654 -23047 10661 -23011
rect 10695 -23047 10699 -23011
rect 10654 -23081 10699 -23047
rect 10654 -23117 10661 -23081
rect 10695 -23117 10699 -23081
rect 10516 -23201 10532 -23167
rect 10566 -23201 10582 -23167
rect 10516 -23309 10532 -23275
rect 10566 -23309 10582 -23275
rect 10397 -23395 10403 -23359
rect 10437 -23395 10442 -23359
rect 10397 -23429 10442 -23395
rect 10397 -23465 10403 -23429
rect 10437 -23465 10442 -23429
rect 10397 -23499 10442 -23465
rect 10397 -23535 10403 -23499
rect 10437 -23535 10442 -23499
rect 10258 -23619 10274 -23585
rect 10308 -23619 10324 -23585
rect 10258 -23727 10274 -23693
rect 10308 -23727 10324 -23693
rect 10140 -23813 10145 -23777
rect 10179 -23813 10185 -23777
rect 10140 -23847 10185 -23813
rect 10140 -23883 10145 -23847
rect 10179 -23883 10185 -23847
rect 10140 -23917 10185 -23883
rect 10140 -23953 10145 -23917
rect 10179 -23953 10185 -23917
rect 10000 -24037 10016 -24003
rect 10050 -24037 10066 -24003
rect 10140 -24071 10185 -23953
rect 10397 -23777 10442 -23535
rect 10654 -23359 10699 -23117
rect 10913 -22941 10958 -22699
rect 11171 -22523 11216 -22281
rect 11171 -22559 11177 -22523
rect 11211 -22559 11216 -22523
rect 11171 -22593 11216 -22559
rect 11171 -22629 11177 -22593
rect 11211 -22629 11216 -22593
rect 11171 -22663 11216 -22629
rect 11171 -22699 11177 -22663
rect 11211 -22699 11216 -22663
rect 11032 -22783 11048 -22749
rect 11082 -22783 11098 -22749
rect 11032 -22891 11048 -22857
rect 11082 -22891 11098 -22857
rect 10913 -22977 10919 -22941
rect 10953 -22977 10958 -22941
rect 10913 -23011 10958 -22977
rect 10913 -23047 10919 -23011
rect 10953 -23047 10958 -23011
rect 10913 -23081 10958 -23047
rect 10913 -23117 10919 -23081
rect 10953 -23117 10958 -23081
rect 10774 -23201 10790 -23167
rect 10824 -23201 10840 -23167
rect 10774 -23309 10790 -23275
rect 10824 -23309 10840 -23275
rect 10654 -23395 10661 -23359
rect 10695 -23395 10699 -23359
rect 10654 -23429 10699 -23395
rect 10654 -23465 10661 -23429
rect 10695 -23465 10699 -23429
rect 10654 -23499 10699 -23465
rect 10654 -23535 10661 -23499
rect 10695 -23535 10699 -23499
rect 10516 -23619 10532 -23585
rect 10566 -23619 10582 -23585
rect 10516 -23727 10532 -23693
rect 10566 -23727 10582 -23693
rect 10397 -23813 10403 -23777
rect 10437 -23813 10442 -23777
rect 10397 -23847 10442 -23813
rect 10397 -23883 10403 -23847
rect 10437 -23883 10442 -23847
rect 10397 -23917 10442 -23883
rect 10397 -23953 10403 -23917
rect 10437 -23953 10442 -23917
rect 10258 -24037 10274 -24003
rect 10308 -24037 10324 -24003
rect 10397 -24071 10442 -23953
rect 10654 -23777 10699 -23535
rect 10913 -23359 10958 -23117
rect 11171 -22941 11216 -22699
rect 11171 -22977 11177 -22941
rect 11211 -22977 11216 -22941
rect 11171 -23011 11216 -22977
rect 11171 -23047 11177 -23011
rect 11211 -23047 11216 -23011
rect 11171 -23081 11216 -23047
rect 11171 -23117 11177 -23081
rect 11211 -23117 11216 -23081
rect 11032 -23201 11048 -23167
rect 11082 -23201 11098 -23167
rect 11032 -23309 11048 -23275
rect 11082 -23309 11098 -23275
rect 10913 -23395 10919 -23359
rect 10953 -23395 10958 -23359
rect 10913 -23429 10958 -23395
rect 10913 -23465 10919 -23429
rect 10953 -23465 10958 -23429
rect 10913 -23499 10958 -23465
rect 10913 -23535 10919 -23499
rect 10953 -23535 10958 -23499
rect 10774 -23619 10790 -23585
rect 10824 -23619 10840 -23585
rect 10774 -23727 10790 -23693
rect 10824 -23727 10840 -23693
rect 10654 -23813 10661 -23777
rect 10695 -23813 10699 -23777
rect 10654 -23847 10699 -23813
rect 10654 -23883 10661 -23847
rect 10695 -23883 10699 -23847
rect 10654 -23917 10699 -23883
rect 10654 -23953 10661 -23917
rect 10695 -23953 10699 -23917
rect 10516 -24037 10532 -24003
rect 10566 -24037 10582 -24003
rect 10654 -24071 10699 -23953
rect 10913 -23777 10958 -23535
rect 11171 -23359 11216 -23117
rect 11171 -23395 11177 -23359
rect 11211 -23395 11216 -23359
rect 11171 -23429 11216 -23395
rect 11171 -23465 11177 -23429
rect 11211 -23465 11216 -23429
rect 11171 -23499 11216 -23465
rect 11171 -23535 11177 -23499
rect 11211 -23535 11216 -23499
rect 11032 -23619 11048 -23585
rect 11082 -23619 11098 -23585
rect 11032 -23727 11048 -23693
rect 11082 -23727 11098 -23693
rect 10913 -23813 10919 -23777
rect 10953 -23813 10958 -23777
rect 10913 -23847 10958 -23813
rect 10913 -23883 10919 -23847
rect 10953 -23883 10958 -23847
rect 10913 -23917 10958 -23883
rect 10913 -23953 10919 -23917
rect 10953 -23953 10958 -23917
rect 10774 -24037 10790 -24003
rect 10824 -24037 10840 -24003
rect 10913 -24071 10958 -23953
rect 11171 -23777 11216 -23535
rect 11171 -23813 11177 -23777
rect 11211 -23813 11216 -23777
rect 11171 -23847 11216 -23813
rect 11171 -23883 11177 -23847
rect 11211 -23883 11216 -23847
rect 11171 -23917 11216 -23883
rect 11171 -23953 11177 -23917
rect 11211 -23953 11216 -23917
rect 11032 -24037 11048 -24003
rect 11082 -24037 11098 -24003
rect 11171 -24071 11216 -23953
rect 11777 -21269 11822 -21225
rect 11777 -21305 11783 -21269
rect 11817 -21305 11822 -21269
rect 11777 -21339 11822 -21305
rect 11777 -21375 11783 -21339
rect 11817 -21375 11822 -21339
rect 11777 -21409 11822 -21375
rect 11777 -21445 11783 -21409
rect 11817 -21445 11822 -21409
rect 11777 -21687 11822 -21445
rect 12035 -21269 12080 -21225
rect 12035 -21305 12041 -21269
rect 12075 -21305 12080 -21269
rect 12035 -21339 12080 -21305
rect 12035 -21375 12041 -21339
rect 12075 -21375 12080 -21339
rect 12035 -21409 12080 -21375
rect 12035 -21445 12041 -21409
rect 12075 -21445 12080 -21409
rect 11896 -21529 11912 -21495
rect 11946 -21529 11962 -21495
rect 11896 -21637 11912 -21603
rect 11946 -21637 11962 -21603
rect 11777 -21723 11783 -21687
rect 11817 -21723 11822 -21687
rect 11777 -21757 11822 -21723
rect 11777 -21793 11783 -21757
rect 11817 -21793 11822 -21757
rect 11777 -21827 11822 -21793
rect 11777 -21863 11783 -21827
rect 11817 -21863 11822 -21827
rect 11777 -22105 11822 -21863
rect 12035 -21687 12080 -21445
rect 12292 -21269 12337 -21225
rect 12292 -21305 12299 -21269
rect 12333 -21305 12337 -21269
rect 12292 -21339 12337 -21305
rect 12292 -21375 12299 -21339
rect 12333 -21375 12337 -21339
rect 12292 -21410 12337 -21375
rect 12292 -21446 12299 -21410
rect 12333 -21446 12337 -21410
rect 12154 -21529 12170 -21495
rect 12204 -21529 12220 -21495
rect 12154 -21637 12170 -21603
rect 12204 -21637 12220 -21603
rect 12035 -21723 12041 -21687
rect 12075 -21723 12080 -21687
rect 12035 -21757 12080 -21723
rect 12035 -21793 12041 -21757
rect 12075 -21793 12080 -21757
rect 12035 -21827 12080 -21793
rect 12035 -21863 12041 -21827
rect 12075 -21863 12080 -21827
rect 11896 -21947 11912 -21913
rect 11946 -21947 11962 -21913
rect 11896 -22055 11912 -22021
rect 11946 -22055 11962 -22021
rect 11777 -22141 11783 -22105
rect 11817 -22141 11822 -22105
rect 11777 -22175 11822 -22141
rect 11777 -22211 11783 -22175
rect 11817 -22211 11822 -22175
rect 11777 -22245 11822 -22211
rect 11777 -22281 11783 -22245
rect 11817 -22281 11822 -22245
rect 11777 -22523 11822 -22281
rect 12035 -22105 12080 -21863
rect 12292 -21687 12337 -21446
rect 12552 -21269 12597 -21225
rect 12552 -21305 12557 -21269
rect 12591 -21305 12597 -21269
rect 12552 -21339 12597 -21305
rect 12552 -21375 12557 -21339
rect 12591 -21375 12597 -21339
rect 12552 -21409 12597 -21375
rect 12552 -21445 12557 -21409
rect 12591 -21445 12597 -21409
rect 12412 -21529 12428 -21495
rect 12462 -21529 12478 -21495
rect 12412 -21637 12428 -21603
rect 12462 -21637 12478 -21603
rect 12292 -21723 12299 -21687
rect 12333 -21723 12337 -21687
rect 12292 -21757 12337 -21723
rect 12292 -21793 12299 -21757
rect 12333 -21793 12337 -21757
rect 12292 -21828 12337 -21793
rect 12292 -21864 12299 -21828
rect 12333 -21864 12337 -21828
rect 12154 -21947 12170 -21913
rect 12204 -21947 12220 -21913
rect 12154 -22055 12170 -22021
rect 12204 -22055 12220 -22021
rect 12035 -22141 12041 -22105
rect 12075 -22141 12080 -22105
rect 12035 -22175 12080 -22141
rect 12035 -22211 12041 -22175
rect 12075 -22211 12080 -22175
rect 12035 -22245 12080 -22211
rect 12035 -22281 12041 -22245
rect 12075 -22281 12080 -22245
rect 11896 -22365 11912 -22331
rect 11946 -22365 11962 -22331
rect 11896 -22473 11912 -22439
rect 11946 -22473 11962 -22439
rect 11777 -22559 11783 -22523
rect 11817 -22559 11822 -22523
rect 11777 -22593 11822 -22559
rect 11777 -22629 11783 -22593
rect 11817 -22629 11822 -22593
rect 11777 -22663 11822 -22629
rect 11777 -22699 11783 -22663
rect 11817 -22699 11822 -22663
rect 11777 -22941 11822 -22699
rect 12035 -22523 12080 -22281
rect 12292 -22105 12337 -21864
rect 12552 -21687 12597 -21445
rect 12810 -21269 12855 -21225
rect 12810 -21305 12815 -21269
rect 12849 -21305 12855 -21269
rect 12810 -21339 12855 -21305
rect 12810 -21375 12815 -21339
rect 12849 -21375 12855 -21339
rect 12810 -21409 12855 -21375
rect 12810 -21445 12815 -21409
rect 12849 -21445 12855 -21409
rect 12670 -21529 12686 -21495
rect 12720 -21529 12736 -21495
rect 12670 -21637 12686 -21603
rect 12720 -21637 12736 -21603
rect 12552 -21723 12557 -21687
rect 12591 -21723 12597 -21687
rect 12552 -21757 12597 -21723
rect 12552 -21793 12557 -21757
rect 12591 -21793 12597 -21757
rect 12552 -21827 12597 -21793
rect 12552 -21863 12557 -21827
rect 12591 -21863 12597 -21827
rect 12412 -21947 12428 -21913
rect 12462 -21947 12478 -21913
rect 12412 -22055 12428 -22021
rect 12462 -22055 12478 -22021
rect 12292 -22141 12299 -22105
rect 12333 -22141 12337 -22105
rect 12292 -22175 12337 -22141
rect 12292 -22211 12299 -22175
rect 12333 -22211 12337 -22175
rect 12292 -22246 12337 -22211
rect 12292 -22282 12299 -22246
rect 12333 -22282 12337 -22246
rect 12154 -22365 12170 -22331
rect 12204 -22365 12220 -22331
rect 12154 -22473 12170 -22439
rect 12204 -22473 12220 -22439
rect 12035 -22559 12041 -22523
rect 12075 -22559 12080 -22523
rect 12035 -22593 12080 -22559
rect 12035 -22629 12041 -22593
rect 12075 -22629 12080 -22593
rect 12035 -22663 12080 -22629
rect 12035 -22699 12041 -22663
rect 12075 -22699 12080 -22663
rect 11896 -22783 11912 -22749
rect 11946 -22783 11962 -22749
rect 11896 -22891 11912 -22857
rect 11946 -22891 11962 -22857
rect 11777 -22977 11783 -22941
rect 11817 -22977 11822 -22941
rect 11777 -23011 11822 -22977
rect 11777 -23047 11783 -23011
rect 11817 -23047 11822 -23011
rect 11777 -23081 11822 -23047
rect 11777 -23117 11783 -23081
rect 11817 -23117 11822 -23081
rect 11777 -23359 11822 -23117
rect 12035 -22941 12080 -22699
rect 12292 -22523 12337 -22282
rect 12552 -22105 12597 -21863
rect 12810 -21687 12855 -21445
rect 13067 -21269 13112 -21225
rect 13067 -21305 13073 -21269
rect 13107 -21305 13112 -21269
rect 13067 -21339 13112 -21305
rect 13067 -21375 13073 -21339
rect 13107 -21375 13112 -21339
rect 13067 -21409 13112 -21375
rect 13067 -21445 13073 -21409
rect 13107 -21445 13112 -21409
rect 12928 -21529 12944 -21495
rect 12978 -21529 12994 -21495
rect 12928 -21637 12944 -21603
rect 12978 -21637 12994 -21603
rect 12810 -21723 12815 -21687
rect 12849 -21723 12855 -21687
rect 12810 -21757 12855 -21723
rect 12810 -21793 12815 -21757
rect 12849 -21793 12855 -21757
rect 12810 -21827 12855 -21793
rect 12810 -21863 12815 -21827
rect 12849 -21863 12855 -21827
rect 12670 -21947 12686 -21913
rect 12720 -21947 12736 -21913
rect 12670 -22055 12686 -22021
rect 12720 -22055 12736 -22021
rect 12552 -22141 12557 -22105
rect 12591 -22141 12597 -22105
rect 12552 -22175 12597 -22141
rect 12552 -22211 12557 -22175
rect 12591 -22211 12597 -22175
rect 12552 -22245 12597 -22211
rect 12552 -22281 12557 -22245
rect 12591 -22281 12597 -22245
rect 12412 -22365 12428 -22331
rect 12462 -22365 12478 -22331
rect 12412 -22473 12428 -22439
rect 12462 -22473 12478 -22439
rect 12292 -22559 12299 -22523
rect 12333 -22559 12337 -22523
rect 12292 -22593 12337 -22559
rect 12292 -22629 12299 -22593
rect 12333 -22629 12337 -22593
rect 12292 -22664 12337 -22629
rect 12292 -22700 12299 -22664
rect 12333 -22700 12337 -22664
rect 12154 -22783 12170 -22749
rect 12204 -22783 12220 -22749
rect 12154 -22891 12170 -22857
rect 12204 -22891 12220 -22857
rect 12035 -22977 12041 -22941
rect 12075 -22977 12080 -22941
rect 12035 -23011 12080 -22977
rect 12035 -23047 12041 -23011
rect 12075 -23047 12080 -23011
rect 12035 -23081 12080 -23047
rect 12035 -23117 12041 -23081
rect 12075 -23117 12080 -23081
rect 11896 -23201 11912 -23167
rect 11946 -23201 11962 -23167
rect 11896 -23309 11912 -23275
rect 11946 -23309 11962 -23275
rect 11777 -23395 11783 -23359
rect 11817 -23395 11822 -23359
rect 11777 -23429 11822 -23395
rect 11777 -23465 11783 -23429
rect 11817 -23465 11822 -23429
rect 11777 -23499 11822 -23465
rect 11777 -23535 11783 -23499
rect 11817 -23535 11822 -23499
rect 11777 -23777 11822 -23535
rect 12035 -23359 12080 -23117
rect 12292 -22941 12337 -22700
rect 12552 -22523 12597 -22281
rect 12810 -22105 12855 -21863
rect 13067 -21687 13112 -21445
rect 13324 -21269 13369 -21225
rect 13324 -21305 13331 -21269
rect 13365 -21305 13369 -21269
rect 13324 -21339 13369 -21305
rect 13324 -21375 13331 -21339
rect 13365 -21375 13369 -21339
rect 13324 -21409 13369 -21375
rect 13324 -21445 13331 -21409
rect 13365 -21445 13369 -21409
rect 13186 -21529 13202 -21495
rect 13236 -21529 13252 -21495
rect 13186 -21637 13202 -21603
rect 13236 -21637 13252 -21603
rect 13067 -21723 13073 -21687
rect 13107 -21723 13112 -21687
rect 13067 -21757 13112 -21723
rect 13067 -21793 13073 -21757
rect 13107 -21793 13112 -21757
rect 13067 -21827 13112 -21793
rect 13067 -21863 13073 -21827
rect 13107 -21863 13112 -21827
rect 12928 -21947 12944 -21913
rect 12978 -21947 12994 -21913
rect 12928 -22055 12944 -22021
rect 12978 -22055 12994 -22021
rect 12810 -22141 12815 -22105
rect 12849 -22141 12855 -22105
rect 12810 -22175 12855 -22141
rect 12810 -22211 12815 -22175
rect 12849 -22211 12855 -22175
rect 12810 -22245 12855 -22211
rect 12810 -22281 12815 -22245
rect 12849 -22281 12855 -22245
rect 12670 -22365 12686 -22331
rect 12720 -22365 12736 -22331
rect 12670 -22473 12686 -22439
rect 12720 -22473 12736 -22439
rect 12552 -22559 12557 -22523
rect 12591 -22559 12597 -22523
rect 12552 -22593 12597 -22559
rect 12552 -22629 12557 -22593
rect 12591 -22629 12597 -22593
rect 12552 -22663 12597 -22629
rect 12552 -22699 12557 -22663
rect 12591 -22699 12597 -22663
rect 12412 -22783 12428 -22749
rect 12462 -22783 12478 -22749
rect 12412 -22891 12428 -22857
rect 12462 -22891 12478 -22857
rect 12292 -22977 12299 -22941
rect 12333 -22977 12337 -22941
rect 12292 -23011 12337 -22977
rect 12292 -23047 12299 -23011
rect 12333 -23047 12337 -23011
rect 12292 -23082 12337 -23047
rect 12292 -23118 12299 -23082
rect 12333 -23118 12337 -23082
rect 12154 -23201 12170 -23167
rect 12204 -23201 12220 -23167
rect 12154 -23309 12170 -23275
rect 12204 -23309 12220 -23275
rect 12035 -23395 12041 -23359
rect 12075 -23395 12080 -23359
rect 12035 -23429 12080 -23395
rect 12035 -23465 12041 -23429
rect 12075 -23465 12080 -23429
rect 12035 -23499 12080 -23465
rect 12035 -23535 12041 -23499
rect 12075 -23535 12080 -23499
rect 11896 -23619 11912 -23585
rect 11946 -23619 11962 -23585
rect 11896 -23727 11912 -23693
rect 11946 -23727 11962 -23693
rect 11777 -23813 11783 -23777
rect 11817 -23813 11822 -23777
rect 11777 -23847 11822 -23813
rect 11777 -23883 11783 -23847
rect 11817 -23883 11822 -23847
rect 11777 -23917 11822 -23883
rect 11777 -23953 11783 -23917
rect 11817 -23953 11822 -23917
rect 11777 -24195 11822 -23953
rect 12035 -23777 12080 -23535
rect 12292 -23359 12337 -23118
rect 12552 -22941 12597 -22699
rect 12810 -22523 12855 -22281
rect 13067 -22105 13112 -21863
rect 13324 -21687 13369 -21445
rect 13583 -21269 13628 -21225
rect 13583 -21305 13589 -21269
rect 13623 -21305 13628 -21269
rect 13583 -21339 13628 -21305
rect 13583 -21375 13589 -21339
rect 13623 -21375 13628 -21339
rect 13583 -21409 13628 -21375
rect 13583 -21445 13589 -21409
rect 13623 -21445 13628 -21409
rect 13444 -21529 13460 -21495
rect 13494 -21529 13510 -21495
rect 13444 -21637 13460 -21603
rect 13494 -21637 13510 -21603
rect 13324 -21723 13331 -21687
rect 13365 -21723 13369 -21687
rect 13324 -21757 13369 -21723
rect 13324 -21793 13331 -21757
rect 13365 -21793 13369 -21757
rect 13324 -21827 13369 -21793
rect 13324 -21863 13331 -21827
rect 13365 -21863 13369 -21827
rect 13186 -21947 13202 -21913
rect 13236 -21947 13252 -21913
rect 13186 -22055 13202 -22021
rect 13236 -22055 13252 -22021
rect 13067 -22141 13073 -22105
rect 13107 -22141 13112 -22105
rect 13067 -22175 13112 -22141
rect 13067 -22211 13073 -22175
rect 13107 -22211 13112 -22175
rect 13067 -22245 13112 -22211
rect 13067 -22281 13073 -22245
rect 13107 -22281 13112 -22245
rect 12928 -22365 12944 -22331
rect 12978 -22365 12994 -22331
rect 12928 -22473 12944 -22439
rect 12978 -22473 12994 -22439
rect 12810 -22559 12815 -22523
rect 12849 -22559 12855 -22523
rect 12810 -22593 12855 -22559
rect 12810 -22629 12815 -22593
rect 12849 -22629 12855 -22593
rect 12810 -22663 12855 -22629
rect 12810 -22699 12815 -22663
rect 12849 -22699 12855 -22663
rect 12670 -22783 12686 -22749
rect 12720 -22783 12736 -22749
rect 12670 -22891 12686 -22857
rect 12720 -22891 12736 -22857
rect 12552 -22977 12557 -22941
rect 12591 -22977 12597 -22941
rect 12552 -23011 12597 -22977
rect 12552 -23047 12557 -23011
rect 12591 -23047 12597 -23011
rect 12552 -23081 12597 -23047
rect 12552 -23117 12557 -23081
rect 12591 -23117 12597 -23081
rect 12412 -23201 12428 -23167
rect 12462 -23201 12478 -23167
rect 12412 -23309 12428 -23275
rect 12462 -23309 12478 -23275
rect 12292 -23395 12299 -23359
rect 12333 -23395 12337 -23359
rect 12292 -23429 12337 -23395
rect 12292 -23465 12299 -23429
rect 12333 -23465 12337 -23429
rect 12292 -23500 12337 -23465
rect 12292 -23536 12299 -23500
rect 12333 -23536 12337 -23500
rect 12154 -23619 12170 -23585
rect 12204 -23619 12220 -23585
rect 12154 -23727 12170 -23693
rect 12204 -23727 12220 -23693
rect 12035 -23813 12041 -23777
rect 12075 -23813 12080 -23777
rect 12035 -23847 12080 -23813
rect 12035 -23883 12041 -23847
rect 12075 -23883 12080 -23847
rect 12035 -23917 12080 -23883
rect 12035 -23953 12041 -23917
rect 12075 -23953 12080 -23917
rect 11896 -24037 11912 -24003
rect 11946 -24037 11962 -24003
rect 12035 -24071 12080 -23953
rect 12292 -23777 12337 -23536
rect 12552 -23359 12597 -23117
rect 12810 -22941 12855 -22699
rect 13067 -22523 13112 -22281
rect 13324 -22105 13369 -21863
rect 13583 -21687 13628 -21445
rect 13841 -21269 13886 -21083
rect 16500 -21084 16549 -21082
rect 14559 -21218 14575 -21184
rect 14609 -21218 14625 -21184
rect 14817 -21218 14833 -21184
rect 14867 -21218 14883 -21184
rect 15075 -21218 15091 -21184
rect 15125 -21218 15141 -21184
rect 15333 -21218 15349 -21184
rect 15383 -21218 15399 -21184
rect 15591 -21218 15607 -21184
rect 15641 -21218 15657 -21184
rect 15849 -21218 15865 -21184
rect 15899 -21218 15915 -21184
rect 16107 -21218 16123 -21184
rect 16157 -21218 16173 -21184
rect 16365 -21218 16381 -21184
rect 16415 -21218 16431 -21184
rect 13841 -21305 13847 -21269
rect 13881 -21305 13886 -21269
rect 13841 -21339 13886 -21305
rect 13841 -21375 13847 -21339
rect 13881 -21375 13886 -21339
rect 13841 -21409 13886 -21375
rect 13841 -21445 13847 -21409
rect 13881 -21445 13886 -21409
rect 13702 -21529 13718 -21495
rect 13752 -21529 13768 -21495
rect 13702 -21637 13718 -21603
rect 13752 -21637 13768 -21603
rect 13583 -21723 13589 -21687
rect 13623 -21723 13628 -21687
rect 13583 -21757 13628 -21723
rect 13583 -21793 13589 -21757
rect 13623 -21793 13628 -21757
rect 13583 -21827 13628 -21793
rect 13583 -21863 13589 -21827
rect 13623 -21863 13628 -21827
rect 13444 -21947 13460 -21913
rect 13494 -21947 13510 -21913
rect 13444 -22055 13460 -22021
rect 13494 -22055 13510 -22021
rect 13324 -22141 13331 -22105
rect 13365 -22141 13369 -22105
rect 13324 -22175 13369 -22141
rect 13324 -22211 13331 -22175
rect 13365 -22211 13369 -22175
rect 13324 -22245 13369 -22211
rect 13324 -22281 13331 -22245
rect 13365 -22281 13369 -22245
rect 13186 -22365 13202 -22331
rect 13236 -22365 13252 -22331
rect 13186 -22473 13202 -22439
rect 13236 -22473 13252 -22439
rect 13067 -22559 13073 -22523
rect 13107 -22559 13112 -22523
rect 13067 -22593 13112 -22559
rect 13067 -22629 13073 -22593
rect 13107 -22629 13112 -22593
rect 13067 -22663 13112 -22629
rect 13067 -22699 13073 -22663
rect 13107 -22699 13112 -22663
rect 12928 -22783 12944 -22749
rect 12978 -22783 12994 -22749
rect 12928 -22891 12944 -22857
rect 12978 -22891 12994 -22857
rect 12810 -22977 12815 -22941
rect 12849 -22977 12855 -22941
rect 12810 -23011 12855 -22977
rect 12810 -23047 12815 -23011
rect 12849 -23047 12855 -23011
rect 12810 -23081 12855 -23047
rect 12810 -23117 12815 -23081
rect 12849 -23117 12855 -23081
rect 12670 -23201 12686 -23167
rect 12720 -23201 12736 -23167
rect 12670 -23309 12686 -23275
rect 12720 -23309 12736 -23275
rect 12552 -23395 12557 -23359
rect 12591 -23395 12597 -23359
rect 12552 -23429 12597 -23395
rect 12552 -23465 12557 -23429
rect 12591 -23465 12597 -23429
rect 12552 -23499 12597 -23465
rect 12552 -23535 12557 -23499
rect 12591 -23535 12597 -23499
rect 12412 -23619 12428 -23585
rect 12462 -23619 12478 -23585
rect 12412 -23727 12428 -23693
rect 12462 -23727 12478 -23693
rect 12292 -23813 12299 -23777
rect 12333 -23813 12337 -23777
rect 12292 -23847 12337 -23813
rect 12292 -23883 12299 -23847
rect 12333 -23883 12337 -23847
rect 12292 -23918 12337 -23883
rect 12292 -23954 12299 -23918
rect 12333 -23954 12337 -23918
rect 12154 -24037 12170 -24003
rect 12204 -24037 12220 -24003
rect 12292 -24071 12337 -23954
rect 12552 -23777 12597 -23535
rect 12810 -23359 12855 -23117
rect 13067 -22941 13112 -22699
rect 13324 -22523 13369 -22281
rect 13583 -22105 13628 -21863
rect 13841 -21687 13886 -21445
rect 13841 -21723 13847 -21687
rect 13881 -21723 13886 -21687
rect 13841 -21757 13886 -21723
rect 13841 -21793 13847 -21757
rect 13881 -21793 13886 -21757
rect 13841 -21827 13886 -21793
rect 13841 -21863 13847 -21827
rect 13881 -21863 13886 -21827
rect 13702 -21947 13718 -21913
rect 13752 -21947 13768 -21913
rect 13702 -22055 13718 -22021
rect 13752 -22055 13768 -22021
rect 13583 -22141 13589 -22105
rect 13623 -22141 13628 -22105
rect 13583 -22175 13628 -22141
rect 13583 -22211 13589 -22175
rect 13623 -22211 13628 -22175
rect 13583 -22245 13628 -22211
rect 13583 -22281 13589 -22245
rect 13623 -22281 13628 -22245
rect 13444 -22365 13460 -22331
rect 13494 -22365 13510 -22331
rect 13444 -22473 13460 -22439
rect 13494 -22473 13510 -22439
rect 13324 -22559 13331 -22523
rect 13365 -22559 13369 -22523
rect 13324 -22593 13369 -22559
rect 13324 -22629 13331 -22593
rect 13365 -22629 13369 -22593
rect 13324 -22663 13369 -22629
rect 13324 -22699 13331 -22663
rect 13365 -22699 13369 -22663
rect 13186 -22783 13202 -22749
rect 13236 -22783 13252 -22749
rect 13186 -22891 13202 -22857
rect 13236 -22891 13252 -22857
rect 13067 -22977 13073 -22941
rect 13107 -22977 13112 -22941
rect 13067 -23011 13112 -22977
rect 13067 -23047 13073 -23011
rect 13107 -23047 13112 -23011
rect 13067 -23081 13112 -23047
rect 13067 -23117 13073 -23081
rect 13107 -23117 13112 -23081
rect 12928 -23201 12944 -23167
rect 12978 -23201 12994 -23167
rect 12928 -23309 12944 -23275
rect 12978 -23309 12994 -23275
rect 12810 -23395 12815 -23359
rect 12849 -23395 12855 -23359
rect 12810 -23429 12855 -23395
rect 12810 -23465 12815 -23429
rect 12849 -23465 12855 -23429
rect 12810 -23499 12855 -23465
rect 12810 -23535 12815 -23499
rect 12849 -23535 12855 -23499
rect 12670 -23619 12686 -23585
rect 12720 -23619 12736 -23585
rect 12670 -23727 12686 -23693
rect 12720 -23727 12736 -23693
rect 12552 -23813 12557 -23777
rect 12591 -23813 12597 -23777
rect 12552 -23847 12597 -23813
rect 12552 -23883 12557 -23847
rect 12591 -23883 12597 -23847
rect 12552 -23917 12597 -23883
rect 12552 -23953 12557 -23917
rect 12591 -23953 12597 -23917
rect 12412 -24037 12428 -24003
rect 12462 -24037 12478 -24003
rect 12552 -24071 12597 -23953
rect 12810 -23777 12855 -23535
rect 13067 -23359 13112 -23117
rect 13324 -22941 13369 -22699
rect 13583 -22523 13628 -22281
rect 13841 -22105 13886 -21863
rect 13841 -22141 13847 -22105
rect 13881 -22141 13886 -22105
rect 13841 -22175 13886 -22141
rect 13841 -22211 13847 -22175
rect 13881 -22211 13886 -22175
rect 13841 -22245 13886 -22211
rect 13841 -22281 13847 -22245
rect 13881 -22281 13886 -22245
rect 13702 -22365 13718 -22331
rect 13752 -22365 13768 -22331
rect 13702 -22473 13718 -22439
rect 13752 -22473 13768 -22439
rect 13583 -22559 13589 -22523
rect 13623 -22559 13628 -22523
rect 13583 -22593 13628 -22559
rect 13583 -22629 13589 -22593
rect 13623 -22629 13628 -22593
rect 13583 -22663 13628 -22629
rect 13583 -22699 13589 -22663
rect 13623 -22699 13628 -22663
rect 13444 -22783 13460 -22749
rect 13494 -22783 13510 -22749
rect 13444 -22891 13460 -22857
rect 13494 -22891 13510 -22857
rect 13324 -22977 13331 -22941
rect 13365 -22977 13369 -22941
rect 13324 -23011 13369 -22977
rect 13324 -23047 13331 -23011
rect 13365 -23047 13369 -23011
rect 13324 -23081 13369 -23047
rect 13324 -23117 13331 -23081
rect 13365 -23117 13369 -23081
rect 13186 -23201 13202 -23167
rect 13236 -23201 13252 -23167
rect 13186 -23309 13202 -23275
rect 13236 -23309 13252 -23275
rect 13067 -23395 13073 -23359
rect 13107 -23395 13112 -23359
rect 13067 -23429 13112 -23395
rect 13067 -23465 13073 -23429
rect 13107 -23465 13112 -23429
rect 13067 -23499 13112 -23465
rect 13067 -23535 13073 -23499
rect 13107 -23535 13112 -23499
rect 12928 -23619 12944 -23585
rect 12978 -23619 12994 -23585
rect 12928 -23727 12944 -23693
rect 12978 -23727 12994 -23693
rect 12810 -23813 12815 -23777
rect 12849 -23813 12855 -23777
rect 12810 -23847 12855 -23813
rect 12810 -23883 12815 -23847
rect 12849 -23883 12855 -23847
rect 12810 -23917 12855 -23883
rect 12810 -23953 12815 -23917
rect 12849 -23953 12855 -23917
rect 12670 -24037 12686 -24003
rect 12720 -24037 12736 -24003
rect 12810 -24071 12855 -23953
rect 13067 -23777 13112 -23535
rect 13324 -23359 13369 -23117
rect 13583 -22941 13628 -22699
rect 13841 -22523 13886 -22281
rect 13841 -22559 13847 -22523
rect 13881 -22559 13886 -22523
rect 13841 -22593 13886 -22559
rect 13841 -22629 13847 -22593
rect 13881 -22629 13886 -22593
rect 13841 -22663 13886 -22629
rect 13841 -22699 13847 -22663
rect 13881 -22699 13886 -22663
rect 13702 -22783 13718 -22749
rect 13752 -22783 13768 -22749
rect 13702 -22891 13718 -22857
rect 13752 -22891 13768 -22857
rect 13583 -22977 13589 -22941
rect 13623 -22977 13628 -22941
rect 13583 -23011 13628 -22977
rect 13583 -23047 13589 -23011
rect 13623 -23047 13628 -23011
rect 13583 -23081 13628 -23047
rect 13583 -23117 13589 -23081
rect 13623 -23117 13628 -23081
rect 13444 -23201 13460 -23167
rect 13494 -23201 13510 -23167
rect 13444 -23309 13460 -23275
rect 13494 -23309 13510 -23275
rect 13324 -23395 13331 -23359
rect 13365 -23395 13369 -23359
rect 13324 -23429 13369 -23395
rect 13324 -23465 13331 -23429
rect 13365 -23465 13369 -23429
rect 13324 -23499 13369 -23465
rect 13324 -23535 13331 -23499
rect 13365 -23535 13369 -23499
rect 13186 -23619 13202 -23585
rect 13236 -23619 13252 -23585
rect 13186 -23727 13202 -23693
rect 13236 -23727 13252 -23693
rect 13067 -23813 13073 -23777
rect 13107 -23813 13112 -23777
rect 13067 -23847 13112 -23813
rect 13067 -23883 13073 -23847
rect 13107 -23883 13112 -23847
rect 13067 -23917 13112 -23883
rect 13067 -23953 13073 -23917
rect 13107 -23953 13112 -23917
rect 12928 -24037 12944 -24003
rect 12978 -24037 12994 -24003
rect 13067 -24071 13112 -23953
rect 13324 -23777 13369 -23535
rect 13583 -23359 13628 -23117
rect 13841 -22941 13886 -22699
rect 13841 -22977 13847 -22941
rect 13881 -22977 13886 -22941
rect 13841 -23011 13886 -22977
rect 13841 -23047 13847 -23011
rect 13881 -23047 13886 -23011
rect 13841 -23081 13886 -23047
rect 13841 -23117 13847 -23081
rect 13881 -23117 13886 -23081
rect 13702 -23201 13718 -23167
rect 13752 -23201 13768 -23167
rect 13702 -23309 13718 -23275
rect 13752 -23309 13768 -23275
rect 13583 -23395 13589 -23359
rect 13623 -23395 13628 -23359
rect 13583 -23429 13628 -23395
rect 13583 -23465 13589 -23429
rect 13623 -23465 13628 -23429
rect 13583 -23499 13628 -23465
rect 13583 -23535 13589 -23499
rect 13623 -23535 13628 -23499
rect 13444 -23619 13460 -23585
rect 13494 -23619 13510 -23585
rect 13444 -23727 13460 -23693
rect 13494 -23727 13510 -23693
rect 13324 -23813 13331 -23777
rect 13365 -23813 13369 -23777
rect 13324 -23847 13369 -23813
rect 13324 -23883 13331 -23847
rect 13365 -23883 13369 -23847
rect 13324 -23917 13369 -23883
rect 13324 -23953 13331 -23917
rect 13365 -23953 13369 -23917
rect 13186 -24037 13202 -24003
rect 13236 -24037 13252 -24003
rect 13324 -24071 13369 -23953
rect 13583 -23777 13628 -23535
rect 13841 -23359 13886 -23117
rect 13841 -23395 13847 -23359
rect 13881 -23395 13886 -23359
rect 13841 -23429 13886 -23395
rect 13841 -23465 13847 -23429
rect 13881 -23465 13886 -23429
rect 13841 -23499 13886 -23465
rect 13841 -23535 13847 -23499
rect 13881 -23535 13886 -23499
rect 13702 -23619 13718 -23585
rect 13752 -23619 13768 -23585
rect 13702 -23727 13718 -23693
rect 13752 -23727 13768 -23693
rect 13583 -23813 13589 -23777
rect 13623 -23813 13628 -23777
rect 13583 -23847 13628 -23813
rect 13583 -23883 13589 -23847
rect 13623 -23883 13628 -23847
rect 13583 -23917 13628 -23883
rect 13583 -23953 13589 -23917
rect 13623 -23953 13628 -23917
rect 13444 -24037 13460 -24003
rect 13494 -24037 13510 -24003
rect 13583 -24071 13628 -23953
rect 13841 -23777 13886 -23535
rect 13841 -23813 13847 -23777
rect 13881 -23813 13886 -23777
rect 13841 -23847 13886 -23813
rect 13841 -23883 13847 -23847
rect 13881 -23883 13886 -23847
rect 13841 -23917 13886 -23883
rect 13841 -23953 13847 -23917
rect 13881 -23953 13886 -23917
rect 13702 -24037 13718 -24003
rect 13752 -24037 13768 -24003
rect 13841 -24071 13886 -23953
rect 14440 -21268 14485 -21224
rect 14440 -21304 14446 -21268
rect 14480 -21304 14485 -21268
rect 14440 -21338 14485 -21304
rect 14440 -21374 14446 -21338
rect 14480 -21374 14485 -21338
rect 14440 -21408 14485 -21374
rect 14440 -21444 14446 -21408
rect 14480 -21444 14485 -21408
rect 14440 -21686 14485 -21444
rect 14698 -21268 14743 -21224
rect 14698 -21304 14704 -21268
rect 14738 -21304 14743 -21268
rect 14698 -21338 14743 -21304
rect 14698 -21374 14704 -21338
rect 14738 -21374 14743 -21338
rect 14698 -21408 14743 -21374
rect 14698 -21444 14704 -21408
rect 14738 -21444 14743 -21408
rect 14559 -21528 14575 -21494
rect 14609 -21528 14625 -21494
rect 14559 -21636 14575 -21602
rect 14609 -21636 14625 -21602
rect 14440 -21722 14446 -21686
rect 14480 -21722 14485 -21686
rect 14440 -21756 14485 -21722
rect 14440 -21792 14446 -21756
rect 14480 -21792 14485 -21756
rect 14440 -21826 14485 -21792
rect 14440 -21862 14446 -21826
rect 14480 -21862 14485 -21826
rect 14440 -22104 14485 -21862
rect 14698 -21686 14743 -21444
rect 14955 -21268 15000 -21224
rect 14955 -21304 14962 -21268
rect 14996 -21304 15000 -21268
rect 14955 -21338 15000 -21304
rect 14955 -21374 14962 -21338
rect 14996 -21374 15000 -21338
rect 14955 -21409 15000 -21374
rect 14955 -21445 14962 -21409
rect 14996 -21445 15000 -21409
rect 14817 -21528 14833 -21494
rect 14867 -21528 14883 -21494
rect 14817 -21636 14833 -21602
rect 14867 -21636 14883 -21602
rect 14698 -21722 14704 -21686
rect 14738 -21722 14743 -21686
rect 14698 -21756 14743 -21722
rect 14698 -21792 14704 -21756
rect 14738 -21792 14743 -21756
rect 14698 -21826 14743 -21792
rect 14698 -21862 14704 -21826
rect 14738 -21862 14743 -21826
rect 14559 -21946 14575 -21912
rect 14609 -21946 14625 -21912
rect 14559 -22054 14575 -22020
rect 14609 -22054 14625 -22020
rect 14440 -22140 14446 -22104
rect 14480 -22140 14485 -22104
rect 14440 -22174 14485 -22140
rect 14440 -22210 14446 -22174
rect 14480 -22210 14485 -22174
rect 14440 -22244 14485 -22210
rect 14440 -22280 14446 -22244
rect 14480 -22280 14485 -22244
rect 14440 -22522 14485 -22280
rect 14698 -22104 14743 -21862
rect 14955 -21686 15000 -21445
rect 15215 -21268 15260 -21224
rect 15215 -21304 15220 -21268
rect 15254 -21304 15260 -21268
rect 15215 -21338 15260 -21304
rect 15215 -21374 15220 -21338
rect 15254 -21374 15260 -21338
rect 15215 -21408 15260 -21374
rect 15215 -21444 15220 -21408
rect 15254 -21444 15260 -21408
rect 15075 -21528 15091 -21494
rect 15125 -21528 15141 -21494
rect 15075 -21636 15091 -21602
rect 15125 -21636 15141 -21602
rect 14955 -21722 14962 -21686
rect 14996 -21722 15000 -21686
rect 14955 -21756 15000 -21722
rect 14955 -21792 14962 -21756
rect 14996 -21792 15000 -21756
rect 14955 -21827 15000 -21792
rect 14955 -21863 14962 -21827
rect 14996 -21863 15000 -21827
rect 14817 -21946 14833 -21912
rect 14867 -21946 14883 -21912
rect 14817 -22054 14833 -22020
rect 14867 -22054 14883 -22020
rect 14698 -22140 14704 -22104
rect 14738 -22140 14743 -22104
rect 14698 -22174 14743 -22140
rect 14698 -22210 14704 -22174
rect 14738 -22210 14743 -22174
rect 14698 -22244 14743 -22210
rect 14698 -22280 14704 -22244
rect 14738 -22280 14743 -22244
rect 14559 -22364 14575 -22330
rect 14609 -22364 14625 -22330
rect 14559 -22472 14575 -22438
rect 14609 -22472 14625 -22438
rect 14440 -22558 14446 -22522
rect 14480 -22558 14485 -22522
rect 14440 -22592 14485 -22558
rect 14440 -22628 14446 -22592
rect 14480 -22628 14485 -22592
rect 14440 -22662 14485 -22628
rect 14440 -22698 14446 -22662
rect 14480 -22698 14485 -22662
rect 14440 -22940 14485 -22698
rect 14698 -22522 14743 -22280
rect 14955 -22104 15000 -21863
rect 15215 -21686 15260 -21444
rect 15473 -21268 15518 -21224
rect 15473 -21304 15478 -21268
rect 15512 -21304 15518 -21268
rect 15473 -21338 15518 -21304
rect 15473 -21374 15478 -21338
rect 15512 -21374 15518 -21338
rect 15473 -21408 15518 -21374
rect 15473 -21444 15478 -21408
rect 15512 -21444 15518 -21408
rect 15333 -21528 15349 -21494
rect 15383 -21528 15399 -21494
rect 15333 -21636 15349 -21602
rect 15383 -21636 15399 -21602
rect 15215 -21722 15220 -21686
rect 15254 -21722 15260 -21686
rect 15215 -21756 15260 -21722
rect 15215 -21792 15220 -21756
rect 15254 -21792 15260 -21756
rect 15215 -21826 15260 -21792
rect 15215 -21862 15220 -21826
rect 15254 -21862 15260 -21826
rect 15075 -21946 15091 -21912
rect 15125 -21946 15141 -21912
rect 15075 -22054 15091 -22020
rect 15125 -22054 15141 -22020
rect 14955 -22140 14962 -22104
rect 14996 -22140 15000 -22104
rect 14955 -22174 15000 -22140
rect 14955 -22210 14962 -22174
rect 14996 -22210 15000 -22174
rect 14955 -22245 15000 -22210
rect 14955 -22281 14962 -22245
rect 14996 -22281 15000 -22245
rect 14817 -22364 14833 -22330
rect 14867 -22364 14883 -22330
rect 14817 -22472 14833 -22438
rect 14867 -22472 14883 -22438
rect 14698 -22558 14704 -22522
rect 14738 -22558 14743 -22522
rect 14698 -22592 14743 -22558
rect 14698 -22628 14704 -22592
rect 14738 -22628 14743 -22592
rect 14698 -22662 14743 -22628
rect 14698 -22698 14704 -22662
rect 14738 -22698 14743 -22662
rect 14559 -22782 14575 -22748
rect 14609 -22782 14625 -22748
rect 14559 -22890 14575 -22856
rect 14609 -22890 14625 -22856
rect 14440 -22976 14446 -22940
rect 14480 -22976 14485 -22940
rect 14440 -23010 14485 -22976
rect 14440 -23046 14446 -23010
rect 14480 -23046 14485 -23010
rect 14440 -23080 14485 -23046
rect 14440 -23116 14446 -23080
rect 14480 -23116 14485 -23080
rect 14440 -23358 14485 -23116
rect 14698 -22940 14743 -22698
rect 14955 -22522 15000 -22281
rect 15215 -22104 15260 -21862
rect 15473 -21686 15518 -21444
rect 15730 -21268 15775 -21224
rect 15730 -21304 15736 -21268
rect 15770 -21304 15775 -21268
rect 15730 -21338 15775 -21304
rect 15730 -21374 15736 -21338
rect 15770 -21374 15775 -21338
rect 15730 -21408 15775 -21374
rect 15730 -21444 15736 -21408
rect 15770 -21444 15775 -21408
rect 15591 -21528 15607 -21494
rect 15641 -21528 15657 -21494
rect 15591 -21636 15607 -21602
rect 15641 -21636 15657 -21602
rect 15473 -21722 15478 -21686
rect 15512 -21722 15518 -21686
rect 15473 -21756 15518 -21722
rect 15473 -21792 15478 -21756
rect 15512 -21792 15518 -21756
rect 15473 -21826 15518 -21792
rect 15473 -21862 15478 -21826
rect 15512 -21862 15518 -21826
rect 15333 -21946 15349 -21912
rect 15383 -21946 15399 -21912
rect 15333 -22054 15349 -22020
rect 15383 -22054 15399 -22020
rect 15215 -22140 15220 -22104
rect 15254 -22140 15260 -22104
rect 15215 -22174 15260 -22140
rect 15215 -22210 15220 -22174
rect 15254 -22210 15260 -22174
rect 15215 -22244 15260 -22210
rect 15215 -22280 15220 -22244
rect 15254 -22280 15260 -22244
rect 15075 -22364 15091 -22330
rect 15125 -22364 15141 -22330
rect 15075 -22472 15091 -22438
rect 15125 -22472 15141 -22438
rect 14955 -22558 14962 -22522
rect 14996 -22558 15000 -22522
rect 14955 -22592 15000 -22558
rect 14955 -22628 14962 -22592
rect 14996 -22628 15000 -22592
rect 14955 -22663 15000 -22628
rect 14955 -22699 14962 -22663
rect 14996 -22699 15000 -22663
rect 14817 -22782 14833 -22748
rect 14867 -22782 14883 -22748
rect 14817 -22890 14833 -22856
rect 14867 -22890 14883 -22856
rect 14698 -22976 14704 -22940
rect 14738 -22976 14743 -22940
rect 14698 -23010 14743 -22976
rect 14698 -23046 14704 -23010
rect 14738 -23046 14743 -23010
rect 14698 -23080 14743 -23046
rect 14698 -23116 14704 -23080
rect 14738 -23116 14743 -23080
rect 14559 -23200 14575 -23166
rect 14609 -23200 14625 -23166
rect 14559 -23308 14575 -23274
rect 14609 -23308 14625 -23274
rect 14440 -23394 14446 -23358
rect 14480 -23394 14485 -23358
rect 14440 -23428 14485 -23394
rect 14440 -23464 14446 -23428
rect 14480 -23464 14485 -23428
rect 14440 -23498 14485 -23464
rect 14440 -23534 14446 -23498
rect 14480 -23534 14485 -23498
rect 14440 -23776 14485 -23534
rect 14698 -23358 14743 -23116
rect 14955 -22940 15000 -22699
rect 15215 -22522 15260 -22280
rect 15473 -22104 15518 -21862
rect 15730 -21686 15775 -21444
rect 15987 -21268 16032 -21224
rect 15987 -21304 15994 -21268
rect 16028 -21304 16032 -21268
rect 15987 -21338 16032 -21304
rect 15987 -21374 15994 -21338
rect 16028 -21374 16032 -21338
rect 15987 -21408 16032 -21374
rect 15987 -21444 15994 -21408
rect 16028 -21444 16032 -21408
rect 15849 -21528 15865 -21494
rect 15899 -21528 15915 -21494
rect 15849 -21636 15865 -21602
rect 15899 -21636 15915 -21602
rect 15730 -21722 15736 -21686
rect 15770 -21722 15775 -21686
rect 15730 -21756 15775 -21722
rect 15730 -21792 15736 -21756
rect 15770 -21792 15775 -21756
rect 15730 -21826 15775 -21792
rect 15730 -21862 15736 -21826
rect 15770 -21862 15775 -21826
rect 15591 -21946 15607 -21912
rect 15641 -21946 15657 -21912
rect 15591 -22054 15607 -22020
rect 15641 -22054 15657 -22020
rect 15473 -22140 15478 -22104
rect 15512 -22140 15518 -22104
rect 15473 -22174 15518 -22140
rect 15473 -22210 15478 -22174
rect 15512 -22210 15518 -22174
rect 15473 -22244 15518 -22210
rect 15473 -22280 15478 -22244
rect 15512 -22280 15518 -22244
rect 15333 -22364 15349 -22330
rect 15383 -22364 15399 -22330
rect 15333 -22472 15349 -22438
rect 15383 -22472 15399 -22438
rect 15215 -22558 15220 -22522
rect 15254 -22558 15260 -22522
rect 15215 -22592 15260 -22558
rect 15215 -22628 15220 -22592
rect 15254 -22628 15260 -22592
rect 15215 -22662 15260 -22628
rect 15215 -22698 15220 -22662
rect 15254 -22698 15260 -22662
rect 15075 -22782 15091 -22748
rect 15125 -22782 15141 -22748
rect 15075 -22890 15091 -22856
rect 15125 -22890 15141 -22856
rect 14955 -22976 14962 -22940
rect 14996 -22976 15000 -22940
rect 14955 -23010 15000 -22976
rect 14955 -23046 14962 -23010
rect 14996 -23046 15000 -23010
rect 14955 -23081 15000 -23046
rect 14955 -23117 14962 -23081
rect 14996 -23117 15000 -23081
rect 14817 -23200 14833 -23166
rect 14867 -23200 14883 -23166
rect 14817 -23308 14833 -23274
rect 14867 -23308 14883 -23274
rect 14698 -23394 14704 -23358
rect 14738 -23394 14743 -23358
rect 14698 -23428 14743 -23394
rect 14698 -23464 14704 -23428
rect 14738 -23464 14743 -23428
rect 14698 -23498 14743 -23464
rect 14698 -23534 14704 -23498
rect 14738 -23534 14743 -23498
rect 14559 -23618 14575 -23584
rect 14609 -23618 14625 -23584
rect 14559 -23726 14575 -23692
rect 14609 -23726 14625 -23692
rect 14440 -23812 14446 -23776
rect 14480 -23812 14485 -23776
rect 14440 -23846 14485 -23812
rect 14440 -23882 14446 -23846
rect 14480 -23882 14485 -23846
rect 14440 -23916 14485 -23882
rect 14440 -23952 14446 -23916
rect 14480 -23952 14485 -23916
rect 14440 -24194 14485 -23952
rect 14698 -23776 14743 -23534
rect 14955 -23358 15000 -23117
rect 15215 -22940 15260 -22698
rect 15473 -22522 15518 -22280
rect 15730 -22104 15775 -21862
rect 15987 -21686 16032 -21444
rect 16246 -21268 16291 -21224
rect 16246 -21304 16252 -21268
rect 16286 -21304 16291 -21268
rect 16246 -21338 16291 -21304
rect 16246 -21374 16252 -21338
rect 16286 -21374 16291 -21338
rect 16246 -21408 16291 -21374
rect 16246 -21444 16252 -21408
rect 16286 -21444 16291 -21408
rect 16107 -21528 16123 -21494
rect 16157 -21528 16173 -21494
rect 16107 -21636 16123 -21602
rect 16157 -21636 16173 -21602
rect 15987 -21722 15994 -21686
rect 16028 -21722 16032 -21686
rect 15987 -21756 16032 -21722
rect 15987 -21792 15994 -21756
rect 16028 -21792 16032 -21756
rect 15987 -21826 16032 -21792
rect 15987 -21862 15994 -21826
rect 16028 -21862 16032 -21826
rect 15849 -21946 15865 -21912
rect 15899 -21946 15915 -21912
rect 15849 -22054 15865 -22020
rect 15899 -22054 15915 -22020
rect 15730 -22140 15736 -22104
rect 15770 -22140 15775 -22104
rect 15730 -22174 15775 -22140
rect 15730 -22210 15736 -22174
rect 15770 -22210 15775 -22174
rect 15730 -22244 15775 -22210
rect 15730 -22280 15736 -22244
rect 15770 -22280 15775 -22244
rect 15591 -22364 15607 -22330
rect 15641 -22364 15657 -22330
rect 15591 -22472 15607 -22438
rect 15641 -22472 15657 -22438
rect 15473 -22558 15478 -22522
rect 15512 -22558 15518 -22522
rect 15473 -22592 15518 -22558
rect 15473 -22628 15478 -22592
rect 15512 -22628 15518 -22592
rect 15473 -22662 15518 -22628
rect 15473 -22698 15478 -22662
rect 15512 -22698 15518 -22662
rect 15333 -22782 15349 -22748
rect 15383 -22782 15399 -22748
rect 15333 -22890 15349 -22856
rect 15383 -22890 15399 -22856
rect 15215 -22976 15220 -22940
rect 15254 -22976 15260 -22940
rect 15215 -23010 15260 -22976
rect 15215 -23046 15220 -23010
rect 15254 -23046 15260 -23010
rect 15215 -23080 15260 -23046
rect 15215 -23116 15220 -23080
rect 15254 -23116 15260 -23080
rect 15075 -23200 15091 -23166
rect 15125 -23200 15141 -23166
rect 15075 -23308 15091 -23274
rect 15125 -23308 15141 -23274
rect 14955 -23394 14962 -23358
rect 14996 -23394 15000 -23358
rect 14955 -23428 15000 -23394
rect 14955 -23464 14962 -23428
rect 14996 -23464 15000 -23428
rect 14955 -23499 15000 -23464
rect 14955 -23535 14962 -23499
rect 14996 -23535 15000 -23499
rect 14817 -23618 14833 -23584
rect 14867 -23618 14883 -23584
rect 14817 -23726 14833 -23692
rect 14867 -23726 14883 -23692
rect 14698 -23812 14704 -23776
rect 14738 -23812 14743 -23776
rect 14698 -23846 14743 -23812
rect 14698 -23882 14704 -23846
rect 14738 -23882 14743 -23846
rect 14698 -23916 14743 -23882
rect 14698 -23952 14704 -23916
rect 14738 -23952 14743 -23916
rect 14559 -24036 14575 -24002
rect 14609 -24036 14625 -24002
rect 14698 -24070 14743 -23952
rect 14955 -23776 15000 -23535
rect 15215 -23358 15260 -23116
rect 15473 -22940 15518 -22698
rect 15730 -22522 15775 -22280
rect 15987 -22104 16032 -21862
rect 16246 -21686 16291 -21444
rect 16504 -21268 16549 -21084
rect 16504 -21304 16510 -21268
rect 16544 -21304 16549 -21268
rect 16504 -21338 16549 -21304
rect 16504 -21374 16510 -21338
rect 16544 -21374 16549 -21338
rect 16504 -21408 16549 -21374
rect 16504 -21444 16510 -21408
rect 16544 -21444 16549 -21408
rect 16365 -21528 16381 -21494
rect 16415 -21528 16431 -21494
rect 16365 -21636 16381 -21602
rect 16415 -21636 16431 -21602
rect 16246 -21722 16252 -21686
rect 16286 -21722 16291 -21686
rect 16246 -21756 16291 -21722
rect 16246 -21792 16252 -21756
rect 16286 -21792 16291 -21756
rect 16246 -21826 16291 -21792
rect 16246 -21862 16252 -21826
rect 16286 -21862 16291 -21826
rect 16107 -21946 16123 -21912
rect 16157 -21946 16173 -21912
rect 16107 -22054 16123 -22020
rect 16157 -22054 16173 -22020
rect 15987 -22140 15994 -22104
rect 16028 -22140 16032 -22104
rect 15987 -22174 16032 -22140
rect 15987 -22210 15994 -22174
rect 16028 -22210 16032 -22174
rect 15987 -22244 16032 -22210
rect 15987 -22280 15994 -22244
rect 16028 -22280 16032 -22244
rect 15849 -22364 15865 -22330
rect 15899 -22364 15915 -22330
rect 15849 -22472 15865 -22438
rect 15899 -22472 15915 -22438
rect 15730 -22558 15736 -22522
rect 15770 -22558 15775 -22522
rect 15730 -22592 15775 -22558
rect 15730 -22628 15736 -22592
rect 15770 -22628 15775 -22592
rect 15730 -22662 15775 -22628
rect 15730 -22698 15736 -22662
rect 15770 -22698 15775 -22662
rect 15591 -22782 15607 -22748
rect 15641 -22782 15657 -22748
rect 15591 -22890 15607 -22856
rect 15641 -22890 15657 -22856
rect 15473 -22976 15478 -22940
rect 15512 -22976 15518 -22940
rect 15473 -23010 15518 -22976
rect 15473 -23046 15478 -23010
rect 15512 -23046 15518 -23010
rect 15473 -23080 15518 -23046
rect 15473 -23116 15478 -23080
rect 15512 -23116 15518 -23080
rect 15333 -23200 15349 -23166
rect 15383 -23200 15399 -23166
rect 15333 -23308 15349 -23274
rect 15383 -23308 15399 -23274
rect 15215 -23394 15220 -23358
rect 15254 -23394 15260 -23358
rect 15215 -23428 15260 -23394
rect 15215 -23464 15220 -23428
rect 15254 -23464 15260 -23428
rect 15215 -23498 15260 -23464
rect 15215 -23534 15220 -23498
rect 15254 -23534 15260 -23498
rect 15075 -23618 15091 -23584
rect 15125 -23618 15141 -23584
rect 15075 -23726 15091 -23692
rect 15125 -23726 15141 -23692
rect 14955 -23812 14962 -23776
rect 14996 -23812 15000 -23776
rect 14955 -23846 15000 -23812
rect 14955 -23882 14962 -23846
rect 14996 -23882 15000 -23846
rect 14955 -23917 15000 -23882
rect 14955 -23953 14962 -23917
rect 14996 -23953 15000 -23917
rect 14817 -24036 14833 -24002
rect 14867 -24036 14883 -24002
rect 14955 -24070 15000 -23953
rect 15215 -23776 15260 -23534
rect 15473 -23358 15518 -23116
rect 15730 -22940 15775 -22698
rect 15987 -22522 16032 -22280
rect 16246 -22104 16291 -21862
rect 16504 -21686 16549 -21444
rect 16504 -21722 16510 -21686
rect 16544 -21722 16549 -21686
rect 16504 -21756 16549 -21722
rect 16504 -21792 16510 -21756
rect 16544 -21792 16549 -21756
rect 16504 -21826 16549 -21792
rect 16504 -21862 16510 -21826
rect 16544 -21862 16549 -21826
rect 16365 -21946 16381 -21912
rect 16415 -21946 16431 -21912
rect 16365 -22054 16381 -22020
rect 16415 -22054 16431 -22020
rect 16246 -22140 16252 -22104
rect 16286 -22140 16291 -22104
rect 16246 -22174 16291 -22140
rect 16246 -22210 16252 -22174
rect 16286 -22210 16291 -22174
rect 16246 -22244 16291 -22210
rect 16246 -22280 16252 -22244
rect 16286 -22280 16291 -22244
rect 16107 -22364 16123 -22330
rect 16157 -22364 16173 -22330
rect 16107 -22472 16123 -22438
rect 16157 -22472 16173 -22438
rect 15987 -22558 15994 -22522
rect 16028 -22558 16032 -22522
rect 15987 -22592 16032 -22558
rect 15987 -22628 15994 -22592
rect 16028 -22628 16032 -22592
rect 15987 -22662 16032 -22628
rect 15987 -22698 15994 -22662
rect 16028 -22698 16032 -22662
rect 15849 -22782 15865 -22748
rect 15899 -22782 15915 -22748
rect 15849 -22890 15865 -22856
rect 15899 -22890 15915 -22856
rect 15730 -22976 15736 -22940
rect 15770 -22976 15775 -22940
rect 15730 -23010 15775 -22976
rect 15730 -23046 15736 -23010
rect 15770 -23046 15775 -23010
rect 15730 -23080 15775 -23046
rect 15730 -23116 15736 -23080
rect 15770 -23116 15775 -23080
rect 15591 -23200 15607 -23166
rect 15641 -23200 15657 -23166
rect 15591 -23308 15607 -23274
rect 15641 -23308 15657 -23274
rect 15473 -23394 15478 -23358
rect 15512 -23394 15518 -23358
rect 15473 -23428 15518 -23394
rect 15473 -23464 15478 -23428
rect 15512 -23464 15518 -23428
rect 15473 -23498 15518 -23464
rect 15473 -23534 15478 -23498
rect 15512 -23534 15518 -23498
rect 15333 -23618 15349 -23584
rect 15383 -23618 15399 -23584
rect 15333 -23726 15349 -23692
rect 15383 -23726 15399 -23692
rect 15215 -23812 15220 -23776
rect 15254 -23812 15260 -23776
rect 15215 -23846 15260 -23812
rect 15215 -23882 15220 -23846
rect 15254 -23882 15260 -23846
rect 15215 -23916 15260 -23882
rect 15215 -23952 15220 -23916
rect 15254 -23952 15260 -23916
rect 15075 -24036 15091 -24002
rect 15125 -24036 15141 -24002
rect 15215 -24070 15260 -23952
rect 15473 -23776 15518 -23534
rect 15730 -23358 15775 -23116
rect 15987 -22940 16032 -22698
rect 16246 -22522 16291 -22280
rect 16504 -22104 16549 -21862
rect 16504 -22140 16510 -22104
rect 16544 -22140 16549 -22104
rect 16504 -22174 16549 -22140
rect 16504 -22210 16510 -22174
rect 16544 -22210 16549 -22174
rect 16504 -22244 16549 -22210
rect 16504 -22280 16510 -22244
rect 16544 -22280 16549 -22244
rect 16365 -22364 16381 -22330
rect 16415 -22364 16431 -22330
rect 16365 -22472 16381 -22438
rect 16415 -22472 16431 -22438
rect 16246 -22558 16252 -22522
rect 16286 -22558 16291 -22522
rect 16246 -22592 16291 -22558
rect 16246 -22628 16252 -22592
rect 16286 -22628 16291 -22592
rect 16246 -22662 16291 -22628
rect 16246 -22698 16252 -22662
rect 16286 -22698 16291 -22662
rect 16107 -22782 16123 -22748
rect 16157 -22782 16173 -22748
rect 16107 -22890 16123 -22856
rect 16157 -22890 16173 -22856
rect 15987 -22976 15994 -22940
rect 16028 -22976 16032 -22940
rect 15987 -23010 16032 -22976
rect 15987 -23046 15994 -23010
rect 16028 -23046 16032 -23010
rect 15987 -23080 16032 -23046
rect 15987 -23116 15994 -23080
rect 16028 -23116 16032 -23080
rect 15849 -23200 15865 -23166
rect 15899 -23200 15915 -23166
rect 15849 -23308 15865 -23274
rect 15899 -23308 15915 -23274
rect 15730 -23394 15736 -23358
rect 15770 -23394 15775 -23358
rect 15730 -23428 15775 -23394
rect 15730 -23464 15736 -23428
rect 15770 -23464 15775 -23428
rect 15730 -23498 15775 -23464
rect 15730 -23534 15736 -23498
rect 15770 -23534 15775 -23498
rect 15591 -23618 15607 -23584
rect 15641 -23618 15657 -23584
rect 15591 -23726 15607 -23692
rect 15641 -23726 15657 -23692
rect 15473 -23812 15478 -23776
rect 15512 -23812 15518 -23776
rect 15473 -23846 15518 -23812
rect 15473 -23882 15478 -23846
rect 15512 -23882 15518 -23846
rect 15473 -23916 15518 -23882
rect 15473 -23952 15478 -23916
rect 15512 -23952 15518 -23916
rect 15333 -24036 15349 -24002
rect 15383 -24036 15399 -24002
rect 15473 -24070 15518 -23952
rect 15730 -23776 15775 -23534
rect 15987 -23358 16032 -23116
rect 16246 -22940 16291 -22698
rect 16504 -22522 16549 -22280
rect 16504 -22558 16510 -22522
rect 16544 -22558 16549 -22522
rect 16504 -22592 16549 -22558
rect 16504 -22628 16510 -22592
rect 16544 -22628 16549 -22592
rect 16504 -22662 16549 -22628
rect 16504 -22698 16510 -22662
rect 16544 -22698 16549 -22662
rect 16365 -22782 16381 -22748
rect 16415 -22782 16431 -22748
rect 16365 -22890 16381 -22856
rect 16415 -22890 16431 -22856
rect 16246 -22976 16252 -22940
rect 16286 -22976 16291 -22940
rect 16246 -23010 16291 -22976
rect 16246 -23046 16252 -23010
rect 16286 -23046 16291 -23010
rect 16246 -23080 16291 -23046
rect 16246 -23116 16252 -23080
rect 16286 -23116 16291 -23080
rect 16107 -23200 16123 -23166
rect 16157 -23200 16173 -23166
rect 16107 -23308 16123 -23274
rect 16157 -23308 16173 -23274
rect 15987 -23394 15994 -23358
rect 16028 -23394 16032 -23358
rect 15987 -23428 16032 -23394
rect 15987 -23464 15994 -23428
rect 16028 -23464 16032 -23428
rect 15987 -23498 16032 -23464
rect 15987 -23534 15994 -23498
rect 16028 -23534 16032 -23498
rect 15849 -23618 15865 -23584
rect 15899 -23618 15915 -23584
rect 15849 -23726 15865 -23692
rect 15899 -23726 15915 -23692
rect 15730 -23812 15736 -23776
rect 15770 -23812 15775 -23776
rect 15730 -23846 15775 -23812
rect 15730 -23882 15736 -23846
rect 15770 -23882 15775 -23846
rect 15730 -23916 15775 -23882
rect 15730 -23952 15736 -23916
rect 15770 -23952 15775 -23916
rect 15591 -24036 15607 -24002
rect 15641 -24036 15657 -24002
rect 15730 -24070 15775 -23952
rect 15987 -23776 16032 -23534
rect 16246 -23358 16291 -23116
rect 16504 -22940 16549 -22698
rect 16504 -22976 16510 -22940
rect 16544 -22976 16549 -22940
rect 16504 -23010 16549 -22976
rect 16504 -23046 16510 -23010
rect 16544 -23046 16549 -23010
rect 16504 -23080 16549 -23046
rect 16504 -23116 16510 -23080
rect 16544 -23116 16549 -23080
rect 16365 -23200 16381 -23166
rect 16415 -23200 16431 -23166
rect 16365 -23308 16381 -23274
rect 16415 -23308 16431 -23274
rect 16246 -23394 16252 -23358
rect 16286 -23394 16291 -23358
rect 16246 -23428 16291 -23394
rect 16246 -23464 16252 -23428
rect 16286 -23464 16291 -23428
rect 16246 -23498 16291 -23464
rect 16246 -23534 16252 -23498
rect 16286 -23534 16291 -23498
rect 16107 -23618 16123 -23584
rect 16157 -23618 16173 -23584
rect 16107 -23726 16123 -23692
rect 16157 -23726 16173 -23692
rect 15987 -23812 15994 -23776
rect 16028 -23812 16032 -23776
rect 15987 -23846 16032 -23812
rect 15987 -23882 15994 -23846
rect 16028 -23882 16032 -23846
rect 15987 -23916 16032 -23882
rect 15987 -23952 15994 -23916
rect 16028 -23952 16032 -23916
rect 15849 -24036 15865 -24002
rect 15899 -24036 15915 -24002
rect 15987 -24070 16032 -23952
rect 16246 -23776 16291 -23534
rect 16504 -23358 16549 -23116
rect 16504 -23394 16510 -23358
rect 16544 -23394 16549 -23358
rect 16504 -23428 16549 -23394
rect 16504 -23464 16510 -23428
rect 16544 -23464 16549 -23428
rect 16504 -23498 16549 -23464
rect 16504 -23534 16510 -23498
rect 16544 -23534 16549 -23498
rect 16365 -23618 16381 -23584
rect 16415 -23618 16431 -23584
rect 16365 -23726 16381 -23692
rect 16415 -23726 16431 -23692
rect 16246 -23812 16252 -23776
rect 16286 -23812 16291 -23776
rect 16246 -23846 16291 -23812
rect 16246 -23882 16252 -23846
rect 16286 -23882 16291 -23846
rect 16246 -23916 16291 -23882
rect 16246 -23952 16252 -23916
rect 16286 -23952 16291 -23916
rect 16107 -24036 16123 -24002
rect 16157 -24036 16173 -24002
rect 16246 -24070 16291 -23952
rect 16504 -23776 16549 -23534
rect 16504 -23812 16510 -23776
rect 16544 -23812 16549 -23776
rect 16504 -23846 16549 -23812
rect 16504 -23882 16510 -23846
rect 16544 -23882 16549 -23846
rect 16504 -23916 16549 -23882
rect 16504 -23952 16510 -23916
rect 16544 -23952 16549 -23916
rect 16365 -24036 16381 -24002
rect 16415 -24036 16431 -24002
rect 16504 -24070 16549 -23952
rect 9107 -24290 10333 -24195
rect 11777 -24290 13003 -24195
rect 14440 -24289 15666 -24194
rect 9106 -24379 9122 -24345
rect 9156 -24379 9172 -24345
rect 9646 -24379 9662 -24345
rect 9696 -24379 9712 -24345
rect 10126 -24379 10137 -24345
rect 10187 -24379 10192 -24345
rect 8967 -24431 9029 -24409
rect 8967 -24465 8993 -24431
rect 9027 -24465 9029 -24431
rect 8967 -24499 9029 -24465
rect 8967 -24535 8993 -24499
rect 9027 -24535 9029 -24499
rect 8967 -24569 9029 -24535
rect 8967 -24603 8993 -24569
rect 9027 -24603 9029 -24569
rect 8967 -24645 9029 -24603
rect 9245 -24431 9313 -24411
rect 9245 -24465 9251 -24431
rect 9285 -24465 9313 -24431
rect 9245 -24499 9313 -24465
rect 9245 -24535 9251 -24499
rect 9285 -24535 9313 -24499
rect 9245 -24569 9313 -24535
rect 9245 -24603 9251 -24569
rect 9285 -24603 9313 -24569
rect 9245 -24647 9313 -24603
rect 9507 -24431 9569 -24409
rect 9507 -24465 9533 -24431
rect 9567 -24465 9569 -24431
rect 9507 -24499 9569 -24465
rect 9507 -24535 9533 -24499
rect 9567 -24535 9569 -24499
rect 9507 -24569 9569 -24535
rect 9507 -24603 9533 -24569
rect 9567 -24603 9569 -24569
rect 9507 -24645 9569 -24603
rect 9785 -24431 9853 -24411
rect 9785 -24465 9791 -24431
rect 9825 -24465 9853 -24431
rect 9785 -24499 9853 -24465
rect 9785 -24535 9791 -24499
rect 9825 -24535 9853 -24499
rect 9785 -24569 9853 -24535
rect 9785 -24603 9791 -24569
rect 9825 -24603 9853 -24569
rect 9785 -24647 9853 -24603
rect 9987 -24431 10049 -24409
rect 9987 -24465 10013 -24431
rect 10047 -24465 10049 -24431
rect 9987 -24499 10049 -24465
rect 9987 -24535 10013 -24499
rect 10047 -24535 10049 -24499
rect 9987 -24569 10049 -24535
rect 9987 -24603 10013 -24569
rect 10047 -24603 10049 -24569
rect 9106 -24689 9122 -24655
rect 9156 -24689 9172 -24655
rect 9646 -24689 9662 -24655
rect 9696 -24689 9712 -24655
rect 9987 -24774 10049 -24603
rect 10265 -24431 10333 -24290
rect 10629 -24377 10645 -24343
rect 10679 -24377 10695 -24343
rect 11139 -24367 11155 -24333
rect 11189 -24367 11205 -24333
rect 11776 -24379 11792 -24345
rect 11826 -24379 11842 -24345
rect 12316 -24379 12332 -24345
rect 12366 -24379 12382 -24345
rect 12796 -24379 12807 -24345
rect 12857 -24379 12862 -24345
rect 10265 -24465 10271 -24431
rect 10305 -24465 10333 -24431
rect 10265 -24499 10333 -24465
rect 10265 -24535 10271 -24499
rect 10305 -24535 10333 -24499
rect 10265 -24569 10333 -24535
rect 10265 -24603 10271 -24569
rect 10305 -24603 10333 -24569
rect 10265 -24647 10333 -24603
rect 10490 -24429 10552 -24407
rect 10490 -24463 10516 -24429
rect 10550 -24463 10552 -24429
rect 10490 -24497 10552 -24463
rect 10490 -24533 10516 -24497
rect 10550 -24533 10552 -24497
rect 10490 -24567 10552 -24533
rect 10490 -24601 10516 -24567
rect 10550 -24601 10552 -24567
rect 10490 -24643 10552 -24601
rect 10768 -24429 10836 -24409
rect 10768 -24463 10774 -24429
rect 10808 -24463 10836 -24429
rect 10768 -24497 10836 -24463
rect 10768 -24533 10774 -24497
rect 10808 -24533 10836 -24497
rect 10768 -24567 10836 -24533
rect 10768 -24601 10774 -24567
rect 10808 -24601 10836 -24567
rect 10768 -24645 10836 -24601
rect 11000 -24419 11062 -24397
rect 11000 -24453 11026 -24419
rect 11060 -24453 11062 -24419
rect 11000 -24487 11062 -24453
rect 11000 -24523 11026 -24487
rect 11060 -24523 11062 -24487
rect 11000 -24557 11062 -24523
rect 11000 -24591 11026 -24557
rect 11060 -24591 11062 -24557
rect 11000 -24633 11062 -24591
rect 11278 -24419 11346 -24399
rect 11278 -24453 11284 -24419
rect 11318 -24453 11346 -24419
rect 11278 -24487 11346 -24453
rect 11278 -24523 11284 -24487
rect 11318 -24523 11346 -24487
rect 11278 -24557 11346 -24523
rect 11278 -24591 11284 -24557
rect 11318 -24591 11346 -24557
rect 11278 -24635 11346 -24591
rect 11637 -24431 11699 -24409
rect 11637 -24465 11663 -24431
rect 11697 -24465 11699 -24431
rect 11637 -24499 11699 -24465
rect 11637 -24535 11663 -24499
rect 11697 -24535 11699 -24499
rect 11637 -24569 11699 -24535
rect 11637 -24603 11663 -24569
rect 11697 -24603 11699 -24569
rect 10126 -24689 10138 -24655
rect 10178 -24689 10192 -24655
rect 10629 -24687 10645 -24653
rect 10679 -24687 10695 -24653
rect 11139 -24677 11155 -24643
rect 11189 -24677 11205 -24643
rect 11637 -24645 11699 -24603
rect 11915 -24431 11983 -24411
rect 11915 -24465 11921 -24431
rect 11955 -24465 11983 -24431
rect 11915 -24499 11983 -24465
rect 11915 -24535 11921 -24499
rect 11955 -24535 11983 -24499
rect 11915 -24569 11983 -24535
rect 11915 -24603 11921 -24569
rect 11955 -24603 11983 -24569
rect 11915 -24647 11983 -24603
rect 12177 -24431 12239 -24409
rect 12177 -24465 12203 -24431
rect 12237 -24465 12239 -24431
rect 12177 -24499 12239 -24465
rect 12177 -24535 12203 -24499
rect 12237 -24535 12239 -24499
rect 12177 -24569 12239 -24535
rect 12177 -24603 12203 -24569
rect 12237 -24603 12239 -24569
rect 12177 -24645 12239 -24603
rect 12455 -24431 12523 -24411
rect 12455 -24465 12461 -24431
rect 12495 -24465 12523 -24431
rect 12455 -24499 12523 -24465
rect 12455 -24535 12461 -24499
rect 12495 -24535 12523 -24499
rect 12455 -24569 12523 -24535
rect 12455 -24603 12461 -24569
rect 12495 -24603 12523 -24569
rect 12455 -24647 12523 -24603
rect 12657 -24431 12719 -24409
rect 12657 -24465 12683 -24431
rect 12717 -24465 12719 -24431
rect 12657 -24499 12719 -24465
rect 12657 -24535 12683 -24499
rect 12717 -24535 12719 -24499
rect 12657 -24569 12719 -24535
rect 12657 -24603 12683 -24569
rect 12717 -24603 12719 -24569
rect 11776 -24689 11792 -24655
rect 11826 -24689 11842 -24655
rect 12316 -24689 12332 -24655
rect 12366 -24689 12382 -24655
rect 12657 -24715 12719 -24603
rect 12935 -24431 13003 -24290
rect 13299 -24377 13315 -24343
rect 13349 -24377 13365 -24343
rect 13809 -24367 13825 -24333
rect 13859 -24367 13875 -24333
rect 14439 -24378 14455 -24344
rect 14489 -24378 14505 -24344
rect 14979 -24378 14995 -24344
rect 15029 -24378 15045 -24344
rect 15459 -24378 15470 -24344
rect 15520 -24378 15525 -24344
rect 12935 -24465 12941 -24431
rect 12975 -24465 13003 -24431
rect 12935 -24499 13003 -24465
rect 12935 -24535 12941 -24499
rect 12975 -24535 13003 -24499
rect 12935 -24569 13003 -24535
rect 12935 -24603 12941 -24569
rect 12975 -24603 13003 -24569
rect 12935 -24647 13003 -24603
rect 13160 -24429 13222 -24407
rect 13160 -24463 13186 -24429
rect 13220 -24463 13222 -24429
rect 13160 -24497 13222 -24463
rect 13160 -24533 13186 -24497
rect 13220 -24533 13222 -24497
rect 13160 -24567 13222 -24533
rect 13160 -24601 13186 -24567
rect 13220 -24601 13222 -24567
rect 13160 -24643 13222 -24601
rect 13438 -24429 13506 -24409
rect 13438 -24463 13444 -24429
rect 13478 -24463 13506 -24429
rect 13438 -24497 13506 -24463
rect 13438 -24533 13444 -24497
rect 13478 -24533 13506 -24497
rect 13438 -24567 13506 -24533
rect 13438 -24601 13444 -24567
rect 13478 -24601 13506 -24567
rect 13438 -24645 13506 -24601
rect 13670 -24419 13732 -24397
rect 13670 -24453 13696 -24419
rect 13730 -24453 13732 -24419
rect 13670 -24487 13732 -24453
rect 13670 -24523 13696 -24487
rect 13730 -24523 13732 -24487
rect 13670 -24557 13732 -24523
rect 13670 -24591 13696 -24557
rect 13730 -24591 13732 -24557
rect 13670 -24633 13732 -24591
rect 13948 -24419 14016 -24399
rect 13948 -24453 13954 -24419
rect 13988 -24453 14016 -24419
rect 13948 -24487 14016 -24453
rect 13948 -24523 13954 -24487
rect 13988 -24523 14016 -24487
rect 13948 -24557 14016 -24523
rect 13948 -24591 13954 -24557
rect 13988 -24591 14016 -24557
rect 13948 -24635 14016 -24591
rect 14300 -24430 14362 -24408
rect 14300 -24464 14326 -24430
rect 14360 -24464 14362 -24430
rect 14300 -24498 14362 -24464
rect 14300 -24534 14326 -24498
rect 14360 -24534 14362 -24498
rect 14300 -24568 14362 -24534
rect 14300 -24602 14326 -24568
rect 14360 -24602 14362 -24568
rect 12796 -24689 12808 -24655
rect 12852 -24689 12862 -24655
rect 13299 -24687 13315 -24653
rect 13349 -24687 13365 -24653
rect 13809 -24677 13825 -24643
rect 13859 -24677 13875 -24643
rect 14300 -24644 14362 -24602
rect 14578 -24430 14646 -24410
rect 14578 -24464 14584 -24430
rect 14618 -24464 14646 -24430
rect 14578 -24498 14646 -24464
rect 14578 -24534 14584 -24498
rect 14618 -24534 14646 -24498
rect 14578 -24568 14646 -24534
rect 14578 -24602 14584 -24568
rect 14618 -24602 14646 -24568
rect 14578 -24646 14646 -24602
rect 14840 -24430 14902 -24408
rect 14840 -24464 14866 -24430
rect 14900 -24464 14902 -24430
rect 14840 -24498 14902 -24464
rect 14840 -24534 14866 -24498
rect 14900 -24534 14902 -24498
rect 14840 -24568 14902 -24534
rect 14840 -24602 14866 -24568
rect 14900 -24602 14902 -24568
rect 14840 -24644 14902 -24602
rect 15118 -24430 15186 -24410
rect 15118 -24464 15124 -24430
rect 15158 -24464 15186 -24430
rect 15118 -24498 15186 -24464
rect 15118 -24534 15124 -24498
rect 15158 -24534 15186 -24498
rect 15118 -24568 15186 -24534
rect 15118 -24602 15124 -24568
rect 15158 -24602 15186 -24568
rect 15118 -24646 15186 -24602
rect 15320 -24430 15382 -24408
rect 15320 -24464 15346 -24430
rect 15380 -24464 15382 -24430
rect 15320 -24498 15382 -24464
rect 15320 -24534 15346 -24498
rect 15380 -24534 15382 -24498
rect 15320 -24568 15382 -24534
rect 15320 -24602 15346 -24568
rect 15380 -24602 15382 -24568
rect 14439 -24688 14455 -24654
rect 14489 -24688 14505 -24654
rect 14979 -24688 14995 -24654
rect 15029 -24688 15045 -24654
rect 12656 -24774 12719 -24715
rect 15320 -24774 15382 -24602
rect 15598 -24430 15666 -24289
rect 15962 -24376 15978 -24342
rect 16012 -24376 16028 -24342
rect 16472 -24366 16488 -24332
rect 16522 -24366 16538 -24332
rect 15598 -24464 15604 -24430
rect 15638 -24464 15666 -24430
rect 15598 -24498 15666 -24464
rect 15598 -24534 15604 -24498
rect 15638 -24534 15666 -24498
rect 15598 -24568 15666 -24534
rect 15598 -24602 15604 -24568
rect 15638 -24602 15666 -24568
rect 15598 -24646 15666 -24602
rect 15823 -24428 15885 -24406
rect 15823 -24462 15849 -24428
rect 15883 -24462 15885 -24428
rect 15823 -24496 15885 -24462
rect 15823 -24532 15849 -24496
rect 15883 -24532 15885 -24496
rect 15823 -24566 15885 -24532
rect 15823 -24600 15849 -24566
rect 15883 -24600 15885 -24566
rect 15823 -24642 15885 -24600
rect 16101 -24428 16169 -24408
rect 16101 -24462 16107 -24428
rect 16141 -24462 16169 -24428
rect 16101 -24496 16169 -24462
rect 16101 -24532 16107 -24496
rect 16141 -24532 16169 -24496
rect 16101 -24566 16169 -24532
rect 16101 -24600 16107 -24566
rect 16141 -24600 16169 -24566
rect 16101 -24644 16169 -24600
rect 16333 -24418 16395 -24396
rect 16333 -24452 16359 -24418
rect 16393 -24452 16395 -24418
rect 16333 -24486 16395 -24452
rect 16333 -24522 16359 -24486
rect 16393 -24522 16395 -24486
rect 16333 -24556 16395 -24522
rect 16333 -24590 16359 -24556
rect 16393 -24590 16395 -24556
rect 16333 -24632 16395 -24590
rect 16611 -24418 16679 -24398
rect 16611 -24452 16617 -24418
rect 16651 -24452 16679 -24418
rect 16611 -24486 16679 -24452
rect 16611 -24522 16617 -24486
rect 16651 -24522 16679 -24486
rect 16611 -24556 16679 -24522
rect 16611 -24590 16617 -24556
rect 16651 -24590 16679 -24556
rect 16611 -24634 16679 -24590
rect 15459 -24688 15470 -24654
rect 15514 -24688 15525 -24654
rect 15962 -24686 15978 -24652
rect 16012 -24686 16028 -24652
rect 16472 -24676 16488 -24642
rect 16522 -24676 16538 -24642
rect 8823 -24781 16813 -24774
rect 8820 -24875 9972 -24781
rect 10064 -24875 12642 -24781
rect 12734 -24875 15308 -24781
rect 15400 -24875 16880 -24781
rect 8820 -24969 16880 -24875
rect 18096 -7550 19420 -7505
rect 18036 -7584 18052 -7550
rect 17990 -7634 18024 -7618
rect 17990 -9026 18024 -9010
rect 18096 -9060 19420 -7584
rect 19913 -7550 21244 -7505
rect 21278 -7584 21294 -7550
rect 18036 -9094 18052 -9060
rect 17990 -9144 18024 -9128
rect 17990 -10536 18024 -10520
rect 18096 -10570 19420 -9094
rect 18036 -10604 18052 -10570
rect 17990 -10654 18024 -10638
rect 17990 -12046 18024 -12030
rect 18096 -12080 19420 -10604
rect 18036 -12114 18052 -12080
rect 17990 -12164 18024 -12148
rect 17990 -13556 18024 -13540
rect 18096 -13590 19420 -12114
rect 18036 -13624 18052 -13590
rect 17990 -13674 18024 -13658
rect 17990 -15066 18024 -15050
rect 18096 -15100 19420 -13624
rect 18036 -15134 18052 -15100
rect 17990 -15184 18024 -15168
rect 17990 -16576 18024 -16560
rect 18096 -16610 19420 -15134
rect 18036 -16644 18052 -16610
rect 17990 -16694 18024 -16678
rect 17990 -18086 18024 -18070
rect 18096 -18120 19420 -16644
rect 18036 -18154 18052 -18120
rect 17990 -18204 18024 -18188
rect 17990 -19596 18024 -19580
rect 18096 -19630 19420 -18154
rect 18036 -19664 18052 -19630
rect 17990 -19714 18024 -19698
rect 17990 -21106 18024 -21090
rect 18096 -21140 19420 -19664
rect 18036 -21174 18052 -21140
rect 17990 -21224 18024 -21208
rect 17990 -22616 18024 -22600
rect 18096 -22650 19420 -21174
rect 18036 -22684 18052 -22650
rect 17990 -22734 18024 -22718
rect 17990 -24126 18024 -24110
rect 18096 -24160 19420 -22684
rect 18036 -24194 18052 -24160
rect 17990 -24244 18024 -24228
rect 17990 -25636 18024 -25620
rect 18096 -25670 19420 -24194
rect 18036 -25704 18052 -25670
rect 18096 -25720 19420 -25704
rect 19642 -7634 19691 -7617
rect 19642 -9010 19648 -7634
rect 19682 -9010 19691 -7634
rect 19642 -9144 19691 -9010
rect 19642 -10520 19648 -9144
rect 19682 -10520 19691 -9144
rect 19642 -10654 19691 -10520
rect 19642 -12030 19648 -10654
rect 19682 -12030 19691 -10654
rect 19642 -12164 19691 -12030
rect 19642 -13540 19648 -12164
rect 19682 -13540 19691 -12164
rect 19642 -13674 19691 -13540
rect 19642 -15050 19648 -13674
rect 19682 -15050 19691 -13674
rect 19642 -15184 19691 -15050
rect 19642 -16560 19648 -15184
rect 19682 -16560 19691 -15184
rect 19642 -16694 19691 -16560
rect 19642 -18070 19648 -16694
rect 19682 -18070 19691 -16694
rect 19642 -18204 19691 -18070
rect 19642 -19580 19648 -18204
rect 19682 -19580 19691 -18204
rect 19642 -19714 19691 -19580
rect 19642 -21090 19648 -19714
rect 19682 -21090 19691 -19714
rect 19642 -21224 19691 -21090
rect 19642 -22600 19648 -21224
rect 19682 -22600 19691 -21224
rect 19642 -22734 19691 -22600
rect 19642 -24110 19648 -22734
rect 19682 -24110 19691 -22734
rect 19642 -24244 19691 -24110
rect 19642 -25620 19648 -24244
rect 19682 -25620 19691 -24244
rect 19642 -25720 19691 -25620
rect 19913 -7670 21244 -7584
rect 21306 -7634 21340 -7618
rect 19913 -9060 21240 -7670
rect 21306 -9026 21340 -9010
rect 21278 -9094 21294 -9060
rect 19913 -10570 21240 -9094
rect 21306 -9144 21340 -9128
rect 21306 -10536 21340 -10520
rect 21278 -10604 21294 -10570
rect 19913 -12080 21240 -10604
rect 21306 -10654 21340 -10638
rect 21306 -12046 21340 -12030
rect 21278 -12114 21294 -12080
rect 19913 -13590 21240 -12114
rect 21306 -12164 21340 -12148
rect 21306 -13556 21340 -13540
rect 21278 -13624 21294 -13590
rect 19913 -15100 21240 -13624
rect 21306 -13674 21340 -13658
rect 21306 -15066 21340 -15050
rect 21278 -15134 21294 -15100
rect 19913 -16610 21240 -15134
rect 21306 -15184 21340 -15168
rect 21306 -16576 21340 -16560
rect 21278 -16644 21294 -16610
rect 19913 -18120 21240 -16644
rect 21306 -16694 21340 -16678
rect 21306 -18086 21340 -18070
rect 21278 -18154 21294 -18120
rect 19913 -19630 21240 -18154
rect 21306 -18204 21340 -18188
rect 21306 -19596 21340 -19580
rect 21278 -19664 21294 -19630
rect 19913 -21140 21240 -19664
rect 21306 -19714 21340 -19698
rect 21306 -21106 21340 -21090
rect 21278 -21174 21294 -21140
rect 19913 -22650 21240 -21174
rect 21306 -21224 21340 -21208
rect 21306 -22616 21340 -22600
rect 21278 -22684 21294 -22650
rect 19913 -24160 21240 -22684
rect 21306 -22734 21340 -22718
rect 21306 -24126 21340 -24110
rect 21278 -24194 21294 -24160
rect 19913 -25670 21240 -24194
rect 21306 -24244 21340 -24228
rect 21306 -25636 21340 -25620
rect 21278 -25704 21294 -25670
rect 19913 -25720 21240 -25704
<< viali >>
rect -18978 55462 -17592 56190
rect -14978 55462 -13592 56190
rect -10978 55462 -9592 56190
rect -6978 55462 -5592 56190
rect -2978 55462 -1592 56190
rect 1022 55462 2408 56190
rect 5022 55462 6408 56190
rect 9022 55462 10408 56190
rect 13022 55462 14408 56190
rect 17022 55462 18408 56190
rect 21022 55462 22408 56190
rect 25022 55462 26408 56190
rect 29022 55462 30408 56190
rect 33022 55462 34408 56190
rect 37022 55462 38408 56190
rect -20714 53298 -19328 54026
rect 37064 52260 38450 52988
rect -20714 49298 -19328 50026
rect -16240 49265 -16202 49662
rect -15922 49265 -15884 49662
rect -15604 49265 -15566 49662
rect -15286 49265 -15248 49662
rect 37064 48260 38450 48988
rect -20714 45298 -19328 46026
rect -16240 44108 -16202 44505
rect -15922 44108 -15884 44505
rect -15604 44108 -15566 44505
rect -15286 44108 -15248 44505
rect 37064 44260 38450 44988
rect -15530 42384 -15458 42386
rect -20714 41298 -19328 42026
rect -16188 41987 -16150 42384
rect -15852 41952 -15848 42384
rect -15848 41952 -15780 42384
rect -15530 41954 -15460 42384
rect -15460 41954 -15458 42384
rect -15116 41951 -15078 42348
rect 37064 40260 38450 40988
rect -20714 37298 -19328 38026
rect -16188 36830 -16150 37227
rect -15850 36794 -15848 37226
rect -15848 36794 -15778 37226
rect -15532 36794 -15530 37222
rect -15530 36794 -15460 37222
rect -15532 36790 -15460 36794
rect -15116 36794 -15078 37191
rect 37064 36260 38450 36988
rect -16196 35487 -16158 35884
rect -15876 35490 -15874 35922
rect -15874 35490 -15804 35922
rect -15556 35490 -15486 35922
rect -15486 35490 -15484 35922
rect -15170 35505 -15132 35902
rect -20714 33298 -19328 34026
rect 37064 32260 38450 32988
rect -16196 30330 -16158 30727
rect -15876 30332 -15874 30764
rect -15874 30332 -15804 30764
rect -15804 30332 -15802 30764
rect -15876 30330 -15802 30332
rect -15558 30332 -15556 30764
rect -15556 30332 -15486 30764
rect -15486 30332 -15484 30764
rect -15558 30330 -15484 30332
rect -15170 30348 -15132 30745
rect -20714 29298 -19328 30026
rect -16174 28735 -16136 29132
rect -15856 28735 -15818 29132
rect -15538 28735 -15500 29132
rect -15220 28735 -15182 29132
rect 37064 28260 38450 28988
rect -20714 25298 -19328 26026
rect 37064 24260 38450 24988
rect -16174 23578 -16136 23975
rect -15856 23578 -15818 23975
rect -15538 23578 -15500 23975
rect -15220 23578 -15182 23975
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -94610 20212 -94576 20556
rect -94610 19524 -94576 20212
rect -94610 19180 -94576 19524
rect -92952 20212 -92918 20556
rect -92952 19524 -92918 20212
rect -92952 19180 -92918 19524
rect -96044 17274 -95512 17740
rect -94610 18576 -94576 18920
rect -94610 17888 -94576 18576
rect -94610 17544 -94576 17888
rect -91294 20212 -91260 20556
rect -91294 19524 -91260 20212
rect -91294 19180 -91260 19524
rect -92952 18576 -92918 18920
rect -92952 17888 -92918 18576
rect -92952 17544 -92918 17888
rect -94608 16830 -94574 17174
rect -94608 16142 -94574 16830
rect -94608 15798 -94574 16142
rect -96044 15274 -95512 15740
rect -89636 20212 -89602 20556
rect -89636 19524 -89602 20212
rect -89636 19180 -89602 19524
rect -91294 18576 -91260 18920
rect -91294 17888 -91260 18576
rect -91294 17544 -91260 17888
rect -92950 16830 -92916 17174
rect -92950 16142 -92916 16830
rect -92950 15798 -92916 16142
rect -94608 15194 -94574 15538
rect -94608 14506 -94574 15194
rect -94608 14162 -94574 14506
rect -87978 20212 -87944 20556
rect -87978 19524 -87944 20212
rect -87978 19180 -87944 19524
rect -89636 18576 -89602 18920
rect -89636 17888 -89602 18576
rect -89636 17544 -89602 17888
rect -91292 16830 -91258 17174
rect -91292 16142 -91258 16830
rect -91292 15798 -91258 16142
rect -92950 15194 -92916 15538
rect -92950 14506 -92916 15194
rect -92950 14162 -92916 14506
rect -96044 13274 -95512 13740
rect -94608 13558 -94574 13902
rect -94608 12870 -94574 13558
rect -94608 12526 -94574 12870
rect -86320 20212 -86286 20556
rect -86320 19524 -86286 20212
rect -86320 19180 -86286 19524
rect -87978 18576 -87944 18920
rect -87978 17888 -87944 18576
rect -87978 17544 -87944 17888
rect -89634 16830 -89600 17174
rect -89634 16142 -89600 16830
rect -89634 15798 -89600 16142
rect -91292 15194 -91258 15538
rect -91292 14506 -91258 15194
rect -91292 14162 -91258 14506
rect -92950 13558 -92916 13902
rect -92950 12870 -92916 13558
rect -92950 12526 -92916 12870
rect -96044 11274 -95512 11740
rect -94608 11922 -94574 12266
rect -94608 11234 -94574 11922
rect -94608 10890 -94574 11234
rect -84662 20212 -84628 20556
rect -84662 19524 -84628 20212
rect -84662 19180 -84628 19524
rect -86320 18576 -86286 18920
rect -86320 17888 -86286 18576
rect -86320 17544 -86286 17888
rect -87976 16830 -87942 17174
rect -87976 16142 -87942 16830
rect -87976 15798 -87942 16142
rect -89634 15194 -89600 15538
rect -89634 14506 -89600 15194
rect -89634 14162 -89600 14506
rect -91292 13558 -91258 13902
rect -91292 12870 -91258 13558
rect -91292 12526 -91258 12870
rect -92950 11922 -92916 12266
rect -92950 11234 -92916 11922
rect -92950 10890 -92916 11234
rect -96044 9274 -95512 9740
rect -94608 10284 -94574 10628
rect -94608 9596 -94574 10284
rect -94608 9252 -94574 9596
rect -83004 20212 -82970 20556
rect -83004 19524 -82970 20212
rect -83004 19180 -82970 19524
rect -84662 18576 -84628 18920
rect -84662 17888 -84628 18576
rect -84662 17544 -84628 17888
rect -86318 16830 -86284 17174
rect -86318 16142 -86284 16830
rect -86318 15798 -86284 16142
rect -87976 15194 -87942 15538
rect -87976 14506 -87942 15194
rect -87976 14162 -87942 14506
rect -89634 13558 -89600 13902
rect -89634 12870 -89600 13558
rect -89634 12526 -89600 12870
rect -91292 11922 -91258 12266
rect -91292 11234 -91258 11922
rect -91292 10890 -91258 11234
rect -92950 10284 -92916 10628
rect -92950 9596 -92916 10284
rect -92950 9252 -92916 9596
rect -96044 7274 -95512 7740
rect -94608 8648 -94574 8992
rect -94608 7960 -94574 8648
rect -94608 7616 -94574 7960
rect -81346 20212 -81312 20556
rect -81346 19524 -81312 20212
rect -81346 19180 -81312 19524
rect -83004 18576 -82970 18920
rect -83004 17888 -82970 18576
rect -83004 17544 -82970 17888
rect -84660 16830 -84626 17174
rect -84660 16142 -84626 16830
rect -84660 15798 -84626 16142
rect -86318 15194 -86284 15538
rect -86318 14506 -86284 15194
rect -86318 14162 -86284 14506
rect -87976 13558 -87942 13902
rect -87976 12870 -87942 13558
rect -87976 12526 -87942 12870
rect -89634 11922 -89600 12266
rect -89634 11234 -89600 11922
rect -89634 10890 -89600 11234
rect -91292 10284 -91258 10628
rect -91292 9596 -91258 10284
rect -91292 9252 -91258 9596
rect -92950 8648 -92916 8992
rect -92950 7960 -92916 8648
rect -92950 7616 -92916 7960
rect -94608 7012 -94574 7356
rect -94608 6324 -94574 7012
rect -94608 5980 -94574 6324
rect -96044 5274 -95512 5740
rect -79688 20212 -79654 20556
rect -79688 19524 -79654 20212
rect -79688 19180 -79654 19524
rect -81346 18576 -81312 18920
rect -81346 17888 -81312 18576
rect -81346 17544 -81312 17888
rect -83002 16830 -82968 17174
rect -83002 16142 -82968 16830
rect -83002 15798 -82968 16142
rect -84660 15194 -84626 15538
rect -84660 14506 -84626 15194
rect -84660 14162 -84626 14506
rect -86318 13558 -86284 13902
rect -86318 12870 -86284 13558
rect -86318 12526 -86284 12870
rect -87976 11922 -87942 12266
rect -87976 11234 -87942 11922
rect -87976 10890 -87942 11234
rect -89634 10284 -89600 10628
rect -89634 9596 -89600 10284
rect -89634 9252 -89600 9596
rect -91292 8648 -91258 8992
rect -91292 7960 -91258 8648
rect -91292 7616 -91258 7960
rect -92950 7012 -92916 7356
rect -92950 6324 -92916 7012
rect -92950 5980 -92916 6324
rect -94608 5376 -94574 5720
rect -94608 4688 -94574 5376
rect -94608 4344 -94574 4688
rect -78030 20212 -77996 20556
rect -78030 19524 -77996 20212
rect -78030 19180 -77996 19524
rect -79688 18576 -79654 18920
rect -79688 17888 -79654 18576
rect -79688 17544 -79654 17888
rect -81344 16830 -81310 17174
rect -81344 16142 -81310 16830
rect -81344 15798 -81310 16142
rect -83002 15194 -82968 15538
rect -83002 14506 -82968 15194
rect -83002 14162 -82968 14506
rect -84660 13558 -84626 13902
rect -84660 12870 -84626 13558
rect -84660 12526 -84626 12870
rect -86318 11922 -86284 12266
rect -86318 11234 -86284 11922
rect -86318 10890 -86284 11234
rect -87976 10284 -87942 10628
rect -87976 9596 -87942 10284
rect -87976 9252 -87942 9596
rect -89634 8648 -89600 8992
rect -89634 7960 -89600 8648
rect -89634 7616 -89600 7960
rect -91292 7012 -91258 7356
rect -91292 6324 -91258 7012
rect -91292 5980 -91258 6324
rect -92950 5376 -92916 5720
rect -92950 4688 -92916 5376
rect -92950 4344 -92916 4688
rect -76372 20212 -76338 20556
rect -76372 19524 -76338 20212
rect -76372 19180 -76338 19524
rect -74714 20212 -74680 20556
rect -74714 19524 -74680 20212
rect -74714 19180 -74680 19524
rect -78030 18576 -77996 18920
rect -78030 17888 -77996 18576
rect -78030 17544 -77996 17888
rect -79686 16830 -79652 17174
rect -79686 16142 -79652 16830
rect -79686 15798 -79652 16142
rect -81344 15194 -81310 15538
rect -81344 14506 -81310 15194
rect -81344 14162 -81310 14506
rect -83002 13558 -82968 13902
rect -83002 12870 -82968 13558
rect -83002 12526 -82968 12870
rect -84660 11922 -84626 12266
rect -84660 11234 -84626 11922
rect -84660 10890 -84626 11234
rect -86318 10284 -86284 10628
rect -86318 9596 -86284 10284
rect -86318 9252 -86284 9596
rect -87976 8648 -87942 8992
rect -87976 7960 -87942 8648
rect -87976 7616 -87942 7960
rect -89634 7012 -89600 7356
rect -89634 6324 -89600 7012
rect -89634 5980 -89600 6324
rect -91292 5376 -91258 5720
rect -91292 4688 -91258 5376
rect -91292 4344 -91258 4688
rect -76372 18576 -76338 18920
rect -76372 17888 -76338 18576
rect -76372 17544 -76338 17888
rect -73056 20212 -73022 20556
rect -73056 19524 -73022 20212
rect -73056 19180 -73022 19524
rect -74714 18576 -74680 18920
rect -74714 17888 -74680 18576
rect -74714 17544 -74680 17888
rect -78028 16830 -77994 17174
rect -78028 16142 -77994 16830
rect -78028 15798 -77994 16142
rect -79686 15194 -79652 15538
rect -79686 14506 -79652 15194
rect -79686 14162 -79652 14506
rect -81344 13558 -81310 13902
rect -81344 12870 -81310 13558
rect -81344 12526 -81310 12870
rect -83002 11922 -82968 12266
rect -83002 11234 -82968 11922
rect -83002 10890 -82968 11234
rect -84660 10284 -84626 10628
rect -84660 9596 -84626 10284
rect -84660 9252 -84626 9596
rect -86318 8648 -86284 8992
rect -86318 7960 -86284 8648
rect -86318 7616 -86284 7960
rect -87976 7012 -87942 7356
rect -87976 6324 -87942 7012
rect -87976 5980 -87942 6324
rect -89634 5376 -89600 5720
rect -89634 4688 -89600 5376
rect -89634 4344 -89600 4688
rect -76370 16830 -76336 17174
rect -76370 16142 -76336 16830
rect -76370 15798 -76336 16142
rect -71398 20212 -71364 20556
rect -71398 19524 -71364 20212
rect -71398 19180 -71364 19524
rect -73056 18576 -73022 18920
rect -73056 17888 -73022 18576
rect -73056 17544 -73022 17888
rect -74712 16830 -74678 17174
rect -74712 16142 -74678 16830
rect -74712 15798 -74678 16142
rect -78028 15194 -77994 15538
rect -78028 14506 -77994 15194
rect -78028 14162 -77994 14506
rect -79686 13558 -79652 13902
rect -79686 12870 -79652 13558
rect -79686 12526 -79652 12870
rect -81344 11922 -81310 12266
rect -81344 11234 -81310 11922
rect -81344 10890 -81310 11234
rect -83002 10284 -82968 10628
rect -83002 9596 -82968 10284
rect -83002 9252 -82968 9596
rect -84660 8648 -84626 8992
rect -84660 7960 -84626 8648
rect -84660 7616 -84626 7960
rect -86318 7012 -86284 7356
rect -86318 6324 -86284 7012
rect -86318 5980 -86284 6324
rect -87976 5376 -87942 5720
rect -87976 4688 -87942 5376
rect -87976 4344 -87942 4688
rect -76370 15194 -76336 15538
rect -76370 14506 -76336 15194
rect -76370 14162 -76336 14506
rect -69740 20212 -69706 20556
rect -69740 19524 -69706 20212
rect -69740 19180 -69706 19524
rect -71398 18576 -71364 18920
rect -71398 17888 -71364 18576
rect -71398 17544 -71364 17888
rect -73054 16830 -73020 17174
rect -73054 16142 -73020 16830
rect -73054 15798 -73020 16142
rect -74712 15194 -74678 15538
rect -74712 14506 -74678 15194
rect -74712 14162 -74678 14506
rect -78028 13558 -77994 13902
rect -78028 12870 -77994 13558
rect -78028 12526 -77994 12870
rect -79686 11922 -79652 12266
rect -79686 11234 -79652 11922
rect -79686 10890 -79652 11234
rect -81344 10284 -81310 10628
rect -81344 9596 -81310 10284
rect -81344 9252 -81310 9596
rect -83002 8648 -82968 8992
rect -83002 7960 -82968 8648
rect -83002 7616 -82968 7960
rect -84660 7012 -84626 7356
rect -84660 6324 -84626 7012
rect -84660 5980 -84626 6324
rect -86318 5376 -86284 5720
rect -86318 4688 -86284 5376
rect -86318 4344 -86284 4688
rect -76370 13558 -76336 13902
rect -76370 12870 -76336 13558
rect -76370 12526 -76336 12870
rect -68082 20212 -68048 20556
rect -68082 19524 -68048 20212
rect -68082 19180 -68048 19524
rect -69740 18576 -69706 18920
rect -69740 17888 -69706 18576
rect -69740 17544 -69706 17888
rect -71396 16830 -71362 17174
rect -71396 16142 -71362 16830
rect -71396 15798 -71362 16142
rect -73054 15194 -73020 15538
rect -73054 14506 -73020 15194
rect -73054 14162 -73020 14506
rect -74712 13558 -74678 13902
rect -74712 12870 -74678 13558
rect -74712 12526 -74678 12870
rect -78028 11922 -77994 12266
rect -78028 11234 -77994 11922
rect -78028 10890 -77994 11234
rect -79686 10284 -79652 10628
rect -79686 9596 -79652 10284
rect -79686 9252 -79652 9596
rect -81344 8648 -81310 8992
rect -81344 7960 -81310 8648
rect -81344 7616 -81310 7960
rect -83002 7012 -82968 7356
rect -83002 6324 -82968 7012
rect -83002 5980 -82968 6324
rect -84660 5376 -84626 5720
rect -84660 4688 -84626 5376
rect -84660 4344 -84626 4688
rect -76370 11922 -76336 12266
rect -76370 11234 -76336 11922
rect -76370 10890 -76336 11234
rect -66424 20212 -66390 20556
rect -66424 19524 -66390 20212
rect -66424 19180 -66390 19524
rect -68082 18576 -68048 18920
rect -68082 17888 -68048 18576
rect -68082 17544 -68048 17888
rect -69738 16830 -69704 17174
rect -69738 16142 -69704 16830
rect -69738 15798 -69704 16142
rect -71396 15194 -71362 15538
rect -71396 14506 -71362 15194
rect -71396 14162 -71362 14506
rect -73054 13558 -73020 13902
rect -73054 12870 -73020 13558
rect -73054 12526 -73020 12870
rect -74712 11922 -74678 12266
rect -74712 11234 -74678 11922
rect -74712 10890 -74678 11234
rect -78028 10284 -77994 10628
rect -78028 9596 -77994 10284
rect -78028 9252 -77994 9596
rect -79686 8648 -79652 8992
rect -79686 7960 -79652 8648
rect -79686 7616 -79652 7960
rect -81344 7012 -81310 7356
rect -81344 6324 -81310 7012
rect -81344 5980 -81310 6324
rect -83002 5376 -82968 5720
rect -83002 4688 -82968 5376
rect -83002 4344 -82968 4688
rect -76370 10284 -76336 10628
rect -76370 9596 -76336 10284
rect -76370 9252 -76336 9596
rect -64766 20212 -64732 20556
rect -64766 19524 -64732 20212
rect -64766 19180 -64732 19524
rect -66424 18576 -66390 18920
rect -66424 17888 -66390 18576
rect -66424 17544 -66390 17888
rect -68080 16830 -68046 17174
rect -68080 16142 -68046 16830
rect -68080 15798 -68046 16142
rect -69738 15194 -69704 15538
rect -69738 14506 -69704 15194
rect -69738 14162 -69704 14506
rect -71396 13558 -71362 13902
rect -71396 12870 -71362 13558
rect -71396 12526 -71362 12870
rect -73054 11922 -73020 12266
rect -73054 11234 -73020 11922
rect -73054 10890 -73020 11234
rect -74712 10284 -74678 10628
rect -74712 9596 -74678 10284
rect -74712 9252 -74678 9596
rect -78028 8648 -77994 8992
rect -78028 7960 -77994 8648
rect -78028 7616 -77994 7960
rect -79686 7012 -79652 7356
rect -79686 6324 -79652 7012
rect -79686 5980 -79652 6324
rect -81344 5376 -81310 5720
rect -81344 4688 -81310 5376
rect -81344 4344 -81310 4688
rect -76370 8648 -76336 8992
rect -76370 7960 -76336 8648
rect -76370 7616 -76336 7960
rect -63108 20212 -63074 20556
rect -63108 19524 -63074 20212
rect -63108 19180 -63074 19524
rect -64766 18576 -64732 18920
rect -64766 17888 -64732 18576
rect -64766 17544 -64732 17888
rect -66422 16830 -66388 17174
rect -66422 16142 -66388 16830
rect -66422 15798 -66388 16142
rect -68080 15194 -68046 15538
rect -68080 14506 -68046 15194
rect -68080 14162 -68046 14506
rect -69738 13558 -69704 13902
rect -69738 12870 -69704 13558
rect -69738 12526 -69704 12870
rect -71396 11922 -71362 12266
rect -71396 11234 -71362 11922
rect -71396 10890 -71362 11234
rect -73054 10284 -73020 10628
rect -73054 9596 -73020 10284
rect -73054 9252 -73020 9596
rect -74712 8648 -74678 8992
rect -74712 7960 -74678 8648
rect -74712 7616 -74678 7960
rect -78028 7012 -77994 7356
rect -78028 6324 -77994 7012
rect -78028 5980 -77994 6324
rect -79686 5376 -79652 5720
rect -79686 4688 -79652 5376
rect -79686 4344 -79652 4688
rect -76370 7012 -76336 7356
rect -76370 6324 -76336 7012
rect -76370 5980 -76336 6324
rect -61450 20212 -61416 20556
rect -61450 19524 -61416 20212
rect -61450 19180 -61416 19524
rect -63108 18576 -63074 18920
rect -63108 17888 -63074 18576
rect -63108 17544 -63074 17888
rect -64764 16830 -64730 17174
rect -64764 16142 -64730 16830
rect -64764 15798 -64730 16142
rect -66422 15194 -66388 15538
rect -66422 14506 -66388 15194
rect -66422 14162 -66388 14506
rect -68080 13558 -68046 13902
rect -68080 12870 -68046 13558
rect -68080 12526 -68046 12870
rect -69738 11922 -69704 12266
rect -69738 11234 -69704 11922
rect -69738 10890 -69704 11234
rect -71396 10284 -71362 10628
rect -71396 9596 -71362 10284
rect -71396 9252 -71362 9596
rect -73054 8648 -73020 8992
rect -73054 7960 -73020 8648
rect -73054 7616 -73020 7960
rect -74712 7012 -74678 7356
rect -74712 6324 -74678 7012
rect -74712 5980 -74678 6324
rect -78028 5376 -77994 5720
rect -78028 4688 -77994 5376
rect -78028 4344 -77994 4688
rect -76370 5376 -76336 5720
rect -76370 4688 -76336 5376
rect -76370 4344 -76336 4688
rect -59792 20212 -59758 20556
rect -59792 19524 -59758 20212
rect -59792 19180 -59758 19524
rect -61450 18576 -61416 18920
rect -61450 17888 -61416 18576
rect -61450 17544 -61416 17888
rect -63106 16830 -63072 17174
rect -63106 16142 -63072 16830
rect -63106 15798 -63072 16142
rect -64764 15194 -64730 15538
rect -64764 14506 -64730 15194
rect -64764 14162 -64730 14506
rect -66422 13558 -66388 13902
rect -66422 12870 -66388 13558
rect -66422 12526 -66388 12870
rect -68080 11922 -68046 12266
rect -68080 11234 -68046 11922
rect -68080 10890 -68046 11234
rect -69738 10284 -69704 10628
rect -69738 9596 -69704 10284
rect -69738 9252 -69704 9596
rect -71396 8648 -71362 8992
rect -71396 7960 -71362 8648
rect -71396 7616 -71362 7960
rect -73054 7012 -73020 7356
rect -73054 6324 -73020 7012
rect -73054 5980 -73020 6324
rect -74712 5376 -74678 5720
rect -74712 4688 -74678 5376
rect -74712 4344 -74678 4688
rect -58134 20212 -58100 20556
rect -58134 19524 -58100 20212
rect -58134 19180 -58100 19524
rect -59792 18576 -59758 18920
rect -59792 17888 -59758 18576
rect -59792 17544 -59758 17888
rect -61448 16830 -61414 17174
rect -61448 16142 -61414 16830
rect -61448 15798 -61414 16142
rect -63106 15194 -63072 15538
rect -63106 14506 -63072 15194
rect -63106 14162 -63072 14506
rect -64764 13558 -64730 13902
rect -64764 12870 -64730 13558
rect -64764 12526 -64730 12870
rect -66422 11922 -66388 12266
rect -66422 11234 -66388 11922
rect -66422 10890 -66388 11234
rect -68080 10284 -68046 10628
rect -68080 9596 -68046 10284
rect -68080 9252 -68046 9596
rect -69738 8648 -69704 8992
rect -69738 7960 -69704 8648
rect -69738 7616 -69704 7960
rect -71396 7012 -71362 7356
rect -71396 6324 -71362 7012
rect -71396 5980 -71362 6324
rect -73054 5376 -73020 5720
rect -73054 4688 -73020 5376
rect -73054 4344 -73020 4688
rect -56476 20212 -56442 20556
rect -56476 19524 -56442 20212
rect -56476 19180 -56442 19524
rect -58134 18576 -58100 18920
rect -58134 17888 -58100 18576
rect -58134 17544 -58100 17888
rect -59790 16830 -59756 17174
rect -59790 16142 -59756 16830
rect -59790 15798 -59756 16142
rect -61448 15194 -61414 15538
rect -61448 14506 -61414 15194
rect -61448 14162 -61414 14506
rect -63106 13558 -63072 13902
rect -63106 12870 -63072 13558
rect -63106 12526 -63072 12870
rect -64764 11922 -64730 12266
rect -64764 11234 -64730 11922
rect -64764 10890 -64730 11234
rect -66422 10284 -66388 10628
rect -66422 9596 -66388 10284
rect -66422 9252 -66388 9596
rect -68080 8648 -68046 8992
rect -68080 7960 -68046 8648
rect -68080 7616 -68046 7960
rect -69738 7012 -69704 7356
rect -69738 6324 -69704 7012
rect -69738 5980 -69704 6324
rect -71396 5376 -71362 5720
rect -71396 4688 -71362 5376
rect -71396 4344 -71362 4688
rect -54818 20212 -54784 20556
rect -54818 19524 -54784 20212
rect -54818 19180 -54784 19524
rect -56476 18576 -56442 18920
rect -56476 17888 -56442 18576
rect -56476 17544 -56442 17888
rect -58132 16830 -58098 17174
rect -58132 16142 -58098 16830
rect -58132 15798 -58098 16142
rect -59790 15194 -59756 15538
rect -59790 14506 -59756 15194
rect -59790 14162 -59756 14506
rect -61448 13558 -61414 13902
rect -61448 12870 -61414 13558
rect -61448 12526 -61414 12870
rect -63106 11922 -63072 12266
rect -63106 11234 -63072 11922
rect -63106 10890 -63072 11234
rect -64764 10284 -64730 10628
rect -64764 9596 -64730 10284
rect -64764 9252 -64730 9596
rect -66422 8648 -66388 8992
rect -66422 7960 -66388 8648
rect -66422 7616 -66388 7960
rect -68080 7012 -68046 7356
rect -68080 6324 -68046 7012
rect -68080 5980 -68046 6324
rect -69738 5376 -69704 5720
rect -69738 4688 -69704 5376
rect -69738 4344 -69704 4688
rect -53160 20212 -53126 20556
rect -53160 19524 -53126 20212
rect -53160 19180 -53126 19524
rect -54818 18576 -54784 18920
rect -54818 17888 -54784 18576
rect -54818 17544 -54784 17888
rect -56474 16830 -56440 17174
rect -56474 16142 -56440 16830
rect -56474 15798 -56440 16142
rect -58132 15194 -58098 15538
rect -58132 14506 -58098 15194
rect -58132 14162 -58098 14506
rect -59790 13558 -59756 13902
rect -59790 12870 -59756 13558
rect -59790 12526 -59756 12870
rect -61448 11922 -61414 12266
rect -61448 11234 -61414 11922
rect -61448 10890 -61414 11234
rect -63106 10284 -63072 10628
rect -63106 9596 -63072 10284
rect -63106 9252 -63072 9596
rect -64764 8648 -64730 8992
rect -64764 7960 -64730 8648
rect -64764 7616 -64730 7960
rect -66422 7012 -66388 7356
rect -66422 6324 -66388 7012
rect -66422 5980 -66388 6324
rect -68080 5376 -68046 5720
rect -68080 4688 -68046 5376
rect -68080 4344 -68046 4688
rect -51502 20212 -51468 20556
rect -51502 19524 -51468 20212
rect -51502 19180 -51468 19524
rect -53160 18576 -53126 18920
rect -53160 17888 -53126 18576
rect -53160 17544 -53126 17888
rect -54816 16830 -54782 17174
rect -54816 16142 -54782 16830
rect -54816 15798 -54782 16142
rect -56474 15194 -56440 15538
rect -56474 14506 -56440 15194
rect -56474 14162 -56440 14506
rect -58132 13558 -58098 13902
rect -58132 12870 -58098 13558
rect -58132 12526 -58098 12870
rect -59790 11922 -59756 12266
rect -59790 11234 -59756 11922
rect -59790 10890 -59756 11234
rect -61448 10284 -61414 10628
rect -61448 9596 -61414 10284
rect -61448 9252 -61414 9596
rect -63106 8648 -63072 8992
rect -63106 7960 -63072 8648
rect -63106 7616 -63072 7960
rect -64764 7012 -64730 7356
rect -64764 6324 -64730 7012
rect -64764 5980 -64730 6324
rect -66422 5376 -66388 5720
rect -66422 4688 -66388 5376
rect -66422 4344 -66388 4688
rect -49844 20212 -49810 20556
rect -49844 19524 -49810 20212
rect -49844 19180 -49810 19524
rect -51502 18576 -51468 18920
rect -51502 17888 -51468 18576
rect -51502 17544 -51468 17888
rect -53158 16830 -53124 17174
rect -53158 16142 -53124 16830
rect -53158 15798 -53124 16142
rect -54816 15194 -54782 15538
rect -54816 14506 -54782 15194
rect -54816 14162 -54782 14506
rect -56474 13558 -56440 13902
rect -56474 12870 -56440 13558
rect -56474 12526 -56440 12870
rect -58132 11922 -58098 12266
rect -58132 11234 -58098 11922
rect -58132 10890 -58098 11234
rect -59790 10284 -59756 10628
rect -59790 9596 -59756 10284
rect -59790 9252 -59756 9596
rect -61448 8648 -61414 8992
rect -61448 7960 -61414 8648
rect -61448 7616 -61414 7960
rect -63106 7012 -63072 7356
rect -63106 6324 -63072 7012
rect -63106 5980 -63072 6324
rect -64764 5376 -64730 5720
rect -64764 4688 -64730 5376
rect -64764 4344 -64730 4688
rect -48186 20212 -48152 20556
rect -48186 19524 -48152 20212
rect -48186 19180 -48152 19524
rect -49844 18576 -49810 18920
rect -49844 17888 -49810 18576
rect -49844 17544 -49810 17888
rect -51500 16830 -51466 17174
rect -51500 16142 -51466 16830
rect -51500 15798 -51466 16142
rect -53158 15194 -53124 15538
rect -53158 14506 -53124 15194
rect -53158 14162 -53124 14506
rect -54816 13558 -54782 13902
rect -54816 12870 -54782 13558
rect -54816 12526 -54782 12870
rect -56474 11922 -56440 12266
rect -56474 11234 -56440 11922
rect -56474 10890 -56440 11234
rect -58132 10284 -58098 10628
rect -58132 9596 -58098 10284
rect -58132 9252 -58098 9596
rect -59790 8648 -59756 8992
rect -59790 7960 -59756 8648
rect -59790 7616 -59756 7960
rect -61448 7012 -61414 7356
rect -61448 6324 -61414 7012
rect -61448 5980 -61414 6324
rect -63106 5376 -63072 5720
rect -63106 4688 -63072 5376
rect -63106 4344 -63072 4688
rect -46528 20212 -46494 20556
rect -46528 19524 -46494 20212
rect -46528 19180 -46494 19524
rect -48186 18576 -48152 18920
rect -48186 17888 -48152 18576
rect -48186 17544 -48152 17888
rect -49842 16830 -49808 17174
rect -49842 16142 -49808 16830
rect -49842 15798 -49808 16142
rect -51500 15194 -51466 15538
rect -51500 14506 -51466 15194
rect -51500 14162 -51466 14506
rect -53158 13558 -53124 13902
rect -53158 12870 -53124 13558
rect -53158 12526 -53124 12870
rect -54816 11922 -54782 12266
rect -54816 11234 -54782 11922
rect -54816 10890 -54782 11234
rect -56474 10284 -56440 10628
rect -56474 9596 -56440 10284
rect -56474 9252 -56440 9596
rect -58132 8648 -58098 8992
rect -58132 7960 -58098 8648
rect -58132 7616 -58098 7960
rect -59790 7012 -59756 7356
rect -59790 6324 -59756 7012
rect -59790 5980 -59756 6324
rect -61448 5376 -61414 5720
rect -61448 4688 -61414 5376
rect -61448 4344 -61414 4688
rect -44870 20212 -44836 20556
rect -44870 19524 -44836 20212
rect -44870 19180 -44836 19524
rect -46528 18576 -46494 18920
rect -46528 17888 -46494 18576
rect -46528 17544 -46494 17888
rect -48184 16830 -48150 17174
rect -48184 16142 -48150 16830
rect -48184 15798 -48150 16142
rect -49842 15194 -49808 15538
rect -49842 14506 -49808 15194
rect -49842 14162 -49808 14506
rect -51500 13558 -51466 13902
rect -51500 12870 -51466 13558
rect -51500 12526 -51466 12870
rect -53158 11922 -53124 12266
rect -53158 11234 -53124 11922
rect -53158 10890 -53124 11234
rect -54816 10284 -54782 10628
rect -54816 9596 -54782 10284
rect -54816 9252 -54782 9596
rect -56474 8648 -56440 8992
rect -56474 7960 -56440 8648
rect -56474 7616 -56440 7960
rect -58132 7012 -58098 7356
rect -58132 6324 -58098 7012
rect -58132 5980 -58098 6324
rect -59790 5376 -59756 5720
rect -59790 4688 -59756 5376
rect -59790 4344 -59756 4688
rect -61008 4251 -60994 4264
rect -60994 4251 -60974 4264
rect -61008 4230 -60974 4251
rect -43212 20212 -43178 20556
rect -43212 19524 -43178 20212
rect -43212 19180 -43178 19524
rect -44870 18576 -44836 18920
rect -44870 17888 -44836 18576
rect -44870 17544 -44836 17888
rect -46526 16830 -46492 17174
rect -46526 16142 -46492 16830
rect -46526 15798 -46492 16142
rect -48184 15194 -48150 15538
rect -48184 14506 -48150 15194
rect -48184 14162 -48150 14506
rect -49842 13558 -49808 13902
rect -49842 12870 -49808 13558
rect -49842 12526 -49808 12870
rect -51500 11922 -51466 12266
rect -51500 11234 -51466 11922
rect -51500 10890 -51466 11234
rect -53158 10284 -53124 10628
rect -53158 9596 -53124 10284
rect -53158 9252 -53124 9596
rect -54816 8648 -54782 8992
rect -54816 7960 -54782 8648
rect -54816 7616 -54782 7960
rect -56474 7012 -56440 7356
rect -56474 6324 -56440 7012
rect -56474 5980 -56440 6324
rect -58132 5376 -58098 5720
rect -58132 4688 -58098 5376
rect -58132 4344 -58098 4688
rect -41554 20212 -41520 20556
rect -41554 19524 -41520 20212
rect -41554 19180 -41520 19524
rect -43212 18576 -43178 18920
rect -43212 17888 -43178 18576
rect -43212 17544 -43178 17888
rect -44868 16830 -44834 17174
rect -44868 16142 -44834 16830
rect -44868 15798 -44834 16142
rect -46526 15194 -46492 15538
rect -46526 14506 -46492 15194
rect -46526 14162 -46492 14506
rect -48184 13558 -48150 13902
rect -48184 12870 -48150 13558
rect -48184 12526 -48150 12870
rect -49842 11922 -49808 12266
rect -49842 11234 -49808 11922
rect -49842 10890 -49808 11234
rect -51500 10284 -51466 10628
rect -51500 9596 -51466 10284
rect -51500 9252 -51466 9596
rect -53158 8648 -53124 8992
rect -53158 7960 -53124 8648
rect -53158 7616 -53124 7960
rect -54816 7012 -54782 7356
rect -54816 6324 -54782 7012
rect -54816 5980 -54782 6324
rect -56474 5376 -56440 5720
rect -56474 4688 -56440 5376
rect -56474 4344 -56440 4688
rect -39896 20212 -39862 20556
rect -39896 19524 -39862 20212
rect -39896 19180 -39862 19524
rect -41554 18576 -41520 18920
rect -41554 17888 -41520 18576
rect -41554 17544 -41520 17888
rect -43210 16830 -43176 17174
rect -43210 16142 -43176 16830
rect -43210 15798 -43176 16142
rect -44868 15194 -44834 15538
rect -44868 14506 -44834 15194
rect -44868 14162 -44834 14506
rect -46526 13558 -46492 13902
rect -46526 12870 -46492 13558
rect -46526 12526 -46492 12870
rect -48184 11922 -48150 12266
rect -48184 11234 -48150 11922
rect -48184 10890 -48150 11234
rect -49842 10284 -49808 10628
rect -49842 9596 -49808 10284
rect -49842 9252 -49808 9596
rect -51500 8648 -51466 8992
rect -51500 7960 -51466 8648
rect -51500 7616 -51466 7960
rect -53158 7012 -53124 7356
rect -53158 6324 -53124 7012
rect -53158 5980 -53124 6324
rect -54816 5376 -54782 5720
rect -54816 4688 -54782 5376
rect -54816 4344 -54782 4688
rect -38238 20212 -38204 20556
rect -38238 19524 -38204 20212
rect -38238 19180 -38204 19524
rect -39896 18576 -39862 18920
rect -39896 17888 -39862 18576
rect -39896 17544 -39862 17888
rect -41552 16830 -41518 17174
rect -41552 16142 -41518 16830
rect -41552 15798 -41518 16142
rect -43210 15194 -43176 15538
rect -43210 14506 -43176 15194
rect -43210 14162 -43176 14506
rect -44868 13558 -44834 13902
rect -44868 12870 -44834 13558
rect -44868 12526 -44834 12870
rect -46526 11922 -46492 12266
rect -46526 11234 -46492 11922
rect -46526 10890 -46492 11234
rect -48184 10284 -48150 10628
rect -48184 9596 -48150 10284
rect -48184 9252 -48150 9596
rect -49842 8648 -49808 8992
rect -49842 7960 -49808 8648
rect -49842 7616 -49808 7960
rect -51500 7012 -51466 7356
rect -51500 6324 -51466 7012
rect -51500 5980 -51466 6324
rect -53158 5376 -53124 5720
rect -53158 4688 -53124 5376
rect -53158 4344 -53124 4688
rect -36580 20212 -36546 20556
rect -36580 19524 -36546 20212
rect -36580 19180 -36546 19524
rect -38238 18576 -38204 18920
rect -38238 17888 -38204 18576
rect -38238 17544 -38204 17888
rect -39894 16830 -39860 17174
rect -39894 16142 -39860 16830
rect -39894 15798 -39860 16142
rect -41552 15194 -41518 15538
rect -41552 14506 -41518 15194
rect -41552 14162 -41518 14506
rect -43210 13558 -43176 13902
rect -43210 12870 -43176 13558
rect -43210 12526 -43176 12870
rect -44868 11922 -44834 12266
rect -44868 11234 -44834 11922
rect -44868 10890 -44834 11234
rect -46526 10284 -46492 10628
rect -46526 9596 -46492 10284
rect -46526 9252 -46492 9596
rect -48184 8648 -48150 8992
rect -48184 7960 -48150 8648
rect -48184 7616 -48150 7960
rect -49842 7012 -49808 7356
rect -49842 6324 -49808 7012
rect -49842 5980 -49808 6324
rect -51500 5376 -51466 5720
rect -51500 4688 -51466 5376
rect -51500 4344 -51466 4688
rect -34922 20212 -34888 20556
rect -34922 19524 -34888 20212
rect -34922 19180 -34888 19524
rect -36580 18576 -36546 18920
rect -36580 17888 -36546 18576
rect -36580 17544 -36546 17888
rect -38236 16830 -38202 17174
rect -38236 16142 -38202 16830
rect -38236 15798 -38202 16142
rect -39894 15194 -39860 15538
rect -39894 14506 -39860 15194
rect -39894 14162 -39860 14506
rect -41552 13558 -41518 13902
rect -41552 12870 -41518 13558
rect -41552 12526 -41518 12870
rect -43210 11922 -43176 12266
rect -43210 11234 -43176 11922
rect -43210 10890 -43176 11234
rect -44868 10284 -44834 10628
rect -44868 9596 -44834 10284
rect -44868 9252 -44834 9596
rect -46526 8648 -46492 8992
rect -46526 7960 -46492 8648
rect -46526 7616 -46492 7960
rect -48184 7012 -48150 7356
rect -48184 6324 -48150 7012
rect -48184 5980 -48150 6324
rect -49842 5376 -49808 5720
rect -49842 4688 -49808 5376
rect -49842 4344 -49808 4688
rect -33264 20212 -33230 20556
rect -33264 19524 -33230 20212
rect -33264 19180 -33230 19524
rect -34922 18576 -34888 18920
rect -34922 17888 -34888 18576
rect -34922 17544 -34888 17888
rect -36578 16830 -36544 17174
rect -36578 16142 -36544 16830
rect -36578 15798 -36544 16142
rect -38236 15194 -38202 15538
rect -38236 14506 -38202 15194
rect -38236 14162 -38202 14506
rect -39894 13558 -39860 13902
rect -39894 12870 -39860 13558
rect -39894 12526 -39860 12870
rect -41552 11922 -41518 12266
rect -41552 11234 -41518 11922
rect -41552 10890 -41518 11234
rect -43210 10284 -43176 10628
rect -43210 9596 -43176 10284
rect -43210 9252 -43176 9596
rect -44868 8648 -44834 8992
rect -44868 7960 -44834 8648
rect -44868 7616 -44834 7960
rect -46526 7012 -46492 7356
rect -46526 6324 -46492 7012
rect -46526 5980 -46492 6324
rect -48184 5376 -48150 5720
rect -48184 4688 -48150 5376
rect -48184 4344 -48150 4688
rect -31606 20212 -31572 20556
rect -31606 19524 -31572 20212
rect -31606 19180 -31572 19524
rect -33264 18576 -33230 18920
rect -33264 17888 -33230 18576
rect -33264 17544 -33230 17888
rect -34920 16830 -34886 17174
rect -34920 16142 -34886 16830
rect -34920 15798 -34886 16142
rect -36578 15194 -36544 15538
rect -36578 14506 -36544 15194
rect -36578 14162 -36544 14506
rect -38236 13558 -38202 13902
rect -38236 12870 -38202 13558
rect -38236 12526 -38202 12870
rect -39894 11922 -39860 12266
rect -39894 11234 -39860 11922
rect -39894 10890 -39860 11234
rect -41552 10284 -41518 10628
rect -41552 9596 -41518 10284
rect -41552 9252 -41518 9596
rect -43210 8648 -43176 8992
rect -43210 7960 -43176 8648
rect -43210 7616 -43176 7960
rect -44868 7012 -44834 7356
rect -44868 6324 -44834 7012
rect -44868 5980 -44834 6324
rect -46526 5376 -46492 5720
rect -46526 4688 -46492 5376
rect -46526 4344 -46492 4688
rect -29948 20212 -29914 20556
rect -29948 19524 -29914 20212
rect -29948 19180 -29914 19524
rect -31606 18576 -31572 18920
rect -31606 17888 -31572 18576
rect -31606 17544 -31572 17888
rect -33262 16830 -33228 17174
rect -33262 16142 -33228 16830
rect -33262 15798 -33228 16142
rect -34920 15194 -34886 15538
rect -34920 14506 -34886 15194
rect -34920 14162 -34886 14506
rect -36578 13558 -36544 13902
rect -36578 12870 -36544 13558
rect -36578 12526 -36544 12870
rect -38236 11922 -38202 12266
rect -38236 11234 -38202 11922
rect -38236 10890 -38202 11234
rect -39894 10284 -39860 10628
rect -39894 9596 -39860 10284
rect -39894 9252 -39860 9596
rect -41552 8648 -41518 8992
rect -41552 7960 -41518 8648
rect -41552 7616 -41518 7960
rect -43210 7012 -43176 7356
rect -43210 6324 -43176 7012
rect -43210 5980 -43176 6324
rect -44868 5376 -44834 5720
rect -44868 4688 -44834 5376
rect -44868 4344 -44834 4688
rect -28290 20212 -28256 20556
rect -28290 19524 -28256 20212
rect -28290 19180 -28256 19524
rect -20714 21298 -19328 22026
rect 37064 20260 38450 20988
rect -27644 19274 -27112 19740
rect -29948 18576 -29914 18920
rect -29948 17888 -29914 18576
rect -29948 17544 -29914 17888
rect -31604 16830 -31570 17174
rect -31604 16142 -31570 16830
rect -31604 15798 -31570 16142
rect -33262 15194 -33228 15538
rect -33262 14506 -33228 15194
rect -33262 14162 -33228 14506
rect -34920 13558 -34886 13902
rect -34920 12870 -34886 13558
rect -34920 12526 -34886 12870
rect -36578 11922 -36544 12266
rect -36578 11234 -36544 11922
rect -36578 10890 -36544 11234
rect -38236 10284 -38202 10628
rect -38236 9596 -38202 10284
rect -38236 9252 -38202 9596
rect -39894 8648 -39860 8992
rect -39894 7960 -39860 8648
rect -39894 7616 -39860 7960
rect -41552 7012 -41518 7356
rect -41552 6324 -41518 7012
rect -41552 5980 -41518 6324
rect -43210 5376 -43176 5720
rect -43210 4688 -43176 5376
rect -43210 4344 -43176 4688
rect -28290 18576 -28256 18920
rect -28290 17888 -28256 18576
rect -28290 17544 -28256 17888
rect -29946 16830 -29912 17174
rect -29946 16142 -29912 16830
rect -29946 15798 -29912 16142
rect -31604 15194 -31570 15538
rect -31604 14506 -31570 15194
rect -31604 14162 -31570 14506
rect -33262 13558 -33228 13902
rect -33262 12870 -33228 13558
rect -33262 12526 -33228 12870
rect -34920 11922 -34886 12266
rect -34920 11234 -34886 11922
rect -34920 10890 -34886 11234
rect -36578 10284 -36544 10628
rect -36578 9596 -36544 10284
rect -36578 9252 -36544 9596
rect -38236 8648 -38202 8992
rect -38236 7960 -38202 8648
rect -38236 7616 -38202 7960
rect -39894 7012 -39860 7356
rect -39894 6324 -39860 7012
rect -39894 5980 -39860 6324
rect -41552 5376 -41518 5720
rect -41552 4688 -41518 5376
rect -41552 4344 -41518 4688
rect -27644 17274 -27112 17740
rect -28288 16830 -28254 17174
rect -28288 16142 -28254 16830
rect -28288 15798 -28254 16142
rect -29946 15194 -29912 15538
rect -29946 14506 -29912 15194
rect -29946 14162 -29912 14506
rect -31604 13558 -31570 13902
rect -31604 12870 -31570 13558
rect -31604 12526 -31570 12870
rect -33262 11922 -33228 12266
rect -33262 11234 -33228 11922
rect -33262 10890 -33228 11234
rect -34920 10284 -34886 10628
rect -34920 9596 -34886 10284
rect -34920 9252 -34886 9596
rect -36578 8648 -36544 8992
rect -36578 7960 -36544 8648
rect -36578 7616 -36544 7960
rect -38236 7012 -38202 7356
rect -38236 6324 -38202 7012
rect -38236 5980 -38202 6324
rect -39894 5376 -39860 5720
rect -39894 4688 -39860 5376
rect -39894 4344 -39860 4688
rect -20714 17298 -19328 18026
rect 37064 16260 38450 16988
rect -28288 15194 -28254 15538
rect -28288 14506 -28254 15194
rect -28288 14162 -28254 14506
rect -27644 15274 -27112 15740
rect -29946 13558 -29912 13902
rect -29946 12870 -29912 13558
rect -29946 12526 -29912 12870
rect -31604 11922 -31570 12266
rect -31604 11234 -31570 11922
rect -31604 10890 -31570 11234
rect -33262 10284 -33228 10628
rect -33262 9596 -33228 10284
rect -33262 9252 -33228 9596
rect -34920 8648 -34886 8992
rect -34920 7960 -34886 8648
rect -34920 7616 -34886 7960
rect -36578 7012 -36544 7356
rect -36578 6324 -36544 7012
rect -36578 5980 -36544 6324
rect -38236 5376 -38202 5720
rect -38236 4688 -38202 5376
rect -38236 4344 -38202 4688
rect -28288 13558 -28254 13902
rect -28288 12870 -28254 13558
rect -28288 12526 -28254 12870
rect -18052 14180 -16666 14908
rect -14052 14180 -12666 14908
rect -10052 14180 -8666 14908
rect -6052 14180 -4666 14908
rect -2052 14180 -666 14908
rect 1948 14180 3334 14908
rect 5948 14180 7334 14908
rect 9948 14180 11334 14908
rect 13948 14180 15334 14908
rect 17948 14180 19334 14908
rect 21948 14180 23334 14908
rect 25948 14180 27334 14908
rect 29948 14180 31334 14908
rect 33948 14180 35334 14908
rect -27644 13274 -27112 13740
rect -29946 11922 -29912 12266
rect -29946 11234 -29912 11922
rect -29946 10890 -29912 11234
rect -31604 10284 -31570 10628
rect -31604 9596 -31570 10284
rect -31604 9252 -31570 9596
rect -33262 8648 -33228 8992
rect -33262 7960 -33228 8648
rect -33262 7616 -33228 7960
rect -34920 7012 -34886 7356
rect -34920 6324 -34886 7012
rect -34920 5980 -34886 6324
rect -36578 5376 -36544 5720
rect -36578 4688 -36544 5376
rect -36578 4344 -36544 4688
rect -28288 11922 -28254 12266
rect -28288 11234 -28254 11922
rect -28288 10890 -28254 11234
rect -27644 11274 -27112 11740
rect 18000 11574 18960 12068
rect -29946 10284 -29912 10628
rect -29946 9596 -29912 10284
rect -29946 9252 -29912 9596
rect -31604 8648 -31570 8992
rect -31604 7960 -31570 8648
rect -31604 7616 -31570 7960
rect -33262 7012 -33228 7356
rect -33262 6324 -33228 7012
rect -33262 5980 -33228 6324
rect -34920 5376 -34886 5720
rect -34920 4688 -34886 5376
rect -34920 4344 -34886 4688
rect -28288 10284 -28254 10628
rect -28288 9596 -28254 10284
rect -28288 9252 -28254 9596
rect 142 10748 539 10786
rect 4423 10748 4820 10786
rect 5372 10748 5769 10786
rect 9653 10748 10050 10786
rect 10602 10748 10999 10786
rect 14883 10748 15280 10786
rect 15832 10748 16229 10786
rect 20113 10748 20510 10786
rect 142 10428 539 10466
rect 4423 10428 4820 10466
rect 5372 10428 5769 10466
rect 9653 10428 10050 10466
rect 10602 10428 10999 10466
rect 14883 10428 15280 10466
rect 15832 10428 16229 10466
rect 20113 10428 20510 10466
rect 142 10108 539 10146
rect 4423 10108 4820 10146
rect 5386 10086 5783 10124
rect 9667 10086 10064 10124
rect 10582 10088 10979 10126
rect 14863 10088 15260 10126
rect 15832 10108 16229 10146
rect 20113 10108 20510 10146
rect 142 9788 539 9826
rect 4423 9788 4820 9826
rect 5386 9768 5783 9806
rect 9667 9768 10064 9806
rect 10582 9770 10979 9808
rect 14863 9770 15260 9808
rect 15832 9788 16229 9826
rect 20113 9788 20510 9826
rect -27644 9274 -27112 9740
rect 142 9468 539 9506
rect 4423 9468 4820 9506
rect 5386 9450 5783 9488
rect 9667 9450 10064 9488
rect 10582 9452 10979 9490
rect 14863 9452 15260 9490
rect 15832 9468 16229 9506
rect 20113 9468 20510 9506
rect -29946 8648 -29912 8992
rect -29946 7960 -29912 8648
rect -29946 7616 -29912 7960
rect -31604 7012 -31570 7356
rect -31604 6324 -31570 7012
rect -31604 5980 -31570 6324
rect -33262 5376 -33228 5720
rect -33262 4688 -33228 5376
rect -33262 4344 -33228 4688
rect -28288 8648 -28254 8992
rect -28288 7960 -28254 8648
rect -28288 7616 -28254 7960
rect 142 9148 539 9186
rect 4423 9148 4820 9186
rect 5386 9132 5783 9170
rect 9667 9132 10064 9170
rect 10582 9134 10979 9172
rect 14863 9134 15260 9172
rect 15832 9148 16229 9186
rect 20113 9148 20510 9186
rect 142 8828 539 8866
rect 4423 8828 4820 8866
rect 5386 8814 5783 8852
rect 9667 8814 10064 8852
rect 10582 8816 10979 8854
rect 14863 8816 15260 8854
rect 15832 8828 16229 8866
rect 20113 8828 20510 8866
rect 142 8508 539 8546
rect 4423 8508 4820 8546
rect 5386 8496 5783 8534
rect 9667 8496 10064 8534
rect 10582 8498 10979 8536
rect 14863 8498 15260 8536
rect 15832 8508 16229 8546
rect 20113 8508 20510 8546
rect 142 8188 539 8226
rect 4423 8188 4820 8226
rect 5386 8178 5783 8216
rect 9667 8178 10064 8216
rect 10582 8180 10979 8218
rect 14863 8180 15260 8218
rect 15832 8188 16229 8226
rect 20113 8188 20510 8226
rect 142 7868 539 7906
rect 4423 7868 4820 7906
rect 5386 7860 5783 7898
rect 9667 7860 10064 7898
rect 10582 7862 10979 7900
rect 14863 7862 15260 7900
rect 15832 7868 16229 7906
rect 20113 7868 20510 7906
rect -29946 7012 -29912 7356
rect -29946 6324 -29912 7012
rect -29946 5980 -29912 6324
rect -31604 5376 -31570 5720
rect -31604 4688 -31570 5376
rect -31604 4344 -31570 4688
rect -28288 7012 -28254 7356
rect -28288 6324 -28254 7012
rect -28288 5980 -28254 6324
rect -27644 7274 -27112 7740
rect 142 7548 539 7586
rect 4423 7548 4820 7586
rect 5386 7542 5783 7580
rect 9667 7542 10064 7580
rect 10582 7544 10979 7582
rect 14863 7544 15260 7582
rect 15832 7548 16229 7586
rect 20113 7548 20510 7586
rect -29946 5376 -29912 5720
rect -29946 4688 -29912 5376
rect -29946 4344 -29912 4688
rect 142 7228 539 7266
rect 4423 7228 4820 7266
rect 5406 7196 5803 7234
rect 9687 7196 10084 7234
rect 10602 7226 10999 7264
rect 14883 7226 15280 7264
rect 15832 7228 16229 7266
rect 20113 7228 20510 7266
rect 142 6908 539 6946
rect 4423 6908 4820 6946
rect 5406 6876 5803 6914
rect 9687 6876 10084 6914
rect 10602 6908 10999 6946
rect 14883 6908 15280 6946
rect 15832 6908 16229 6946
rect 20113 6908 20510 6946
rect -28288 5376 -28254 5720
rect -28288 4688 -28254 5376
rect -28288 4344 -28254 4688
rect -27644 5274 -27112 5740
rect 7324 6356 7464 6480
rect 1374 5776 1700 6016
rect 2724 5963 2808 5997
rect 3926 5908 4050 6000
rect 5286 5975 5370 6009
rect -61904 3884 -61870 3918
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect -61770 3784 -61736 3878
rect -61770 3596 -61736 3784
rect -61770 3502 -61736 3596
rect -61674 3784 -61640 3878
rect -61674 3596 -61640 3784
rect -61674 3502 -61640 3596
rect -61578 3784 -61544 3878
rect -61578 3596 -61544 3784
rect -61578 3502 -61544 3596
rect -61482 3784 -61448 3878
rect -61482 3596 -61448 3784
rect -61482 3502 -61448 3596
rect -61386 3784 -61352 3878
rect -61386 3596 -61352 3784
rect -61386 3502 -61352 3596
rect 2620 5172 2654 5660
rect 2878 5172 2912 5660
rect 1074 4932 1108 5026
rect 1074 4744 1108 4932
rect 1074 4650 1108 4744
rect 1162 4932 1196 5026
rect 1162 4744 1196 4932
rect 1162 4650 1196 4744
rect 1306 4930 1340 5024
rect 1306 4742 1340 4930
rect 1306 4648 1340 4742
rect 1394 4930 1428 5024
rect 1394 4742 1428 4930
rect 1394 4648 1428 4742
rect 1534 4928 1568 5022
rect 1534 4740 1568 4928
rect 1534 4646 1568 4740
rect 1622 4928 1656 5022
rect 1622 4740 1656 4928
rect 1622 4646 1656 4740
rect 1752 4930 1786 5024
rect 1752 4742 1786 4930
rect 1752 4648 1786 4742
rect 1840 4930 1874 5024
rect 1840 4742 1874 4930
rect 1840 4648 1874 4742
rect 1098 4344 1132 4388
rect 1098 4256 1132 4344
rect 1098 4212 1132 4256
rect 1186 4344 1220 4388
rect 1186 4256 1220 4344
rect 1186 4212 1220 4256
rect 1314 4346 1348 4390
rect 1314 4258 1348 4346
rect 1314 4214 1348 4258
rect 1402 4346 1436 4390
rect 1402 4258 1436 4346
rect 1402 4214 1436 4258
rect 1532 4346 1566 4390
rect 1532 4258 1566 4346
rect 1532 4214 1566 4258
rect 1620 4346 1654 4390
rect 1620 4258 1654 4346
rect 1620 4214 1654 4258
rect 1754 4344 1788 4388
rect 1754 4256 1788 4344
rect 1754 4212 1788 4256
rect 1842 4344 1876 4388
rect 1842 4256 1876 4344
rect 5182 5184 5216 5672
rect 5440 5184 5474 5672
rect 1842 4212 1876 4256
rect 1426 4130 1466 4168
rect 1704 4130 1738 4164
rect 3668 4070 3862 4246
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect 4682 3790 4876 3966
rect 7630 6306 7682 6406
rect 7810 6318 7862 6402
rect 8534 6326 8612 6424
rect 10312 6320 10400 6452
rect 6262 5854 6588 6094
rect 6260 4950 6294 5044
rect 6260 4762 6294 4950
rect 6260 4668 6294 4762
rect 6348 4950 6382 5044
rect 6348 4762 6382 4950
rect 6348 4668 6382 4762
rect 6492 4948 6526 5042
rect 6492 4760 6526 4948
rect 6492 4666 6526 4760
rect 6580 4948 6614 5042
rect 6580 4760 6614 4948
rect 6580 4666 6614 4760
rect 6720 4946 6754 5040
rect 6720 4758 6754 4946
rect 6720 4664 6754 4758
rect 6808 4946 6842 5040
rect 6808 4758 6842 4946
rect 6808 4664 6842 4758
rect 6938 4948 6972 5042
rect 6938 4760 6972 4948
rect 6938 4666 6972 4760
rect 7026 4948 7060 5042
rect 7026 4760 7060 4948
rect 7026 4666 7060 4760
rect 6284 4362 6318 4406
rect 6284 4274 6318 4362
rect 6284 4230 6318 4274
rect 6372 4362 6406 4406
rect 6372 4274 6406 4362
rect 6372 4230 6406 4274
rect 6500 4364 6534 4408
rect 6500 4276 6534 4364
rect 6500 4232 6534 4276
rect 6588 4364 6622 4408
rect 6588 4276 6622 4364
rect 6588 4232 6622 4276
rect 6718 4364 6752 4408
rect 6718 4276 6752 4364
rect 6718 4232 6752 4276
rect 6806 4364 6840 4408
rect 6806 4276 6840 4364
rect 6806 4232 6840 4276
rect 6940 4362 6974 4406
rect 6940 4274 6974 4362
rect 6940 4230 6974 4274
rect 7028 4362 7062 4406
rect 7028 4274 7062 4362
rect 7028 4230 7062 4274
rect 6612 4148 6652 4186
rect 6890 4148 6924 4182
rect 5854 3958 5916 4026
rect -61818 3190 -61784 3234
rect -61818 3102 -61784 3190
rect -61818 3058 -61784 3102
rect -61722 3190 -61688 3234
rect -61722 3102 -61688 3190
rect -61722 3058 -61688 3102
rect -61626 3190 -61592 3234
rect -61626 3102 -61592 3190
rect -61626 3058 -61592 3102
rect -61530 3190 -61496 3234
rect -61530 3102 -61496 3190
rect -61530 3058 -61496 3102
rect -61434 3190 -61400 3234
rect -61434 3102 -61400 3190
rect -61434 3058 -61400 3102
rect -61864 2826 -61806 2878
rect -61464 2826 -61406 2878
rect 2730 2570 2814 2604
rect 3356 2572 3740 2606
rect 2626 2388 2660 2476
rect 2884 2388 2918 2476
rect 3102 2390 3136 2478
rect 4328 2572 4712 2606
rect 4074 2390 4108 2478
rect 5264 2570 5348 2604
rect 5160 2388 5194 2476
rect 5418 2388 5452 2476
rect 3524 1204 4484 1698
rect 9246 5928 9378 6012
rect 9902 5988 10058 6098
rect 12778 6106 12860 6192
rect 14218 6120 14278 6174
rect 8660 5703 8744 5737
rect 8556 4912 8590 5400
rect 8814 4912 8848 5400
rect 9022 5392 9080 5408
rect 9022 4904 9035 5392
rect 9035 4904 9069 5392
rect 9069 4904 9080 5392
rect 9022 4894 9080 4904
rect 9551 4904 9585 5386
rect 9551 4898 9585 4904
rect 9691 5394 9731 5424
rect 9691 4906 9693 5394
rect 9693 4906 9727 5394
rect 9727 4906 9731 5394
rect 9691 4900 9731 4906
rect 9248 4470 9382 4558
rect 10209 4906 10243 5388
rect 10209 4900 10243 4906
rect 10454 5677 10538 5711
rect 11574 5642 11900 5882
rect 10350 4886 10384 5374
rect 10608 4886 10642 5374
rect 10964 5216 11074 5292
rect 11436 4962 11470 5056
rect 10200 4298 10244 4366
rect 11198 4506 11274 4576
rect 10514 4142 10716 4264
rect 10514 3844 10720 3976
rect 8505 3664 8605 3765
rect 10738 3716 10862 3768
rect 9028 3559 9088 3574
rect 9028 3409 9044 3559
rect 9044 3409 9078 3559
rect 9078 3409 9088 3559
rect 9028 3382 9088 3409
rect 9032 3003 9092 3028
rect 9032 2853 9044 3003
rect 9044 2853 9078 3003
rect 9078 2853 9092 3003
rect 9554 3559 9614 3590
rect 9554 3409 9560 3559
rect 9560 3409 9594 3559
rect 9594 3409 9614 3559
rect 9554 3398 9614 3409
rect 9032 2836 9092 2853
rect 9556 3003 9612 3034
rect 9556 2853 9560 3003
rect 9560 2853 9594 3003
rect 9594 2853 9612 3003
rect 9556 2842 9612 2853
rect 8538 2528 8580 2568
rect 10042 3559 10102 3574
rect 10042 3409 10058 3559
rect 10058 3409 10092 3559
rect 10092 3409 10102 3559
rect 10042 3382 10102 3409
rect 10046 3003 10106 3028
rect 10046 2853 10058 3003
rect 10058 2853 10092 3003
rect 10092 2853 10106 3003
rect 10568 3559 10628 3590
rect 10568 3409 10574 3559
rect 10574 3409 10608 3559
rect 10608 3409 10628 3559
rect 10568 3398 10628 3409
rect 10046 2836 10106 2853
rect 10570 3003 10626 3034
rect 10570 2853 10574 3003
rect 10574 2853 10608 3003
rect 10608 2853 10626 3003
rect 10570 2842 10626 2853
rect 9616 2464 9736 2600
rect 10952 2452 11072 2544
rect 11436 4774 11470 4962
rect 11436 4680 11470 4774
rect 11524 4962 11558 5056
rect 11524 4774 11558 4962
rect 11524 4680 11558 4774
rect 11668 4960 11702 5054
rect 11668 4772 11702 4960
rect 11668 4678 11702 4772
rect 11756 4960 11790 5054
rect 11756 4772 11790 4960
rect 11756 4678 11790 4772
rect 11896 4958 11930 5052
rect 11896 4770 11930 4958
rect 11896 4676 11930 4770
rect 11984 4958 12018 5052
rect 11984 4770 12018 4958
rect 11984 4676 12018 4770
rect 12114 4960 12148 5054
rect 12114 4772 12148 4960
rect 12114 4678 12148 4772
rect 12202 4960 12236 5054
rect 12202 4772 12236 4960
rect 12202 4678 12236 4772
rect 11460 4374 11494 4418
rect 11460 4286 11494 4374
rect 11460 4242 11494 4286
rect 11548 4374 11582 4418
rect 11548 4286 11582 4374
rect 11548 4242 11582 4286
rect 11676 4376 11710 4420
rect 11676 4288 11710 4376
rect 11676 4244 11710 4288
rect 11764 4376 11798 4420
rect 11764 4288 11798 4376
rect 11764 4244 11798 4288
rect 11894 4376 11928 4420
rect 11894 4288 11928 4376
rect 11894 4244 11928 4288
rect 11982 4376 12016 4420
rect 11982 4288 12016 4376
rect 11982 4244 12016 4288
rect 12116 4374 12150 4418
rect 12116 4286 12150 4374
rect 12116 4242 12150 4286
rect 12204 4374 12238 4418
rect 12204 4286 12238 4374
rect 12204 4242 12238 4286
rect 11788 4160 11828 4198
rect 12066 4160 12100 4194
rect 12686 3272 12746 3376
rect 12308 2096 12452 2228
rect 9248 1956 9446 1960
rect 9248 1922 9261 1956
rect 9261 1922 9445 1956
rect 9445 1922 9446 1956
rect 9248 1920 9446 1922
rect 9859 1956 10063 1958
rect 9859 1922 10040 1956
rect 10040 1922 10063 1956
rect 9859 1920 10063 1922
rect 10946 1020 11906 1514
rect 13934 5575 14018 5609
rect 14378 5591 14562 5594
rect 14378 5557 14562 5591
rect 14378 5556 14562 5557
rect 13830 4784 13864 5272
rect 14088 4784 14122 5272
rect 16254 6060 16448 6124
rect 14782 5784 14842 5886
rect 14950 5591 15134 5596
rect 14950 5558 15134 5591
rect 16344 5954 16478 6004
rect 15522 5587 15606 5621
rect 17010 5584 17336 5824
rect 15418 4796 15452 5284
rect 15676 4796 15710 5284
rect 17092 4754 17126 4848
rect 17092 4566 17126 4754
rect 17092 4472 17126 4566
rect 17180 4754 17214 4848
rect 17180 4566 17214 4754
rect 17180 4472 17214 4566
rect 17324 4752 17358 4846
rect 17324 4564 17358 4752
rect 17324 4470 17358 4564
rect 17412 4752 17446 4846
rect 17412 4564 17446 4752
rect 17412 4470 17446 4564
rect 17552 4750 17586 4844
rect 17552 4562 17586 4750
rect 17552 4468 17586 4562
rect 17640 4750 17674 4844
rect 17640 4562 17674 4750
rect 17640 4468 17674 4562
rect 17770 4752 17804 4846
rect 17770 4564 17804 4752
rect 17770 4470 17804 4564
rect 17858 4752 17892 4846
rect 17858 4564 17892 4752
rect 17858 4470 17892 4564
rect 17116 4166 17150 4210
rect 17116 4078 17150 4166
rect 17116 4034 17150 4078
rect 17204 4166 17238 4210
rect 17204 4078 17238 4166
rect 17204 4034 17238 4078
rect 17332 4168 17366 4212
rect 17332 4080 17366 4168
rect 17332 4036 17366 4080
rect 17420 4168 17454 4212
rect 17420 4080 17454 4168
rect 17420 4036 17454 4080
rect 17550 4168 17584 4212
rect 17550 4080 17584 4168
rect 17550 4036 17584 4080
rect 17638 4168 17672 4212
rect 17638 4080 17672 4168
rect 17638 4036 17672 4080
rect 17772 4166 17806 4210
rect 17772 4078 17806 4166
rect 17772 4034 17806 4078
rect 17860 4166 17894 4210
rect 17860 4078 17894 4166
rect 17860 4034 17894 4078
rect 17444 3952 17484 3990
rect 17722 3952 17756 3986
rect 13422 3152 13506 3186
rect 13972 3018 14056 3052
rect 14230 3018 14314 3052
rect 14488 3018 14572 3052
rect 14972 3018 15056 3052
rect 15230 3018 15314 3052
rect 15488 3018 15572 3052
rect 16020 3102 16104 3136
rect 13318 1020 13352 2408
rect 13576 1020 13610 2408
rect 13972 2062 14056 2096
rect 14230 2062 14314 2096
rect 13972 1106 14056 1140
rect 14488 2062 14572 2096
rect 14230 1106 14314 1140
rect 14488 1106 14572 1140
rect 14972 2062 15056 2096
rect 15230 2062 15314 2096
rect 14972 1106 15056 1140
rect 15488 2062 15572 2096
rect 15230 1106 15314 1140
rect 15488 1106 15572 1140
rect 15916 970 15950 2358
rect 16174 970 16208 2358
rect 17578 1338 18538 1832
rect 26138 3246 26538 3638
rect 26886 2482 26920 2794
rect 26974 2482 27008 2794
rect 27090 2520 27124 2832
rect 27178 2832 27212 2834
rect 27178 2520 27212 2832
rect 27498 2490 27532 2802
rect 27586 2490 27620 2802
rect 27702 2528 27736 2840
rect 27790 2840 27824 2842
rect 27790 2528 27824 2840
rect 26690 2190 26780 2264
rect 26886 2072 26920 2196
rect 27078 2072 27112 2196
rect 28076 2486 28110 2798
rect 28164 2486 28198 2798
rect 28280 2524 28314 2836
rect 28368 2836 28402 2838
rect 28368 2524 28402 2836
rect 27498 2080 27532 2204
rect 27690 2080 27724 2204
rect 28650 2494 28684 2806
rect 28738 2494 28772 2806
rect 28854 2532 28888 2844
rect 28942 2844 28976 2846
rect 28942 2532 28976 2844
rect 28076 2076 28110 2200
rect 28268 2076 28302 2200
rect 29228 2494 29262 2806
rect 29316 2494 29350 2806
rect 29432 2532 29466 2844
rect 29520 2844 29554 2846
rect 29520 2532 29554 2844
rect 28650 2084 28684 2208
rect 28842 2084 28876 2208
rect 29806 2494 29840 2806
rect 29894 2494 29928 2806
rect 30010 2532 30044 2844
rect 30098 2844 30132 2846
rect 30098 2532 30132 2844
rect 29228 2084 29262 2208
rect 29420 2084 29454 2208
rect 30388 2498 30422 2810
rect 30476 2498 30510 2810
rect 30592 2536 30626 2848
rect 30680 2848 30714 2850
rect 30680 2536 30714 2848
rect 29806 2084 29840 2208
rect 29998 2084 30032 2208
rect 30964 2494 30998 2806
rect 31052 2494 31086 2806
rect 31168 2532 31202 2844
rect 31256 2844 31290 2846
rect 31256 2532 31290 2844
rect 31534 2490 31568 2802
rect 31622 2490 31656 2802
rect 31738 2528 31772 2840
rect 31826 2840 31860 2842
rect 31826 2528 31860 2840
rect 30388 2088 30422 2212
rect 30580 2088 30614 2212
rect 30964 2084 30998 2208
rect 31156 2084 31190 2208
rect 31320 2012 31382 2074
rect 31534 2080 31568 2204
rect 31726 2080 31760 2204
rect 32424 1746 32904 2206
rect 28280 428 28314 740
rect 28368 428 28402 740
rect 28480 466 28514 778
rect 28568 466 28602 778
rect 28682 426 28716 738
rect 28770 426 28804 738
rect 28280 -78 28314 234
rect 28368 -78 28402 234
rect 28480 -40 28514 272
rect 28568 -40 28602 272
rect 28680 -78 28714 234
rect 28768 -78 28802 234
rect 28280 -586 28314 -274
rect 28368 -586 28402 -274
rect 28480 -548 28514 -236
rect 28568 -548 28602 -236
rect 28680 -586 28714 -274
rect 28768 -586 28802 -274
rect 29808 -266 29842 358
rect 8763 -968 8797 -958
rect 8763 -992 8797 -968
rect 8855 -968 8889 -958
rect 8855 -992 8889 -968
rect 8947 -968 8981 -958
rect 8947 -992 8981 -968
rect 9039 -968 9073 -958
rect 9039 -992 9073 -968
rect 9131 -968 9165 -958
rect 9131 -992 9165 -968
rect 9223 -968 9257 -958
rect 9223 -992 9257 -968
rect 9315 -968 9349 -958
rect 9315 -992 9349 -968
rect 9407 -968 9441 -958
rect 9407 -992 9441 -968
rect 9499 -968 9533 -958
rect 9499 -992 9533 -968
rect 9591 -968 9625 -958
rect 9591 -992 9625 -968
rect 9683 -968 9717 -958
rect 9683 -992 9717 -968
rect 9775 -968 9809 -958
rect 9775 -992 9809 -968
rect 9867 -968 9901 -958
rect 9867 -992 9901 -968
rect 9959 -968 9993 -958
rect 9959 -992 9993 -968
rect 10051 -968 10085 -958
rect 10051 -992 10085 -968
rect 10143 -968 10177 -958
rect 10143 -992 10177 -968
rect 10235 -968 10269 -958
rect 10235 -992 10269 -968
rect 10327 -968 10361 -958
rect 10327 -992 10361 -968
rect 10419 -968 10453 -958
rect 10419 -992 10453 -968
rect 10511 -968 10545 -958
rect 10511 -992 10545 -968
rect 10603 -968 10637 -958
rect 10603 -992 10637 -968
rect 10695 -968 10729 -958
rect 10695 -992 10729 -968
rect 10787 -968 10821 -958
rect 10787 -992 10821 -968
rect 11229 -968 11263 -958
rect 11229 -992 11263 -968
rect 11321 -968 11355 -958
rect 11321 -992 11355 -968
rect 11413 -968 11447 -958
rect 11413 -992 11447 -968
rect 11505 -968 11539 -958
rect 11505 -992 11539 -968
rect 11597 -968 11631 -958
rect 11597 -992 11631 -968
rect 11689 -968 11723 -958
rect 11689 -992 11723 -968
rect 11781 -968 11815 -958
rect 11781 -992 11815 -968
rect 11873 -968 11907 -958
rect 11873 -992 11907 -968
rect 11965 -968 11999 -958
rect 11965 -992 11999 -968
rect 12057 -968 12091 -958
rect 12057 -992 12091 -968
rect 12149 -968 12183 -958
rect 12149 -992 12183 -968
rect 12241 -968 12275 -958
rect 12241 -992 12275 -968
rect 12333 -968 12367 -958
rect 12333 -992 12367 -968
rect 12425 -968 12459 -958
rect 12425 -992 12459 -968
rect 12517 -968 12551 -958
rect 12517 -992 12551 -968
rect 12609 -968 12643 -958
rect 12609 -992 12643 -968
rect 12701 -968 12735 -958
rect 12701 -992 12735 -968
rect 12793 -968 12827 -958
rect 12793 -992 12827 -968
rect 12885 -968 12919 -958
rect 12885 -992 12919 -968
rect 12977 -968 13011 -958
rect 12977 -992 13011 -968
rect 13069 -968 13103 -958
rect 13069 -992 13103 -968
rect 13161 -968 13195 -958
rect 13161 -992 13195 -968
rect 13253 -968 13287 -958
rect 13253 -992 13287 -968
rect 8856 -1289 8868 -1264
rect 8868 -1289 8890 -1264
rect 8856 -1298 8890 -1289
rect 8937 -1144 8971 -1128
rect 8937 -1162 8971 -1144
rect 9039 -1230 9073 -1196
rect 9315 -1162 9349 -1128
rect 9223 -1298 9257 -1264
rect 9939 -1154 9973 -1128
rect 9939 -1162 9970 -1154
rect 9970 -1162 9973 -1154
rect 9495 -1366 9529 -1332
rect 9567 -1350 9591 -1332
rect 9591 -1350 9601 -1332
rect 9567 -1366 9601 -1350
rect 9939 -1280 9973 -1264
rect 9939 -1298 9965 -1280
rect 9965 -1298 9973 -1280
rect 10155 -1278 10189 -1269
rect 10155 -1303 10171 -1278
rect 10171 -1303 10189 -1278
rect 10215 -1366 10249 -1332
rect 10488 -1301 10522 -1266
rect 10783 -1299 10817 -1265
rect 11230 -1270 11264 -1264
rect 11230 -1298 11232 -1270
rect 11232 -1298 11264 -1270
rect 11322 -1289 11334 -1264
rect 11334 -1289 11356 -1264
rect 11322 -1298 11356 -1289
rect 11403 -1144 11437 -1128
rect 11403 -1162 11437 -1144
rect 11505 -1230 11539 -1196
rect 11781 -1162 11815 -1128
rect 11689 -1298 11723 -1264
rect 12405 -1154 12439 -1128
rect 12405 -1162 12436 -1154
rect 12436 -1162 12439 -1154
rect 11961 -1366 11995 -1332
rect 12033 -1350 12057 -1332
rect 12057 -1350 12067 -1332
rect 12033 -1366 12067 -1350
rect 12405 -1280 12439 -1264
rect 12405 -1298 12431 -1280
rect 12431 -1298 12439 -1280
rect 12621 -1278 12655 -1269
rect 12621 -1303 12637 -1278
rect 12637 -1303 12655 -1278
rect 12681 -1366 12715 -1332
rect 13251 -1298 13285 -1264
rect 8763 -1530 8797 -1502
rect 8763 -1536 8797 -1530
rect 8855 -1530 8889 -1502
rect 8855 -1536 8889 -1530
rect 8947 -1530 8981 -1502
rect 8947 -1536 8981 -1530
rect 9039 -1530 9073 -1502
rect 9039 -1536 9073 -1530
rect 9131 -1530 9165 -1502
rect 9131 -1536 9165 -1530
rect 9223 -1530 9257 -1502
rect 9223 -1536 9257 -1530
rect 9315 -1530 9349 -1502
rect 9315 -1536 9349 -1530
rect 9407 -1530 9441 -1502
rect 9407 -1536 9441 -1530
rect 9499 -1530 9533 -1502
rect 9499 -1536 9533 -1530
rect 9591 -1530 9625 -1502
rect 9591 -1536 9625 -1530
rect 9683 -1530 9717 -1502
rect 9683 -1536 9717 -1530
rect 9775 -1530 9809 -1502
rect 9775 -1536 9809 -1530
rect 9867 -1530 9901 -1502
rect 9867 -1536 9901 -1530
rect 9959 -1530 9993 -1502
rect 9959 -1536 9993 -1530
rect 10051 -1530 10085 -1502
rect 10051 -1536 10085 -1530
rect 10143 -1530 10177 -1502
rect 10143 -1536 10177 -1530
rect 10235 -1530 10269 -1502
rect 10235 -1536 10269 -1530
rect 10327 -1530 10361 -1502
rect 10327 -1536 10361 -1530
rect 10419 -1530 10453 -1502
rect 10419 -1536 10453 -1530
rect 10511 -1530 10545 -1502
rect 10511 -1536 10545 -1530
rect 10603 -1530 10637 -1502
rect 10603 -1536 10637 -1530
rect 10695 -1530 10729 -1502
rect 10695 -1536 10729 -1530
rect 10787 -1530 10821 -1502
rect 10787 -1536 10821 -1530
rect 11229 -1529 11263 -1502
rect 11229 -1536 11263 -1529
rect 11321 -1529 11355 -1502
rect 11321 -1536 11355 -1529
rect 11413 -1529 11447 -1502
rect 11413 -1536 11447 -1529
rect 11505 -1529 11539 -1502
rect 11505 -1536 11539 -1529
rect 11597 -1529 11631 -1502
rect 11597 -1536 11631 -1529
rect 11689 -1529 11723 -1502
rect 11689 -1536 11723 -1529
rect 11781 -1529 11815 -1502
rect 11781 -1536 11815 -1529
rect 11873 -1529 11907 -1502
rect 11873 -1536 11907 -1529
rect 11965 -1529 11999 -1502
rect 11965 -1536 11999 -1529
rect 12057 -1529 12091 -1502
rect 12057 -1536 12091 -1529
rect 12149 -1529 12183 -1502
rect 12149 -1536 12183 -1529
rect 12241 -1529 12275 -1502
rect 12241 -1536 12275 -1529
rect 12333 -1529 12367 -1502
rect 12333 -1536 12367 -1529
rect 12425 -1529 12459 -1502
rect 12425 -1536 12459 -1529
rect 12517 -1529 12551 -1502
rect 12517 -1536 12551 -1529
rect 12609 -1529 12643 -1502
rect 12609 -1536 12643 -1529
rect 12701 -1529 12735 -1502
rect 12701 -1536 12735 -1529
rect 12793 -1529 12827 -1502
rect 12793 -1536 12827 -1529
rect 12885 -1529 12919 -1502
rect 12885 -1536 12919 -1529
rect 12977 -1529 13011 -1502
rect 12977 -1536 13011 -1529
rect 13069 -1529 13103 -1502
rect 13069 -1536 13103 -1529
rect 13161 -1529 13195 -1502
rect 13161 -1536 13195 -1529
rect 13253 -1529 13287 -1502
rect 13253 -1536 13287 -1529
rect 10181 -1770 10215 -1760
rect 10181 -1794 10215 -1770
rect 10273 -1770 10307 -1760
rect 10273 -1794 10307 -1770
rect 10365 -1770 10399 -1760
rect 10365 -1794 10399 -1770
rect 11229 -1769 11263 -1760
rect 11229 -1794 11263 -1769
rect 11321 -1769 11355 -1760
rect 11321 -1794 11355 -1769
rect 11413 -1769 11447 -1760
rect 11413 -1794 11447 -1769
rect 11505 -1769 11539 -1760
rect 11505 -1794 11539 -1769
rect 11597 -1769 11631 -1760
rect 11597 -1794 11631 -1769
rect 11689 -1769 11723 -1760
rect 11689 -1794 11723 -1769
rect 11781 -1769 11815 -1760
rect 11781 -1794 11815 -1769
rect 11873 -1769 11907 -1760
rect 11873 -1794 11907 -1769
rect 11965 -1769 11999 -1760
rect 11965 -1794 11999 -1769
rect 12057 -1769 12091 -1760
rect 12057 -1794 12091 -1769
rect 12149 -1769 12183 -1760
rect 12149 -1794 12183 -1769
rect 12241 -1769 12275 -1760
rect 12241 -1794 12275 -1769
rect 12333 -1769 12367 -1760
rect 12333 -1794 12367 -1769
rect 12425 -1769 12459 -1760
rect 12425 -1794 12459 -1769
rect 12517 -1769 12551 -1760
rect 12517 -1794 12551 -1769
rect 12609 -1769 12643 -1760
rect 12609 -1794 12643 -1769
rect 12701 -1769 12735 -1760
rect 12701 -1794 12735 -1769
rect 12793 -1769 12827 -1760
rect 12793 -1794 12827 -1769
rect 12885 -1769 12919 -1760
rect 12885 -1794 12919 -1769
rect 12977 -1769 13011 -1760
rect 12977 -1794 13011 -1769
rect 13069 -1769 13103 -1760
rect 13069 -1794 13103 -1769
rect 13161 -1769 13195 -1760
rect 13161 -1794 13195 -1769
rect 13253 -1769 13287 -1760
rect 13253 -1794 13287 -1769
rect 10181 -2072 10215 -2066
rect 10181 -2100 10189 -2072
rect 10189 -2100 10215 -2072
rect 10273 -2130 10307 -2096
rect 11230 -2066 11265 -2032
rect 11322 -2091 11334 -2066
rect 11334 -2091 11356 -2066
rect 11322 -2100 11356 -2091
rect 11403 -1946 11437 -1930
rect 11403 -1964 11437 -1946
rect 11505 -2062 11539 -2028
rect 11781 -1964 11815 -1930
rect 11689 -2100 11723 -2066
rect 12405 -1956 12439 -1930
rect 12405 -1964 12436 -1956
rect 12436 -1964 12439 -1956
rect 11961 -2168 11995 -2134
rect 12033 -2152 12057 -2134
rect 12057 -2152 12067 -2134
rect 12033 -2168 12067 -2152
rect 12405 -2082 12439 -2066
rect 12405 -2100 12431 -2082
rect 12431 -2100 12439 -2082
rect 12621 -2080 12655 -2071
rect 12621 -2105 12637 -2080
rect 12637 -2105 12655 -2080
rect 12681 -2168 12715 -2134
rect 13249 -2131 13283 -2097
rect 10181 -2330 10215 -2304
rect 10181 -2338 10215 -2330
rect 10273 -2330 10307 -2304
rect 10273 -2338 10307 -2330
rect 10365 -2330 10399 -2304
rect 10365 -2338 10399 -2330
rect 11229 -2332 11263 -2304
rect 11229 -2338 11263 -2332
rect 11321 -2332 11355 -2304
rect 11321 -2338 11355 -2332
rect 11413 -2332 11447 -2304
rect 11413 -2338 11447 -2332
rect 11505 -2332 11539 -2304
rect 11505 -2338 11539 -2332
rect 11597 -2332 11631 -2304
rect 11597 -2338 11631 -2332
rect 11689 -2332 11723 -2304
rect 11689 -2338 11723 -2332
rect 11781 -2332 11815 -2304
rect 11781 -2338 11815 -2332
rect 11873 -2332 11907 -2304
rect 11873 -2338 11907 -2332
rect 11965 -2332 11999 -2304
rect 11965 -2338 11999 -2332
rect 12057 -2332 12091 -2304
rect 12057 -2338 12091 -2332
rect 12149 -2332 12183 -2304
rect 12149 -2338 12183 -2332
rect 12241 -2332 12275 -2304
rect 12241 -2338 12275 -2332
rect 12333 -2332 12367 -2304
rect 12333 -2338 12367 -2332
rect 12425 -2332 12459 -2304
rect 12425 -2338 12459 -2332
rect 12517 -2332 12551 -2304
rect 12517 -2338 12551 -2332
rect 12609 -2332 12643 -2304
rect 12609 -2338 12643 -2332
rect 12701 -2332 12735 -2304
rect 12701 -2338 12735 -2332
rect 12793 -2332 12827 -2304
rect 12793 -2338 12827 -2332
rect 12885 -2332 12919 -2304
rect 12885 -2338 12919 -2332
rect 12977 -2332 13011 -2304
rect 12977 -2338 13011 -2332
rect 13069 -2332 13103 -2304
rect 13069 -2338 13103 -2332
rect 13161 -2332 13195 -2304
rect 13161 -2338 13195 -2332
rect 13253 -2332 13287 -2304
rect 13253 -2338 13287 -2332
rect -9129 -4238 -9095 -4228
rect -9129 -4262 -9095 -4238
rect -9037 -4238 -9003 -4228
rect -9037 -4262 -9003 -4238
rect -8945 -4238 -8911 -4228
rect -8945 -4262 -8911 -4238
rect -8853 -4238 -8819 -4228
rect -8853 -4262 -8819 -4238
rect -8761 -4238 -8727 -4228
rect -8761 -4262 -8727 -4238
rect -8669 -4238 -8635 -4228
rect -8669 -4262 -8635 -4238
rect -8577 -4238 -8543 -4228
rect -8577 -4262 -8543 -4238
rect -8485 -4238 -8451 -4228
rect -8485 -4262 -8451 -4238
rect -8393 -4238 -8359 -4228
rect -8393 -4262 -8359 -4238
rect -8301 -4238 -8267 -4228
rect -8301 -4262 -8267 -4238
rect -8209 -4238 -8175 -4228
rect -8209 -4262 -8175 -4238
rect -8117 -4238 -8083 -4228
rect -8117 -4262 -8083 -4238
rect -8025 -4238 -7991 -4228
rect -8025 -4262 -7991 -4238
rect -7933 -4238 -7899 -4228
rect -7933 -4262 -7899 -4238
rect -7841 -4238 -7807 -4228
rect -7841 -4262 -7807 -4238
rect -7749 -4238 -7715 -4228
rect -7749 -4262 -7715 -4238
rect -7657 -4238 -7623 -4228
rect -7657 -4262 -7623 -4238
rect -7565 -4238 -7531 -4228
rect -7565 -4262 -7531 -4238
rect -7473 -4238 -7439 -4228
rect -7473 -4262 -7439 -4238
rect -7381 -4238 -7347 -4228
rect -7381 -4262 -7347 -4238
rect -7289 -4238 -7255 -4228
rect -7289 -4262 -7255 -4238
rect -7197 -4238 -7163 -4228
rect -7197 -4262 -7163 -4238
rect -7105 -4238 -7071 -4228
rect -7105 -4262 -7071 -4238
rect -7013 -4238 -6979 -4228
rect -7013 -4262 -6979 -4238
rect -6921 -4238 -6887 -4228
rect -6921 -4262 -6887 -4238
rect -6829 -4238 -6795 -4228
rect -6829 -4262 -6795 -4238
rect -6737 -4238 -6703 -4228
rect -6737 -4262 -6703 -4238
rect -6645 -4238 -6611 -4228
rect -6645 -4262 -6611 -4238
rect -6553 -4238 -6519 -4228
rect -6553 -4262 -6519 -4238
rect -6461 -4238 -6427 -4228
rect -6461 -4262 -6427 -4238
rect -6369 -4238 -6335 -4228
rect -6369 -4262 -6335 -4238
rect -6277 -4238 -6243 -4228
rect -6277 -4262 -6243 -4238
rect -6185 -4238 -6151 -4228
rect -6185 -4262 -6151 -4238
rect -6093 -4238 -6059 -4228
rect -6093 -4262 -6059 -4238
rect -6001 -4238 -5967 -4228
rect -6001 -4262 -5967 -4238
rect -5909 -4238 -5875 -4228
rect -5909 -4262 -5875 -4238
rect -5817 -4238 -5783 -4228
rect -5817 -4262 -5783 -4238
rect -5725 -4238 -5691 -4228
rect -5725 -4262 -5691 -4238
rect -5633 -4238 -5599 -4228
rect -5633 -4262 -5599 -4238
rect -5541 -4238 -5507 -4228
rect -5541 -4262 -5507 -4238
rect -5449 -4238 -5415 -4228
rect -5449 -4262 -5415 -4238
rect -5357 -4238 -5323 -4228
rect -5357 -4262 -5323 -4238
rect -5265 -4238 -5231 -4228
rect -5265 -4262 -5231 -4238
rect -5173 -4238 -5139 -4228
rect -5173 -4262 -5139 -4238
rect -5081 -4238 -5047 -4228
rect -5081 -4262 -5047 -4238
rect -4989 -4238 -4955 -4228
rect -4989 -4262 -4955 -4238
rect -4897 -4238 -4863 -4228
rect -4897 -4262 -4863 -4238
rect -4805 -4238 -4771 -4228
rect -4805 -4262 -4771 -4238
rect -4713 -4238 -4679 -4228
rect -4713 -4262 -4679 -4238
rect -4621 -4238 -4587 -4228
rect -4621 -4262 -4587 -4238
rect -4529 -4238 -4495 -4228
rect -4529 -4262 -4495 -4238
rect -4437 -4238 -4403 -4228
rect -4437 -4262 -4403 -4238
rect -4345 -4238 -4311 -4228
rect -4345 -4262 -4311 -4238
rect -4253 -4238 -4219 -4228
rect -4253 -4262 -4219 -4238
rect -4161 -4238 -4127 -4228
rect -4161 -4262 -4127 -4238
rect -4069 -4238 -4035 -4228
rect -4069 -4262 -4035 -4238
rect -3977 -4238 -3943 -4228
rect -3977 -4262 -3943 -4238
rect -3885 -4238 -3851 -4228
rect -3885 -4262 -3851 -4238
rect -3793 -4238 -3759 -4228
rect -3793 -4262 -3759 -4238
rect -3701 -4238 -3667 -4228
rect -3701 -4262 -3667 -4238
rect -3609 -4238 -3575 -4228
rect -3609 -4262 -3575 -4238
rect -3517 -4238 -3483 -4228
rect -3517 -4262 -3483 -4238
rect -3425 -4238 -3391 -4228
rect -3425 -4262 -3391 -4238
rect -3333 -4238 -3299 -4228
rect -3333 -4262 -3299 -4238
rect -3241 -4238 -3207 -4228
rect -3241 -4262 -3207 -4238
rect -3149 -4238 -3115 -4228
rect -3149 -4262 -3115 -4238
rect -3057 -4238 -3023 -4228
rect -3057 -4262 -3023 -4238
rect -2965 -4238 -2931 -4228
rect -2965 -4262 -2931 -4238
rect -2873 -4238 -2839 -4228
rect -2873 -4262 -2839 -4238
rect -2781 -4238 -2747 -4228
rect -2781 -4262 -2747 -4238
rect -2689 -4238 -2655 -4228
rect -2689 -4262 -2655 -4238
rect -2597 -4238 -2563 -4228
rect -2597 -4262 -2563 -4238
rect -2505 -4238 -2471 -4228
rect -2505 -4262 -2471 -4238
rect -2413 -4238 -2379 -4228
rect -2413 -4262 -2379 -4238
rect -2321 -4238 -2287 -4228
rect -2321 -4262 -2287 -4238
rect -2229 -4238 -2195 -4228
rect -2229 -4262 -2195 -4238
rect -2137 -4238 -2103 -4228
rect -2137 -4262 -2103 -4238
rect -2045 -4238 -2011 -4228
rect -2045 -4262 -2011 -4238
rect -1953 -4238 -1919 -4228
rect -1953 -4262 -1919 -4238
rect -1861 -4238 -1827 -4228
rect -1861 -4262 -1827 -4238
rect -1769 -4238 -1735 -4228
rect -1769 -4262 -1735 -4238
rect -1677 -4238 -1643 -4228
rect -1677 -4262 -1643 -4238
rect -1585 -4238 -1551 -4228
rect -1585 -4262 -1551 -4238
rect -1493 -4238 -1459 -4228
rect -1493 -4262 -1459 -4238
rect -1401 -4238 -1367 -4228
rect -1401 -4262 -1367 -4238
rect -1309 -4238 -1275 -4228
rect -1309 -4262 -1275 -4238
rect -1217 -4238 -1183 -4228
rect -1217 -4262 -1183 -4238
rect -1125 -4238 -1091 -4228
rect -1125 -4262 -1091 -4238
rect -1033 -4238 -999 -4228
rect -1033 -4262 -999 -4238
rect -941 -4238 -907 -4228
rect -941 -4262 -907 -4238
rect -849 -4238 -815 -4228
rect -849 -4262 -815 -4238
rect -757 -4238 -723 -4228
rect -757 -4262 -723 -4238
rect -665 -4238 -631 -4228
rect -665 -4262 -631 -4238
rect -573 -4238 -539 -4228
rect -573 -4262 -539 -4238
rect -481 -4238 -447 -4228
rect -481 -4262 -447 -4238
rect -389 -4238 -355 -4228
rect -389 -4262 -355 -4238
rect -297 -4238 -263 -4228
rect -297 -4262 -263 -4238
rect -205 -4238 -171 -4228
rect -205 -4262 -171 -4238
rect -113 -4238 -79 -4228
rect -113 -4262 -79 -4238
rect -21 -4238 13 -4228
rect -21 -4262 13 -4238
rect 71 -4238 105 -4228
rect 71 -4262 105 -4238
rect 163 -4238 197 -4228
rect 163 -4262 197 -4238
rect 255 -4238 289 -4228
rect 255 -4262 289 -4238
rect 347 -4238 381 -4228
rect 347 -4262 381 -4238
rect 439 -4238 473 -4228
rect 439 -4262 473 -4238
rect 531 -4238 565 -4228
rect 531 -4262 565 -4238
rect 623 -4238 657 -4228
rect 623 -4262 657 -4238
rect 715 -4238 749 -4228
rect 715 -4262 749 -4238
rect 807 -4238 841 -4228
rect 807 -4262 841 -4238
rect 899 -4238 933 -4228
rect 899 -4262 933 -4238
rect 991 -4238 1025 -4228
rect 991 -4262 1025 -4238
rect 1083 -4238 1117 -4228
rect 1083 -4262 1117 -4238
rect 1175 -4238 1209 -4228
rect 1175 -4262 1209 -4238
rect 1267 -4238 1301 -4228
rect 1267 -4262 1301 -4238
rect 1359 -4238 1393 -4228
rect 1359 -4262 1393 -4238
rect 1451 -4238 1485 -4228
rect 1451 -4262 1485 -4238
rect 1543 -4238 1577 -4228
rect 1543 -4262 1577 -4238
rect 1635 -4238 1669 -4228
rect 1635 -4262 1669 -4238
rect 1727 -4238 1761 -4228
rect 1727 -4262 1761 -4238
rect 1819 -4238 1853 -4228
rect 1819 -4262 1853 -4238
rect 1911 -4238 1945 -4228
rect 1911 -4262 1945 -4238
rect 2003 -4238 2037 -4228
rect 2003 -4262 2037 -4238
rect 2095 -4238 2129 -4228
rect 2095 -4262 2129 -4238
rect 2187 -4238 2221 -4228
rect 2187 -4262 2221 -4238
rect 2279 -4238 2313 -4228
rect 2279 -4262 2313 -4238
rect 2371 -4238 2405 -4228
rect 2371 -4262 2405 -4238
rect 2463 -4238 2497 -4228
rect 2463 -4262 2497 -4238
rect 2555 -4238 2589 -4228
rect 2555 -4262 2589 -4238
rect 2647 -4238 2681 -4228
rect 2647 -4262 2681 -4238
rect 2739 -4238 2773 -4228
rect 2739 -4262 2773 -4238
rect 2831 -4238 2865 -4228
rect 2831 -4262 2865 -4238
rect 2923 -4238 2957 -4228
rect 2923 -4262 2957 -4238
rect 3015 -4238 3049 -4228
rect 3015 -4262 3049 -4238
rect 3107 -4238 3141 -4228
rect 3107 -4262 3141 -4238
rect 3199 -4238 3233 -4228
rect 3199 -4262 3233 -4238
rect 3291 -4238 3325 -4228
rect 3291 -4262 3325 -4238
rect 3383 -4238 3417 -4228
rect 3383 -4262 3417 -4238
rect 3475 -4238 3509 -4228
rect 3475 -4262 3509 -4238
rect 3567 -4238 3601 -4228
rect 3567 -4262 3601 -4238
rect 3659 -4238 3693 -4228
rect 3659 -4262 3693 -4238
rect 3751 -4238 3785 -4228
rect 3751 -4262 3785 -4238
rect 3843 -4238 3877 -4228
rect 3843 -4262 3877 -4238
rect 3935 -4238 3969 -4228
rect 3935 -4262 3969 -4238
rect 4027 -4238 4061 -4228
rect 4027 -4262 4061 -4238
rect 4119 -4238 4153 -4228
rect 4119 -4262 4153 -4238
rect 4211 -4238 4245 -4228
rect 4211 -4262 4245 -4238
rect 4303 -4238 4337 -4228
rect 4303 -4262 4337 -4238
rect 4395 -4238 4429 -4228
rect 4395 -4262 4429 -4238
rect 4487 -4238 4521 -4228
rect 4487 -4262 4521 -4238
rect 4579 -4238 4613 -4228
rect 4579 -4262 4613 -4238
rect 4671 -4238 4705 -4228
rect 4671 -4262 4705 -4238
rect 4763 -4238 4797 -4228
rect 4763 -4262 4797 -4238
rect 4855 -4238 4889 -4228
rect 4855 -4262 4889 -4238
rect 4947 -4238 4981 -4228
rect 4947 -4262 4981 -4238
rect 5039 -4238 5073 -4228
rect 5039 -4262 5073 -4238
rect 5131 -4238 5165 -4228
rect 5131 -4262 5165 -4238
rect 5223 -4238 5257 -4228
rect 5223 -4262 5257 -4238
rect 5315 -4238 5349 -4228
rect 5315 -4262 5349 -4238
rect 5407 -4238 5441 -4228
rect 5407 -4262 5441 -4238
rect 5499 -4238 5533 -4228
rect 5499 -4262 5533 -4238
rect 5591 -4238 5625 -4228
rect 5591 -4262 5625 -4238
rect 5683 -4238 5717 -4228
rect 5683 -4262 5717 -4238
rect 5775 -4238 5809 -4228
rect 5775 -4262 5809 -4238
rect 5867 -4238 5901 -4228
rect 5867 -4262 5901 -4238
rect 5959 -4238 5993 -4228
rect 5959 -4262 5993 -4238
rect 6051 -4238 6085 -4228
rect 6051 -4262 6085 -4238
rect 6143 -4238 6177 -4228
rect 6143 -4262 6177 -4238
rect 6235 -4238 6269 -4228
rect 6235 -4262 6269 -4238
rect 6327 -4238 6361 -4228
rect 6327 -4262 6361 -4238
rect 6419 -4238 6453 -4228
rect 6419 -4262 6453 -4238
rect 6511 -4238 6545 -4228
rect 6511 -4262 6545 -4238
rect 6603 -4238 6637 -4228
rect 6603 -4262 6637 -4238
rect 6695 -4238 6729 -4228
rect 6695 -4262 6729 -4238
rect 6787 -4238 6821 -4228
rect 6787 -4262 6821 -4238
rect 6879 -4238 6913 -4228
rect 6879 -4262 6913 -4238
rect 6971 -4238 7005 -4228
rect 6971 -4262 7005 -4238
rect 7063 -4238 7097 -4228
rect 7063 -4262 7097 -4238
rect 7155 -4238 7189 -4228
rect 7155 -4262 7189 -4238
rect 7247 -4238 7281 -4228
rect 7247 -4262 7281 -4238
rect 7339 -4238 7373 -4228
rect 7339 -4262 7373 -4238
rect 7431 -4238 7465 -4228
rect 7431 -4262 7465 -4238
rect 7523 -4238 7557 -4228
rect 7523 -4262 7557 -4238
rect 7615 -4238 7649 -4228
rect 7615 -4262 7649 -4238
rect 7707 -4238 7741 -4228
rect 7707 -4262 7741 -4238
rect 7799 -4238 7833 -4228
rect 7799 -4262 7833 -4238
rect 7891 -4238 7925 -4228
rect 7891 -4262 7925 -4238
rect 7983 -4238 8017 -4228
rect 7983 -4262 8017 -4238
rect 8075 -4238 8109 -4228
rect 8075 -4262 8109 -4238
rect 8167 -4238 8201 -4228
rect 8167 -4262 8201 -4238
rect 8259 -4238 8293 -4228
rect 8259 -4262 8293 -4238
rect 8351 -4238 8385 -4228
rect 8351 -4262 8385 -4238
rect 8443 -4238 8477 -4228
rect 8443 -4262 8477 -4238
rect 8535 -4238 8569 -4228
rect 8535 -4262 8569 -4238
rect 8627 -4238 8661 -4228
rect 8627 -4262 8661 -4238
rect 8719 -4238 8753 -4228
rect 8719 -4262 8753 -4238
rect 8811 -4238 8845 -4228
rect 8811 -4262 8845 -4238
rect 8903 -4238 8937 -4228
rect 8903 -4262 8937 -4238
rect 8995 -4238 9029 -4228
rect 8995 -4262 9029 -4238
rect 9087 -4238 9121 -4228
rect 9087 -4262 9121 -4238
rect 9179 -4238 9213 -4228
rect 9179 -4262 9213 -4238
rect 9271 -4238 9305 -4228
rect 9271 -4262 9305 -4238
rect 9363 -4238 9397 -4228
rect 9363 -4262 9397 -4238
rect 9455 -4238 9489 -4228
rect 9455 -4262 9489 -4238
rect 9547 -4238 9581 -4228
rect 9547 -4262 9581 -4238
rect 9639 -4238 9673 -4228
rect 9639 -4262 9673 -4238
rect 9731 -4238 9765 -4228
rect 9731 -4262 9765 -4238
rect 9823 -4238 9857 -4228
rect 9823 -4262 9857 -4238
rect 9915 -4238 9949 -4228
rect 9915 -4262 9949 -4238
rect 10007 -4238 10041 -4228
rect 10007 -4262 10041 -4238
rect 10099 -4238 10133 -4228
rect 10099 -4262 10133 -4238
rect 10191 -4238 10225 -4228
rect 10191 -4262 10225 -4238
rect 10283 -4238 10317 -4228
rect 10283 -4262 10317 -4238
rect 10375 -4238 10409 -4228
rect 10375 -4262 10409 -4238
rect 10467 -4238 10501 -4228
rect 10467 -4262 10501 -4238
rect 10559 -4238 10593 -4228
rect 10559 -4262 10593 -4238
rect 10651 -4238 10685 -4228
rect 10651 -4262 10685 -4238
rect 10743 -4238 10777 -4228
rect 10743 -4262 10777 -4238
rect 10835 -4238 10869 -4228
rect 10835 -4262 10869 -4238
rect 10927 -4238 10961 -4228
rect 10927 -4262 10961 -4238
rect 11019 -4238 11053 -4228
rect 11019 -4262 11053 -4238
rect 11111 -4238 11145 -4228
rect 11111 -4262 11145 -4238
rect 11203 -4238 11237 -4228
rect 11203 -4262 11237 -4238
rect 11295 -4238 11329 -4228
rect 11295 -4262 11329 -4238
rect 11387 -4238 11421 -4228
rect 11387 -4262 11421 -4238
rect 11479 -4238 11513 -4228
rect 11479 -4262 11513 -4238
rect 11571 -4238 11605 -4228
rect 11571 -4262 11605 -4238
rect 11663 -4238 11697 -4228
rect 11663 -4262 11697 -4238
rect 11755 -4238 11789 -4228
rect 11755 -4262 11789 -4238
rect 11847 -4238 11881 -4228
rect 11847 -4262 11881 -4238
rect 11939 -4238 11973 -4228
rect 11939 -4262 11973 -4238
rect 12031 -4238 12065 -4228
rect 12031 -4262 12065 -4238
rect 12123 -4238 12157 -4228
rect 12123 -4262 12157 -4238
rect 12215 -4238 12249 -4228
rect 12215 -4262 12249 -4238
rect 12307 -4238 12341 -4228
rect 12307 -4262 12341 -4238
rect 12399 -4238 12433 -4228
rect 12399 -4262 12433 -4238
rect 12491 -4238 12525 -4228
rect 12491 -4262 12525 -4238
rect 12583 -4238 12617 -4228
rect 12583 -4262 12617 -4238
rect 12675 -4238 12709 -4228
rect 12675 -4262 12709 -4238
rect 12767 -4238 12801 -4228
rect 12767 -4262 12801 -4238
rect 12859 -4238 12893 -4228
rect 12859 -4262 12893 -4238
rect 12951 -4238 12985 -4228
rect 12951 -4262 12985 -4238
rect 13043 -4238 13077 -4228
rect 13043 -4262 13077 -4238
rect 13135 -4238 13169 -4228
rect 13135 -4262 13169 -4238
rect 13227 -4238 13261 -4228
rect 13227 -4262 13261 -4238
rect 13319 -4238 13353 -4228
rect 13319 -4262 13353 -4238
rect 13411 -4238 13445 -4228
rect 13411 -4262 13445 -4238
rect 13503 -4238 13537 -4228
rect 13503 -4262 13537 -4238
rect 13595 -4238 13629 -4228
rect 13595 -4262 13629 -4238
rect 13687 -4238 13721 -4228
rect 13687 -4262 13721 -4238
rect 13779 -4238 13813 -4228
rect 13779 -4262 13813 -4238
rect 13871 -4238 13905 -4228
rect 13871 -4262 13905 -4238
rect 13963 -4238 13997 -4228
rect 13963 -4262 13997 -4238
rect 14055 -4238 14089 -4228
rect 14055 -4262 14089 -4238
rect 14147 -4238 14181 -4228
rect 14147 -4262 14181 -4238
rect 14239 -4238 14273 -4228
rect 14239 -4262 14273 -4238
rect 14331 -4238 14365 -4228
rect 14331 -4262 14365 -4238
rect 14423 -4238 14457 -4228
rect 14423 -4262 14457 -4238
rect 14515 -4238 14549 -4228
rect 14515 -4262 14549 -4238
rect 14607 -4238 14641 -4228
rect 14607 -4262 14641 -4238
rect 14699 -4238 14733 -4228
rect 14699 -4262 14733 -4238
rect 14791 -4238 14825 -4228
rect 14791 -4262 14825 -4238
rect 14883 -4238 14917 -4228
rect 14883 -4262 14917 -4238
rect 14975 -4238 15009 -4228
rect 14975 -4262 15009 -4238
rect 15067 -4238 15101 -4228
rect 15067 -4262 15101 -4238
rect 15159 -4238 15193 -4228
rect 15159 -4262 15193 -4238
rect 15251 -4238 15285 -4228
rect 15251 -4262 15285 -4238
rect 15343 -4238 15377 -4228
rect 15343 -4262 15377 -4238
rect 15435 -4238 15469 -4228
rect 15435 -4262 15469 -4238
rect 15527 -4238 15561 -4228
rect 15527 -4262 15561 -4238
rect 15619 -4238 15653 -4228
rect 15619 -4262 15653 -4238
rect 15711 -4238 15745 -4228
rect 15711 -4262 15745 -4238
rect 15803 -4238 15837 -4228
rect 15803 -4262 15837 -4238
rect 15895 -4238 15929 -4228
rect 15895 -4262 15929 -4238
rect 15987 -4238 16021 -4228
rect 15987 -4262 16021 -4238
rect 16079 -4238 16113 -4228
rect 16079 -4262 16113 -4238
rect 16171 -4238 16205 -4228
rect 16171 -4262 16205 -4238
rect 16263 -4238 16297 -4228
rect 16263 -4262 16297 -4238
rect 16355 -4238 16389 -4228
rect 16355 -4262 16389 -4238
rect 16447 -4238 16481 -4228
rect 16447 -4262 16481 -4238
rect 16539 -4238 16573 -4228
rect 16539 -4262 16573 -4238
rect 16631 -4238 16665 -4228
rect 16631 -4262 16665 -4238
rect 16723 -4238 16757 -4228
rect 16723 -4262 16757 -4238
rect 16815 -4238 16849 -4228
rect 16815 -4262 16849 -4238
rect 16907 -4238 16941 -4228
rect 16907 -4262 16941 -4238
rect 16999 -4238 17033 -4228
rect 16999 -4262 17033 -4238
rect 17091 -4238 17125 -4228
rect 17091 -4262 17125 -4238
rect 17183 -4238 17217 -4228
rect 17183 -4262 17217 -4238
rect 17275 -4238 17309 -4228
rect 17275 -4262 17309 -4238
rect 17367 -4238 17401 -4228
rect 17367 -4262 17401 -4238
rect 17459 -4238 17493 -4228
rect 17459 -4262 17493 -4238
rect 17551 -4238 17585 -4228
rect 17551 -4262 17585 -4238
rect 17643 -4238 17677 -4228
rect 17643 -4262 17677 -4238
rect 17735 -4238 17769 -4228
rect 17735 -4262 17769 -4238
rect 17827 -4238 17861 -4228
rect 17827 -4262 17861 -4238
rect 17919 -4238 17953 -4228
rect 17919 -4262 17953 -4238
rect 18011 -4238 18045 -4228
rect 18011 -4262 18045 -4238
rect 18103 -4238 18137 -4228
rect 18103 -4262 18137 -4238
rect 18195 -4238 18229 -4228
rect 18195 -4262 18229 -4238
rect 18287 -4238 18321 -4228
rect 18287 -4262 18321 -4238
rect 18379 -4238 18413 -4228
rect 18379 -4262 18413 -4238
rect 18471 -4238 18505 -4228
rect 18471 -4262 18505 -4238
rect 18563 -4238 18597 -4228
rect 18563 -4262 18597 -4238
rect 18655 -4238 18689 -4228
rect 18655 -4262 18689 -4238
rect 18747 -4238 18781 -4228
rect 18747 -4262 18781 -4238
rect 18839 -4238 18873 -4228
rect 18839 -4262 18873 -4238
rect 18931 -4238 18965 -4228
rect 18931 -4262 18965 -4238
rect 19023 -4238 19057 -4228
rect 19023 -4262 19057 -4238
rect 19115 -4238 19149 -4228
rect 19115 -4262 19149 -4238
rect 19207 -4238 19241 -4228
rect 19207 -4262 19241 -4238
rect 19299 -4238 19333 -4228
rect 19299 -4262 19333 -4238
rect 19391 -4238 19425 -4228
rect 19391 -4262 19425 -4238
rect 19483 -4238 19517 -4228
rect 19483 -4262 19517 -4238
rect 19575 -4238 19609 -4228
rect 19575 -4262 19609 -4238
rect 19667 -4238 19701 -4228
rect 19667 -4262 19701 -4238
rect 19759 -4238 19793 -4228
rect 19759 -4262 19793 -4238
rect 19851 -4238 19885 -4228
rect 19851 -4262 19885 -4238
rect 19943 -4238 19977 -4228
rect 19943 -4262 19977 -4238
rect 20035 -4238 20069 -4228
rect 20035 -4262 20069 -4238
rect 20127 -4238 20161 -4228
rect 20127 -4262 20161 -4238
rect 20219 -4238 20253 -4228
rect 20219 -4262 20253 -4238
rect 20311 -4238 20345 -4228
rect 20311 -4262 20345 -4238
rect 20403 -4238 20437 -4228
rect 20403 -4262 20437 -4238
rect 20495 -4238 20529 -4228
rect 20495 -4262 20529 -4238
rect 20587 -4238 20621 -4228
rect 20587 -4262 20621 -4238
rect 20679 -4238 20713 -4228
rect 20679 -4262 20713 -4238
rect 20771 -4238 20805 -4228
rect 20771 -4262 20805 -4238
rect 20863 -4238 20897 -4228
rect 20863 -4262 20897 -4238
rect 20955 -4238 20989 -4228
rect 20955 -4262 20989 -4238
rect 21047 -4238 21081 -4228
rect 21047 -4262 21081 -4238
rect 21139 -4238 21173 -4228
rect 21139 -4262 21173 -4238
rect 21231 -4238 21265 -4228
rect 21231 -4262 21265 -4238
rect 21323 -4238 21357 -4228
rect 21323 -4262 21357 -4238
rect 21415 -4238 21449 -4228
rect 21415 -4262 21449 -4238
rect 21507 -4238 21541 -4228
rect 21507 -4262 21541 -4238
rect 21599 -4238 21633 -4228
rect 21599 -4262 21633 -4238
rect 21691 -4238 21725 -4228
rect 21691 -4262 21725 -4238
rect 21783 -4238 21817 -4228
rect 21783 -4262 21817 -4238
rect 21875 -4238 21909 -4228
rect 21875 -4262 21909 -4238
rect 21967 -4238 22001 -4228
rect 21967 -4262 22001 -4238
rect 22059 -4238 22093 -4228
rect 22059 -4262 22093 -4238
rect 22151 -4238 22185 -4228
rect 22151 -4262 22185 -4238
rect 22243 -4238 22277 -4228
rect 22243 -4262 22277 -4238
rect 22335 -4238 22369 -4228
rect 22335 -4262 22369 -4238
rect 22427 -4238 22461 -4228
rect 22427 -4262 22461 -4238
rect 22519 -4238 22553 -4228
rect 22519 -4262 22553 -4238
rect 22611 -4238 22645 -4228
rect 22611 -4262 22645 -4238
rect 22703 -4238 22737 -4228
rect 22703 -4262 22737 -4238
rect 22795 -4238 22829 -4228
rect 22795 -4262 22829 -4238
rect 22887 -4238 22921 -4228
rect 22887 -4262 22921 -4238
rect 22979 -4238 23013 -4228
rect 22979 -4262 23013 -4238
rect 23071 -4238 23105 -4228
rect 23071 -4262 23105 -4238
rect 23163 -4238 23197 -4228
rect 23163 -4262 23197 -4238
rect 23255 -4238 23289 -4228
rect 23255 -4262 23289 -4238
rect 23347 -4238 23381 -4228
rect 23347 -4262 23381 -4238
rect 23439 -4238 23473 -4228
rect 23439 -4262 23473 -4238
rect 23531 -4238 23565 -4228
rect 23531 -4262 23565 -4238
rect 23623 -4238 23657 -4228
rect 23623 -4262 23657 -4238
rect 23715 -4238 23749 -4228
rect 23715 -4262 23749 -4238
rect 23807 -4238 23841 -4228
rect 23807 -4262 23841 -4238
rect 23899 -4238 23933 -4228
rect 23899 -4262 23933 -4238
rect 23991 -4238 24025 -4228
rect 23991 -4262 24025 -4238
rect 24083 -4238 24117 -4228
rect 24083 -4262 24117 -4238
rect 24175 -4238 24209 -4228
rect 24175 -4262 24209 -4238
rect 24267 -4238 24301 -4228
rect 24267 -4262 24301 -4238
rect 24359 -4238 24393 -4228
rect 24359 -4262 24393 -4238
rect 24451 -4238 24485 -4228
rect 24451 -4262 24485 -4238
rect 24543 -4238 24577 -4228
rect 24543 -4262 24577 -4238
rect 24635 -4238 24669 -4228
rect 24635 -4262 24669 -4238
rect 24727 -4238 24761 -4228
rect 24727 -4262 24761 -4238
rect 24819 -4238 24853 -4228
rect 24819 -4262 24853 -4238
rect 24911 -4238 24945 -4228
rect 24911 -4262 24945 -4238
rect 25003 -4238 25037 -4228
rect 25003 -4262 25037 -4238
rect 25095 -4238 25129 -4228
rect 25095 -4262 25129 -4238
rect 25187 -4238 25221 -4228
rect 25187 -4262 25221 -4238
rect 25279 -4238 25313 -4228
rect 25279 -4262 25313 -4238
rect 25371 -4238 25405 -4228
rect 25371 -4262 25405 -4238
rect 25463 -4238 25497 -4228
rect 25463 -4262 25497 -4238
rect 25555 -4238 25589 -4228
rect 25555 -4262 25589 -4238
rect 25647 -4238 25681 -4228
rect 25647 -4262 25681 -4238
rect 25739 -4238 25773 -4228
rect 25739 -4262 25773 -4238
rect 25831 -4238 25865 -4228
rect 25831 -4262 25865 -4238
rect 25923 -4238 25957 -4228
rect 25923 -4262 25957 -4238
rect 26015 -4238 26049 -4228
rect 26015 -4262 26049 -4238
rect 26107 -4238 26141 -4228
rect 26107 -4262 26141 -4238
rect 26199 -4238 26233 -4228
rect 26199 -4262 26233 -4238
rect 26291 -4238 26325 -4228
rect 26291 -4262 26325 -4238
rect 26383 -4238 26417 -4228
rect 26383 -4262 26417 -4238
rect 26475 -4238 26509 -4228
rect 26475 -4262 26509 -4238
rect 26567 -4238 26601 -4228
rect 26567 -4262 26601 -4238
rect 26659 -4238 26693 -4228
rect 26659 -4262 26693 -4238
rect 26751 -4238 26785 -4228
rect 26751 -4262 26785 -4238
rect 26843 -4238 26877 -4228
rect 26843 -4262 26877 -4238
rect 26935 -4238 26969 -4228
rect 26935 -4262 26969 -4238
rect 27027 -4238 27061 -4228
rect 27027 -4262 27061 -4238
rect 27119 -4238 27153 -4228
rect 27119 -4262 27153 -4238
rect 27211 -4238 27245 -4228
rect 27211 -4262 27245 -4238
rect 27303 -4238 27337 -4228
rect 27303 -4262 27337 -4238
rect 27395 -4238 27429 -4228
rect 27395 -4262 27429 -4238
rect 27487 -4238 27521 -4228
rect 27487 -4262 27521 -4238
rect 27579 -4238 27613 -4228
rect 27579 -4262 27613 -4238
rect 27671 -4238 27705 -4228
rect 27671 -4262 27705 -4238
rect 27763 -4238 27797 -4228
rect 27763 -4262 27797 -4238
rect 27855 -4238 27889 -4228
rect 27855 -4262 27889 -4238
rect 27947 -4238 27981 -4228
rect 27947 -4262 27981 -4238
rect 28039 -4238 28073 -4228
rect 28039 -4262 28073 -4238
rect 28131 -4238 28165 -4228
rect 28131 -4262 28165 -4238
rect 28223 -4238 28257 -4228
rect 28223 -4262 28257 -4238
rect 28315 -4238 28349 -4228
rect 28315 -4262 28349 -4238
rect 28407 -4238 28441 -4228
rect 28407 -4262 28441 -4238
rect 28499 -4238 28533 -4228
rect 28499 -4262 28533 -4238
rect 28591 -4238 28625 -4228
rect 28591 -4262 28625 -4238
rect 28683 -4238 28717 -4228
rect 28683 -4262 28717 -4238
rect 28775 -4238 28809 -4228
rect 28775 -4262 28809 -4238
rect 28867 -4238 28901 -4228
rect 28867 -4262 28901 -4238
rect 28959 -4238 28993 -4228
rect 28959 -4262 28993 -4238
rect 29051 -4238 29085 -4228
rect 29051 -4262 29085 -4238
rect 29143 -4238 29177 -4228
rect 29143 -4262 29177 -4238
rect 29235 -4238 29269 -4228
rect 29235 -4262 29269 -4238
rect 29327 -4238 29361 -4228
rect 29327 -4262 29361 -4238
rect 29419 -4238 29453 -4228
rect 29419 -4262 29453 -4238
rect 29511 -4238 29545 -4228
rect 29511 -4262 29545 -4238
rect 29603 -4238 29637 -4228
rect 29603 -4262 29637 -4238
rect 29695 -4238 29729 -4228
rect 29695 -4262 29729 -4238
rect 29787 -4238 29821 -4228
rect 29787 -4262 29821 -4238
rect 29879 -4238 29913 -4228
rect 29879 -4262 29913 -4238
rect 29971 -4238 30005 -4228
rect 29971 -4262 30005 -4238
rect 30063 -4238 30097 -4228
rect 30063 -4262 30097 -4238
rect 30155 -4238 30189 -4228
rect 30155 -4262 30189 -4238
rect 30247 -4238 30281 -4228
rect 30247 -4262 30281 -4238
rect 30339 -4238 30373 -4228
rect 30339 -4262 30373 -4238
rect 30431 -4238 30465 -4228
rect 30431 -4262 30465 -4238
rect 30523 -4238 30557 -4228
rect 30523 -4262 30557 -4238
rect 30615 -4238 30649 -4228
rect 30615 -4262 30649 -4238
rect 30707 -4238 30741 -4228
rect 30707 -4262 30741 -4238
rect 30799 -4238 30833 -4228
rect 30799 -4262 30833 -4238
rect 30891 -4238 30925 -4228
rect 30891 -4262 30925 -4238
rect 30983 -4238 31017 -4228
rect 30983 -4262 31017 -4238
rect 31075 -4238 31109 -4228
rect 31075 -4262 31109 -4238
rect 31167 -4238 31201 -4228
rect 31167 -4262 31201 -4238
rect 31259 -4238 31293 -4228
rect 31259 -4262 31293 -4238
rect 31351 -4238 31385 -4228
rect 31351 -4262 31385 -4238
rect 31443 -4238 31477 -4228
rect 31443 -4262 31477 -4238
rect 31535 -4238 31569 -4228
rect 31535 -4262 31569 -4238
rect 31627 -4238 31661 -4228
rect 31627 -4262 31661 -4238
rect 31719 -4238 31753 -4228
rect 31719 -4262 31753 -4238
rect 31811 -4238 31845 -4228
rect 31811 -4262 31845 -4238
rect 31903 -4238 31937 -4228
rect 31903 -4262 31937 -4238
rect 31995 -4238 32029 -4228
rect 31995 -4262 32029 -4238
rect 32087 -4238 32121 -4228
rect 32087 -4262 32121 -4238
rect 32179 -4238 32213 -4228
rect 32179 -4262 32213 -4238
rect 32271 -4238 32305 -4228
rect 32271 -4262 32305 -4238
rect 32363 -4238 32397 -4228
rect 32363 -4262 32397 -4238
rect 32455 -4238 32489 -4228
rect 32455 -4262 32489 -4238
rect 32547 -4238 32581 -4228
rect 32547 -4262 32581 -4238
rect 32639 -4238 32673 -4228
rect 32639 -4262 32673 -4238
rect 32731 -4238 32765 -4228
rect 32731 -4262 32765 -4238
rect 32823 -4238 32857 -4228
rect 32823 -4262 32857 -4238
rect 32915 -4238 32949 -4228
rect 32915 -4262 32949 -4238
rect 33007 -4238 33041 -4228
rect 33007 -4262 33041 -4238
rect 33099 -4238 33133 -4228
rect 33099 -4262 33133 -4238
rect -9036 -4559 -9024 -4534
rect -9024 -4559 -9002 -4534
rect -9036 -4568 -9002 -4559
rect -8955 -4414 -8921 -4398
rect -8955 -4432 -8921 -4414
rect -8851 -4648 -8813 -4614
rect -8577 -4432 -8543 -4398
rect -8669 -4568 -8635 -4534
rect -7953 -4424 -7919 -4398
rect -7953 -4432 -7922 -4424
rect -7922 -4432 -7919 -4424
rect -8397 -4636 -8363 -4602
rect -8325 -4620 -8301 -4602
rect -8301 -4620 -8291 -4602
rect -8325 -4636 -8291 -4620
rect -7953 -4550 -7919 -4534
rect -7953 -4568 -7927 -4550
rect -7927 -4568 -7919 -4550
rect -7737 -4548 -7703 -4539
rect -7737 -4573 -7721 -4548
rect -7721 -4573 -7703 -4548
rect -7677 -4636 -7643 -4602
rect -7082 -4549 -7044 -4515
rect -6920 -4559 -6908 -4534
rect -6908 -4559 -6886 -4534
rect -6920 -4568 -6886 -4559
rect -6839 -4414 -6805 -4398
rect -6839 -4432 -6805 -4414
rect -6735 -4648 -6697 -4614
rect -6461 -4432 -6427 -4398
rect -6553 -4568 -6519 -4534
rect -5837 -4424 -5803 -4398
rect -5837 -4432 -5806 -4424
rect -5806 -4432 -5803 -4424
rect -6281 -4636 -6247 -4602
rect -6209 -4620 -6185 -4602
rect -6185 -4620 -6175 -4602
rect -6209 -4636 -6175 -4620
rect -5837 -4550 -5803 -4534
rect -5837 -4568 -5811 -4550
rect -5811 -4568 -5803 -4550
rect -5621 -4548 -5587 -4539
rect -5621 -4573 -5605 -4548
rect -5605 -4573 -5587 -4548
rect -5561 -4636 -5527 -4602
rect -4966 -4549 -4928 -4515
rect -4804 -4559 -4792 -4534
rect -4792 -4559 -4770 -4534
rect -4804 -4568 -4770 -4559
rect -4723 -4414 -4689 -4398
rect -4723 -4432 -4689 -4414
rect -4619 -4648 -4581 -4614
rect -4345 -4432 -4311 -4398
rect -4437 -4568 -4403 -4534
rect -3721 -4424 -3687 -4398
rect -3721 -4432 -3690 -4424
rect -3690 -4432 -3687 -4424
rect -4165 -4636 -4131 -4602
rect -4093 -4620 -4069 -4602
rect -4069 -4620 -4059 -4602
rect -4093 -4636 -4059 -4620
rect -3721 -4550 -3687 -4534
rect -3721 -4568 -3695 -4550
rect -3695 -4568 -3687 -4550
rect -3505 -4548 -3471 -4539
rect -3505 -4573 -3489 -4548
rect -3489 -4573 -3471 -4548
rect -3445 -4636 -3411 -4602
rect -2850 -4549 -2812 -4515
rect -2688 -4559 -2676 -4534
rect -2676 -4559 -2654 -4534
rect -2688 -4568 -2654 -4559
rect -2607 -4414 -2573 -4398
rect -2607 -4432 -2573 -4414
rect -2503 -4648 -2465 -4614
rect -2229 -4432 -2195 -4398
rect -2321 -4568 -2287 -4534
rect -1605 -4424 -1571 -4398
rect -1605 -4432 -1574 -4424
rect -1574 -4432 -1571 -4424
rect -2049 -4636 -2015 -4602
rect -1977 -4620 -1953 -4602
rect -1953 -4620 -1943 -4602
rect -1977 -4636 -1943 -4620
rect -1605 -4550 -1571 -4534
rect -1605 -4568 -1579 -4550
rect -1579 -4568 -1571 -4550
rect -1389 -4548 -1355 -4539
rect -1389 -4573 -1373 -4548
rect -1373 -4573 -1355 -4548
rect -1329 -4636 -1295 -4602
rect -734 -4549 -696 -4515
rect -572 -4559 -560 -4534
rect -560 -4559 -538 -4534
rect -572 -4568 -538 -4559
rect -491 -4414 -457 -4398
rect -491 -4432 -457 -4414
rect -387 -4648 -349 -4614
rect -113 -4432 -79 -4398
rect -205 -4568 -171 -4534
rect 511 -4424 545 -4398
rect 511 -4432 542 -4424
rect 542 -4432 545 -4424
rect 67 -4636 101 -4602
rect 139 -4620 163 -4602
rect 163 -4620 173 -4602
rect 139 -4636 173 -4620
rect 511 -4550 545 -4534
rect 511 -4568 537 -4550
rect 537 -4568 545 -4550
rect 727 -4548 761 -4539
rect 727 -4573 743 -4548
rect 743 -4573 761 -4548
rect 787 -4636 821 -4602
rect 1382 -4549 1420 -4515
rect 1544 -4559 1556 -4534
rect 1556 -4559 1578 -4534
rect 1544 -4568 1578 -4559
rect 1625 -4414 1659 -4398
rect 1625 -4432 1659 -4414
rect 1729 -4648 1767 -4614
rect 2003 -4432 2037 -4398
rect 1911 -4568 1945 -4534
rect 2627 -4424 2661 -4398
rect 2627 -4432 2658 -4424
rect 2658 -4432 2661 -4424
rect 2183 -4636 2217 -4602
rect 2255 -4620 2279 -4602
rect 2279 -4620 2289 -4602
rect 2255 -4636 2289 -4620
rect 2627 -4550 2661 -4534
rect 2627 -4568 2653 -4550
rect 2653 -4568 2661 -4550
rect 2843 -4548 2877 -4539
rect 2843 -4573 2859 -4548
rect 2859 -4573 2877 -4548
rect 2903 -4636 2937 -4602
rect 3498 -4549 3536 -4515
rect 3660 -4559 3672 -4534
rect 3672 -4559 3694 -4534
rect 3660 -4568 3694 -4559
rect 3741 -4414 3775 -4398
rect 3741 -4432 3775 -4414
rect 3845 -4648 3883 -4614
rect 4119 -4432 4153 -4398
rect 4027 -4568 4061 -4534
rect 4743 -4424 4777 -4398
rect 4743 -4432 4774 -4424
rect 4774 -4432 4777 -4424
rect 4299 -4636 4333 -4602
rect 4371 -4620 4395 -4602
rect 4395 -4620 4405 -4602
rect 4371 -4636 4405 -4620
rect 4743 -4550 4777 -4534
rect 4743 -4568 4769 -4550
rect 4769 -4568 4777 -4550
rect 4959 -4548 4993 -4539
rect 4959 -4573 4975 -4548
rect 4975 -4573 4993 -4548
rect 5019 -4636 5053 -4602
rect 5614 -4549 5652 -4515
rect 5776 -4559 5788 -4534
rect 5788 -4559 5810 -4534
rect 5776 -4568 5810 -4559
rect 5857 -4414 5891 -4398
rect 5857 -4432 5891 -4414
rect 5961 -4648 5999 -4614
rect 6235 -4432 6269 -4398
rect 6143 -4568 6177 -4534
rect 6859 -4424 6893 -4398
rect 6859 -4432 6890 -4424
rect 6890 -4432 6893 -4424
rect 6415 -4636 6449 -4602
rect 6487 -4620 6511 -4602
rect 6511 -4620 6521 -4602
rect 6487 -4636 6521 -4620
rect 6859 -4550 6893 -4534
rect 6859 -4568 6885 -4550
rect 6885 -4568 6893 -4550
rect 7075 -4548 7109 -4539
rect 7075 -4573 7091 -4548
rect 7091 -4573 7109 -4548
rect 7135 -4636 7169 -4602
rect 7730 -4549 7768 -4515
rect 7892 -4559 7904 -4534
rect 7904 -4559 7926 -4534
rect 7892 -4568 7926 -4559
rect 7973 -4414 8007 -4398
rect 7973 -4432 8007 -4414
rect 8077 -4648 8115 -4614
rect 8351 -4432 8385 -4398
rect 8259 -4568 8293 -4534
rect 8975 -4424 9009 -4398
rect 8975 -4432 9006 -4424
rect 9006 -4432 9009 -4424
rect 8531 -4636 8565 -4602
rect 8603 -4620 8627 -4602
rect 8627 -4620 8637 -4602
rect 8603 -4636 8637 -4620
rect 8975 -4550 9009 -4534
rect 8975 -4568 9001 -4550
rect 9001 -4568 9009 -4550
rect 9191 -4548 9225 -4539
rect 9191 -4573 9207 -4548
rect 9207 -4573 9225 -4548
rect 9251 -4636 9285 -4602
rect 9846 -4549 9884 -4515
rect 10008 -4559 10020 -4534
rect 10020 -4559 10042 -4534
rect 10008 -4568 10042 -4559
rect 10089 -4414 10123 -4398
rect 10089 -4432 10123 -4414
rect 10193 -4648 10231 -4614
rect 10467 -4432 10501 -4398
rect 10375 -4568 10409 -4534
rect 11091 -4424 11125 -4398
rect 11091 -4432 11122 -4424
rect 11122 -4432 11125 -4424
rect 10647 -4636 10681 -4602
rect 10719 -4620 10743 -4602
rect 10743 -4620 10753 -4602
rect 10719 -4636 10753 -4620
rect 11091 -4550 11125 -4534
rect 11091 -4568 11117 -4550
rect 11117 -4568 11125 -4550
rect 11307 -4548 11341 -4539
rect 11307 -4573 11323 -4548
rect 11323 -4573 11341 -4548
rect 11367 -4636 11401 -4602
rect 11962 -4549 12000 -4515
rect 12124 -4559 12136 -4534
rect 12136 -4559 12158 -4534
rect 12124 -4568 12158 -4559
rect 12205 -4414 12239 -4398
rect 12205 -4432 12239 -4414
rect 12309 -4648 12347 -4614
rect 12583 -4432 12617 -4398
rect 12491 -4568 12525 -4534
rect 13207 -4424 13241 -4398
rect 13207 -4432 13238 -4424
rect 13238 -4432 13241 -4424
rect 12763 -4636 12797 -4602
rect 12835 -4620 12859 -4602
rect 12859 -4620 12869 -4602
rect 12835 -4636 12869 -4620
rect 13207 -4550 13241 -4534
rect 13207 -4568 13233 -4550
rect 13233 -4568 13241 -4550
rect 13423 -4548 13457 -4539
rect 13423 -4573 13439 -4548
rect 13439 -4573 13457 -4548
rect 13483 -4636 13517 -4602
rect 14078 -4549 14116 -4515
rect 14240 -4559 14252 -4534
rect 14252 -4559 14274 -4534
rect 14240 -4568 14274 -4559
rect 14321 -4414 14355 -4398
rect 14321 -4432 14355 -4414
rect 14425 -4648 14463 -4614
rect 14699 -4432 14733 -4398
rect 14607 -4568 14641 -4534
rect 15323 -4424 15357 -4398
rect 15323 -4432 15354 -4424
rect 15354 -4432 15357 -4424
rect 14879 -4636 14913 -4602
rect 14951 -4620 14975 -4602
rect 14975 -4620 14985 -4602
rect 14951 -4636 14985 -4620
rect 15323 -4550 15357 -4534
rect 15323 -4568 15349 -4550
rect 15349 -4568 15357 -4550
rect 15539 -4548 15573 -4539
rect 15539 -4573 15555 -4548
rect 15555 -4573 15573 -4548
rect 15599 -4636 15633 -4602
rect 16194 -4549 16232 -4515
rect 16356 -4559 16368 -4534
rect 16368 -4559 16390 -4534
rect 16356 -4568 16390 -4559
rect 16437 -4414 16471 -4398
rect 16437 -4432 16471 -4414
rect 16541 -4648 16579 -4614
rect 16815 -4432 16849 -4398
rect 16723 -4568 16757 -4534
rect 17439 -4424 17473 -4398
rect 17439 -4432 17470 -4424
rect 17470 -4432 17473 -4424
rect 16995 -4636 17029 -4602
rect 17067 -4620 17091 -4602
rect 17091 -4620 17101 -4602
rect 17067 -4636 17101 -4620
rect 17439 -4550 17473 -4534
rect 17439 -4568 17465 -4550
rect 17465 -4568 17473 -4550
rect 17655 -4548 17689 -4539
rect 17655 -4573 17671 -4548
rect 17671 -4573 17689 -4548
rect 17715 -4636 17749 -4602
rect 18310 -4549 18348 -4515
rect 18472 -4559 18484 -4534
rect 18484 -4559 18506 -4534
rect 18472 -4568 18506 -4559
rect 18553 -4414 18587 -4398
rect 18553 -4432 18587 -4414
rect 18657 -4648 18695 -4614
rect 18931 -4432 18965 -4398
rect 18839 -4568 18873 -4534
rect 19555 -4424 19589 -4398
rect 19555 -4432 19586 -4424
rect 19586 -4432 19589 -4424
rect 19111 -4636 19145 -4602
rect 19183 -4620 19207 -4602
rect 19207 -4620 19217 -4602
rect 19183 -4636 19217 -4620
rect 19555 -4550 19589 -4534
rect 19555 -4568 19581 -4550
rect 19581 -4568 19589 -4550
rect 19771 -4548 19805 -4539
rect 19771 -4573 19787 -4548
rect 19787 -4573 19805 -4548
rect 19831 -4636 19865 -4602
rect 20426 -4549 20464 -4515
rect 20588 -4559 20600 -4534
rect 20600 -4559 20622 -4534
rect 20588 -4568 20622 -4559
rect 20669 -4414 20703 -4398
rect 20669 -4432 20703 -4414
rect 20773 -4648 20811 -4614
rect 21047 -4432 21081 -4398
rect 20955 -4568 20989 -4534
rect 21671 -4424 21705 -4398
rect 21671 -4432 21702 -4424
rect 21702 -4432 21705 -4424
rect 21227 -4636 21261 -4602
rect 21299 -4620 21323 -4602
rect 21323 -4620 21333 -4602
rect 21299 -4636 21333 -4620
rect 21671 -4550 21705 -4534
rect 21671 -4568 21697 -4550
rect 21697 -4568 21705 -4550
rect 21887 -4548 21921 -4539
rect 21887 -4573 21903 -4548
rect 21903 -4573 21921 -4548
rect 21947 -4636 21981 -4602
rect 22542 -4549 22580 -4515
rect 22704 -4559 22716 -4534
rect 22716 -4559 22738 -4534
rect 22704 -4568 22738 -4559
rect 22785 -4414 22819 -4398
rect 22785 -4432 22819 -4414
rect 22889 -4648 22927 -4614
rect 23163 -4432 23197 -4398
rect 23071 -4568 23105 -4534
rect 23787 -4424 23821 -4398
rect 23787 -4432 23818 -4424
rect 23818 -4432 23821 -4424
rect 23343 -4636 23377 -4602
rect 23415 -4620 23439 -4602
rect 23439 -4620 23449 -4602
rect 23415 -4636 23449 -4620
rect 23787 -4550 23821 -4534
rect 23787 -4568 23813 -4550
rect 23813 -4568 23821 -4550
rect 24003 -4548 24037 -4539
rect 24003 -4573 24019 -4548
rect 24019 -4573 24037 -4548
rect 24063 -4636 24097 -4602
rect 24658 -4549 24696 -4515
rect 24820 -4559 24832 -4534
rect 24832 -4559 24854 -4534
rect 24820 -4568 24854 -4559
rect 24901 -4414 24935 -4398
rect 24901 -4432 24935 -4414
rect 25005 -4648 25043 -4614
rect 25279 -4432 25313 -4398
rect 25187 -4568 25221 -4534
rect 25903 -4424 25937 -4398
rect 25903 -4432 25934 -4424
rect 25934 -4432 25937 -4424
rect 25459 -4636 25493 -4602
rect 25531 -4620 25555 -4602
rect 25555 -4620 25565 -4602
rect 25531 -4636 25565 -4620
rect 25903 -4550 25937 -4534
rect 25903 -4568 25929 -4550
rect 25929 -4568 25937 -4550
rect 26119 -4548 26153 -4539
rect 26119 -4573 26135 -4548
rect 26135 -4573 26153 -4548
rect 26179 -4636 26213 -4602
rect 26774 -4549 26812 -4515
rect 26936 -4559 26948 -4534
rect 26948 -4559 26970 -4534
rect 26936 -4568 26970 -4559
rect 27017 -4414 27051 -4398
rect 27017 -4432 27051 -4414
rect 27121 -4648 27159 -4614
rect 27395 -4432 27429 -4398
rect 27303 -4568 27337 -4534
rect 28019 -4424 28053 -4398
rect 28019 -4432 28050 -4424
rect 28050 -4432 28053 -4424
rect 27575 -4636 27609 -4602
rect 27647 -4620 27671 -4602
rect 27671 -4620 27681 -4602
rect 27647 -4636 27681 -4620
rect 28019 -4550 28053 -4534
rect 28019 -4568 28045 -4550
rect 28045 -4568 28053 -4550
rect 28235 -4548 28269 -4539
rect 28235 -4573 28251 -4548
rect 28251 -4573 28269 -4548
rect 28295 -4636 28329 -4602
rect 28890 -4549 28928 -4515
rect 29052 -4559 29064 -4534
rect 29064 -4559 29086 -4534
rect 29052 -4568 29086 -4559
rect 29133 -4414 29167 -4398
rect 29133 -4432 29167 -4414
rect 29237 -4648 29275 -4614
rect 29511 -4432 29545 -4398
rect 29419 -4568 29453 -4534
rect 30135 -4424 30169 -4398
rect 30135 -4432 30166 -4424
rect 30166 -4432 30169 -4424
rect 29691 -4636 29725 -4602
rect 29763 -4620 29787 -4602
rect 29787 -4620 29797 -4602
rect 29763 -4636 29797 -4620
rect 30135 -4550 30169 -4534
rect 30135 -4568 30161 -4550
rect 30161 -4568 30169 -4550
rect 30351 -4548 30385 -4539
rect 30351 -4573 30367 -4548
rect 30367 -4573 30385 -4548
rect 30411 -4636 30445 -4602
rect 31006 -4549 31044 -4515
rect 31168 -4559 31180 -4534
rect 31180 -4559 31202 -4534
rect 31168 -4568 31202 -4559
rect 31249 -4414 31283 -4398
rect 31249 -4432 31283 -4414
rect 31353 -4648 31391 -4614
rect 31627 -4432 31661 -4398
rect 31535 -4568 31569 -4534
rect 32251 -4424 32285 -4398
rect 32251 -4432 32282 -4424
rect 32282 -4432 32285 -4424
rect 31807 -4636 31841 -4602
rect 31879 -4620 31903 -4602
rect 31903 -4620 31913 -4602
rect 31879 -4636 31913 -4620
rect 32251 -4550 32285 -4534
rect 32251 -4568 32277 -4550
rect 32277 -4568 32285 -4550
rect 32467 -4548 32501 -4539
rect 32467 -4573 32483 -4548
rect 32483 -4573 32501 -4548
rect 32527 -4636 32561 -4602
rect 33122 -4549 33160 -4515
rect -9129 -4796 -9095 -4772
rect -9129 -4806 -9095 -4796
rect -9037 -4796 -9003 -4772
rect -9037 -4806 -9003 -4796
rect -8945 -4796 -8911 -4772
rect -8945 -4806 -8911 -4796
rect -8853 -4796 -8819 -4772
rect -8853 -4806 -8819 -4796
rect -8761 -4796 -8727 -4772
rect -8761 -4806 -8727 -4796
rect -8669 -4796 -8635 -4772
rect -8669 -4806 -8635 -4796
rect -8577 -4796 -8543 -4772
rect -8577 -4806 -8543 -4796
rect -8485 -4796 -8451 -4772
rect -8485 -4806 -8451 -4796
rect -8393 -4796 -8359 -4772
rect -8393 -4806 -8359 -4796
rect -8301 -4796 -8267 -4772
rect -8301 -4806 -8267 -4796
rect -8209 -4796 -8175 -4772
rect -8209 -4806 -8175 -4796
rect -8117 -4796 -8083 -4772
rect -8117 -4806 -8083 -4796
rect -8025 -4796 -7991 -4772
rect -8025 -4806 -7991 -4796
rect -7933 -4796 -7899 -4772
rect -7933 -4806 -7899 -4796
rect -7841 -4796 -7807 -4772
rect -7841 -4806 -7807 -4796
rect -7749 -4796 -7715 -4772
rect -7749 -4806 -7715 -4796
rect -7657 -4796 -7623 -4772
rect -7657 -4806 -7623 -4796
rect -7565 -4796 -7531 -4772
rect -7565 -4806 -7531 -4796
rect -7473 -4796 -7439 -4772
rect -7473 -4806 -7439 -4796
rect -7381 -4796 -7347 -4772
rect -7381 -4806 -7347 -4796
rect -7289 -4796 -7255 -4772
rect -7289 -4806 -7255 -4796
rect -7197 -4796 -7163 -4772
rect -7197 -4806 -7163 -4796
rect -7105 -4796 -7071 -4772
rect -7105 -4806 -7071 -4796
rect -7013 -4796 -6979 -4772
rect -7013 -4806 -6979 -4796
rect -6921 -4796 -6887 -4772
rect -6921 -4806 -6887 -4796
rect -6829 -4796 -6795 -4772
rect -6829 -4806 -6795 -4796
rect -6737 -4796 -6703 -4772
rect -6737 -4806 -6703 -4796
rect -6645 -4796 -6611 -4772
rect -6645 -4806 -6611 -4796
rect -6553 -4796 -6519 -4772
rect -6553 -4806 -6519 -4796
rect -6461 -4796 -6427 -4772
rect -6461 -4806 -6427 -4796
rect -6369 -4796 -6335 -4772
rect -6369 -4806 -6335 -4796
rect -6277 -4796 -6243 -4772
rect -6277 -4806 -6243 -4796
rect -6185 -4796 -6151 -4772
rect -6185 -4806 -6151 -4796
rect -6093 -4796 -6059 -4772
rect -6093 -4806 -6059 -4796
rect -6001 -4796 -5967 -4772
rect -6001 -4806 -5967 -4796
rect -5909 -4796 -5875 -4772
rect -5909 -4806 -5875 -4796
rect -5817 -4796 -5783 -4772
rect -5817 -4806 -5783 -4796
rect -5725 -4796 -5691 -4772
rect -5725 -4806 -5691 -4796
rect -5633 -4796 -5599 -4772
rect -5633 -4806 -5599 -4796
rect -5541 -4796 -5507 -4772
rect -5541 -4806 -5507 -4796
rect -5449 -4796 -5415 -4772
rect -5449 -4806 -5415 -4796
rect -5357 -4796 -5323 -4772
rect -5357 -4806 -5323 -4796
rect -5265 -4796 -5231 -4772
rect -5265 -4806 -5231 -4796
rect -5173 -4796 -5139 -4772
rect -5173 -4806 -5139 -4796
rect -5081 -4796 -5047 -4772
rect -5081 -4806 -5047 -4796
rect -4989 -4796 -4955 -4772
rect -4989 -4806 -4955 -4796
rect -4897 -4796 -4863 -4772
rect -4897 -4806 -4863 -4796
rect -4805 -4796 -4771 -4772
rect -4805 -4806 -4771 -4796
rect -4713 -4796 -4679 -4772
rect -4713 -4806 -4679 -4796
rect -4621 -4796 -4587 -4772
rect -4621 -4806 -4587 -4796
rect -4529 -4796 -4495 -4772
rect -4529 -4806 -4495 -4796
rect -4437 -4796 -4403 -4772
rect -4437 -4806 -4403 -4796
rect -4345 -4796 -4311 -4772
rect -4345 -4806 -4311 -4796
rect -4253 -4796 -4219 -4772
rect -4253 -4806 -4219 -4796
rect -4161 -4796 -4127 -4772
rect -4161 -4806 -4127 -4796
rect -4069 -4796 -4035 -4772
rect -4069 -4806 -4035 -4796
rect -3977 -4796 -3943 -4772
rect -3977 -4806 -3943 -4796
rect -3885 -4796 -3851 -4772
rect -3885 -4806 -3851 -4796
rect -3793 -4796 -3759 -4772
rect -3793 -4806 -3759 -4796
rect -3701 -4796 -3667 -4772
rect -3701 -4806 -3667 -4796
rect -3609 -4796 -3575 -4772
rect -3609 -4806 -3575 -4796
rect -3517 -4796 -3483 -4772
rect -3517 -4806 -3483 -4796
rect -3425 -4796 -3391 -4772
rect -3425 -4806 -3391 -4796
rect -3333 -4796 -3299 -4772
rect -3333 -4806 -3299 -4796
rect -3241 -4796 -3207 -4772
rect -3241 -4806 -3207 -4796
rect -3149 -4796 -3115 -4772
rect -3149 -4806 -3115 -4796
rect -3057 -4796 -3023 -4772
rect -3057 -4806 -3023 -4796
rect -2965 -4796 -2931 -4772
rect -2965 -4806 -2931 -4796
rect -2873 -4796 -2839 -4772
rect -2873 -4806 -2839 -4796
rect -2781 -4796 -2747 -4772
rect -2781 -4806 -2747 -4796
rect -2689 -4796 -2655 -4772
rect -2689 -4806 -2655 -4796
rect -2597 -4796 -2563 -4772
rect -2597 -4806 -2563 -4796
rect -2505 -4796 -2471 -4772
rect -2505 -4806 -2471 -4796
rect -2413 -4796 -2379 -4772
rect -2413 -4806 -2379 -4796
rect -2321 -4796 -2287 -4772
rect -2321 -4806 -2287 -4796
rect -2229 -4796 -2195 -4772
rect -2229 -4806 -2195 -4796
rect -2137 -4796 -2103 -4772
rect -2137 -4806 -2103 -4796
rect -2045 -4796 -2011 -4772
rect -2045 -4806 -2011 -4796
rect -1953 -4796 -1919 -4772
rect -1953 -4806 -1919 -4796
rect -1861 -4796 -1827 -4772
rect -1861 -4806 -1827 -4796
rect -1769 -4796 -1735 -4772
rect -1769 -4806 -1735 -4796
rect -1677 -4796 -1643 -4772
rect -1677 -4806 -1643 -4796
rect -1585 -4796 -1551 -4772
rect -1585 -4806 -1551 -4796
rect -1493 -4796 -1459 -4772
rect -1493 -4806 -1459 -4796
rect -1401 -4796 -1367 -4772
rect -1401 -4806 -1367 -4796
rect -1309 -4796 -1275 -4772
rect -1309 -4806 -1275 -4796
rect -1217 -4796 -1183 -4772
rect -1217 -4806 -1183 -4796
rect -1125 -4796 -1091 -4772
rect -1125 -4806 -1091 -4796
rect -1033 -4796 -999 -4772
rect -1033 -4806 -999 -4796
rect -941 -4796 -907 -4772
rect -941 -4806 -907 -4796
rect -849 -4796 -815 -4772
rect -849 -4806 -815 -4796
rect -757 -4796 -723 -4772
rect -757 -4806 -723 -4796
rect -665 -4796 -631 -4772
rect -665 -4806 -631 -4796
rect -573 -4796 -539 -4772
rect -573 -4806 -539 -4796
rect -481 -4796 -447 -4772
rect -481 -4806 -447 -4796
rect -389 -4796 -355 -4772
rect -389 -4806 -355 -4796
rect -297 -4796 -263 -4772
rect -297 -4806 -263 -4796
rect -205 -4796 -171 -4772
rect -205 -4806 -171 -4796
rect -113 -4796 -79 -4772
rect -113 -4806 -79 -4796
rect -21 -4796 13 -4772
rect -21 -4806 13 -4796
rect 71 -4796 105 -4772
rect 71 -4806 105 -4796
rect 163 -4796 197 -4772
rect 163 -4806 197 -4796
rect 255 -4796 289 -4772
rect 255 -4806 289 -4796
rect 347 -4796 381 -4772
rect 347 -4806 381 -4796
rect 439 -4796 473 -4772
rect 439 -4806 473 -4796
rect 531 -4796 565 -4772
rect 531 -4806 565 -4796
rect 623 -4796 657 -4772
rect 623 -4806 657 -4796
rect 715 -4796 749 -4772
rect 715 -4806 749 -4796
rect 807 -4796 841 -4772
rect 807 -4806 841 -4796
rect 899 -4796 933 -4772
rect 899 -4806 933 -4796
rect 991 -4796 1025 -4772
rect 991 -4806 1025 -4796
rect 1083 -4796 1117 -4772
rect 1083 -4806 1117 -4796
rect 1175 -4796 1209 -4772
rect 1175 -4806 1209 -4796
rect 1267 -4796 1301 -4772
rect 1267 -4806 1301 -4796
rect 1359 -4796 1393 -4772
rect 1359 -4806 1393 -4796
rect 1451 -4796 1485 -4772
rect 1451 -4806 1485 -4796
rect 1543 -4796 1577 -4772
rect 1543 -4806 1577 -4796
rect 1635 -4796 1669 -4772
rect 1635 -4806 1669 -4796
rect 1727 -4796 1761 -4772
rect 1727 -4806 1761 -4796
rect 1819 -4796 1853 -4772
rect 1819 -4806 1853 -4796
rect 1911 -4796 1945 -4772
rect 1911 -4806 1945 -4796
rect 2003 -4796 2037 -4772
rect 2003 -4806 2037 -4796
rect 2095 -4796 2129 -4772
rect 2095 -4806 2129 -4796
rect 2187 -4796 2221 -4772
rect 2187 -4806 2221 -4796
rect 2279 -4796 2313 -4772
rect 2279 -4806 2313 -4796
rect 2371 -4796 2405 -4772
rect 2371 -4806 2405 -4796
rect 2463 -4796 2497 -4772
rect 2463 -4806 2497 -4796
rect 2555 -4796 2589 -4772
rect 2555 -4806 2589 -4796
rect 2647 -4796 2681 -4772
rect 2647 -4806 2681 -4796
rect 2739 -4796 2773 -4772
rect 2739 -4806 2773 -4796
rect 2831 -4796 2865 -4772
rect 2831 -4806 2865 -4796
rect 2923 -4796 2957 -4772
rect 2923 -4806 2957 -4796
rect 3015 -4796 3049 -4772
rect 3015 -4806 3049 -4796
rect 3107 -4796 3141 -4772
rect 3107 -4806 3141 -4796
rect 3199 -4796 3233 -4772
rect 3199 -4806 3233 -4796
rect 3291 -4796 3325 -4772
rect 3291 -4806 3325 -4796
rect 3383 -4796 3417 -4772
rect 3383 -4806 3417 -4796
rect 3475 -4796 3509 -4772
rect 3475 -4806 3509 -4796
rect 3567 -4796 3601 -4772
rect 3567 -4806 3601 -4796
rect 3659 -4796 3693 -4772
rect 3659 -4806 3693 -4796
rect 3751 -4796 3785 -4772
rect 3751 -4806 3785 -4796
rect 3843 -4796 3877 -4772
rect 3843 -4806 3877 -4796
rect 3935 -4796 3969 -4772
rect 3935 -4806 3969 -4796
rect 4027 -4796 4061 -4772
rect 4027 -4806 4061 -4796
rect 4119 -4796 4153 -4772
rect 4119 -4806 4153 -4796
rect 4211 -4796 4245 -4772
rect 4211 -4806 4245 -4796
rect 4303 -4796 4337 -4772
rect 4303 -4806 4337 -4796
rect 4395 -4796 4429 -4772
rect 4395 -4806 4429 -4796
rect 4487 -4796 4521 -4772
rect 4487 -4806 4521 -4796
rect 4579 -4796 4613 -4772
rect 4579 -4806 4613 -4796
rect 4671 -4796 4705 -4772
rect 4671 -4806 4705 -4796
rect 4763 -4796 4797 -4772
rect 4763 -4806 4797 -4796
rect 4855 -4796 4889 -4772
rect 4855 -4806 4889 -4796
rect 4947 -4796 4981 -4772
rect 4947 -4806 4981 -4796
rect 5039 -4796 5073 -4772
rect 5039 -4806 5073 -4796
rect 5131 -4796 5165 -4772
rect 5131 -4806 5165 -4796
rect 5223 -4796 5257 -4772
rect 5223 -4806 5257 -4796
rect 5315 -4796 5349 -4772
rect 5315 -4806 5349 -4796
rect 5407 -4796 5441 -4772
rect 5407 -4806 5441 -4796
rect 5499 -4796 5533 -4772
rect 5499 -4806 5533 -4796
rect 5591 -4796 5625 -4772
rect 5591 -4806 5625 -4796
rect 5683 -4796 5717 -4772
rect 5683 -4806 5717 -4796
rect 5775 -4796 5809 -4772
rect 5775 -4806 5809 -4796
rect 5867 -4796 5901 -4772
rect 5867 -4806 5901 -4796
rect 5959 -4796 5993 -4772
rect 5959 -4806 5993 -4796
rect 6051 -4796 6085 -4772
rect 6051 -4806 6085 -4796
rect 6143 -4796 6177 -4772
rect 6143 -4806 6177 -4796
rect 6235 -4796 6269 -4772
rect 6235 -4806 6269 -4796
rect 6327 -4796 6361 -4772
rect 6327 -4806 6361 -4796
rect 6419 -4796 6453 -4772
rect 6419 -4806 6453 -4796
rect 6511 -4796 6545 -4772
rect 6511 -4806 6545 -4796
rect 6603 -4796 6637 -4772
rect 6603 -4806 6637 -4796
rect 6695 -4796 6729 -4772
rect 6695 -4806 6729 -4796
rect 6787 -4796 6821 -4772
rect 6787 -4806 6821 -4796
rect 6879 -4796 6913 -4772
rect 6879 -4806 6913 -4796
rect 6971 -4796 7005 -4772
rect 6971 -4806 7005 -4796
rect 7063 -4796 7097 -4772
rect 7063 -4806 7097 -4796
rect 7155 -4796 7189 -4772
rect 7155 -4806 7189 -4796
rect 7247 -4796 7281 -4772
rect 7247 -4806 7281 -4796
rect 7339 -4796 7373 -4772
rect 7339 -4806 7373 -4796
rect 7431 -4796 7465 -4772
rect 7431 -4806 7465 -4796
rect 7523 -4796 7557 -4772
rect 7523 -4806 7557 -4796
rect 7615 -4796 7649 -4772
rect 7615 -4806 7649 -4796
rect 7707 -4796 7741 -4772
rect 7707 -4806 7741 -4796
rect 7799 -4796 7833 -4772
rect 7799 -4806 7833 -4796
rect 7891 -4796 7925 -4772
rect 7891 -4806 7925 -4796
rect 7983 -4796 8017 -4772
rect 7983 -4806 8017 -4796
rect 8075 -4796 8109 -4772
rect 8075 -4806 8109 -4796
rect 8167 -4796 8201 -4772
rect 8167 -4806 8201 -4796
rect 8259 -4796 8293 -4772
rect 8259 -4806 8293 -4796
rect 8351 -4796 8385 -4772
rect 8351 -4806 8385 -4796
rect 8443 -4796 8477 -4772
rect 8443 -4806 8477 -4796
rect 8535 -4796 8569 -4772
rect 8535 -4806 8569 -4796
rect 8627 -4796 8661 -4772
rect 8627 -4806 8661 -4796
rect 8719 -4796 8753 -4772
rect 8719 -4806 8753 -4796
rect 8811 -4796 8845 -4772
rect 8811 -4806 8845 -4796
rect 8903 -4796 8937 -4772
rect 8903 -4806 8937 -4796
rect 8995 -4796 9029 -4772
rect 8995 -4806 9029 -4796
rect 9087 -4796 9121 -4772
rect 9087 -4806 9121 -4796
rect 9179 -4796 9213 -4772
rect 9179 -4806 9213 -4796
rect 9271 -4796 9305 -4772
rect 9271 -4806 9305 -4796
rect 9363 -4796 9397 -4772
rect 9363 -4806 9397 -4796
rect 9455 -4796 9489 -4772
rect 9455 -4806 9489 -4796
rect 9547 -4796 9581 -4772
rect 9547 -4806 9581 -4796
rect 9639 -4796 9673 -4772
rect 9639 -4806 9673 -4796
rect 9731 -4796 9765 -4772
rect 9731 -4806 9765 -4796
rect 9823 -4796 9857 -4772
rect 9823 -4806 9857 -4796
rect 9915 -4796 9949 -4772
rect 9915 -4806 9949 -4796
rect 10007 -4796 10041 -4772
rect 10007 -4806 10041 -4796
rect 10099 -4796 10133 -4772
rect 10099 -4806 10133 -4796
rect 10191 -4796 10225 -4772
rect 10191 -4806 10225 -4796
rect 10283 -4796 10317 -4772
rect 10283 -4806 10317 -4796
rect 10375 -4796 10409 -4772
rect 10375 -4806 10409 -4796
rect 10467 -4796 10501 -4772
rect 10467 -4806 10501 -4796
rect 10559 -4796 10593 -4772
rect 10559 -4806 10593 -4796
rect 10651 -4796 10685 -4772
rect 10651 -4806 10685 -4796
rect 10743 -4796 10777 -4772
rect 10743 -4806 10777 -4796
rect 10835 -4796 10869 -4772
rect 10835 -4806 10869 -4796
rect 10927 -4796 10961 -4772
rect 10927 -4806 10961 -4796
rect 11019 -4796 11053 -4772
rect 11019 -4806 11053 -4796
rect 11111 -4796 11145 -4772
rect 11111 -4806 11145 -4796
rect 11203 -4796 11237 -4772
rect 11203 -4806 11237 -4796
rect 11295 -4796 11329 -4772
rect 11295 -4806 11329 -4796
rect 11387 -4796 11421 -4772
rect 11387 -4806 11421 -4796
rect 11479 -4796 11513 -4772
rect 11479 -4806 11513 -4796
rect 11571 -4796 11605 -4772
rect 11571 -4806 11605 -4796
rect 11663 -4796 11697 -4772
rect 11663 -4806 11697 -4796
rect 11755 -4796 11789 -4772
rect 11755 -4806 11789 -4796
rect 11847 -4796 11881 -4772
rect 11847 -4806 11881 -4796
rect 11939 -4796 11973 -4772
rect 11939 -4806 11973 -4796
rect 12031 -4796 12065 -4772
rect 12031 -4806 12065 -4796
rect 12123 -4796 12157 -4772
rect 12123 -4806 12157 -4796
rect 12215 -4796 12249 -4772
rect 12215 -4806 12249 -4796
rect 12307 -4796 12341 -4772
rect 12307 -4806 12341 -4796
rect 12399 -4796 12433 -4772
rect 12399 -4806 12433 -4796
rect 12491 -4796 12525 -4772
rect 12491 -4806 12525 -4796
rect 12583 -4796 12617 -4772
rect 12583 -4806 12617 -4796
rect 12675 -4796 12709 -4772
rect 12675 -4806 12709 -4796
rect 12767 -4796 12801 -4772
rect 12767 -4806 12801 -4796
rect 12859 -4796 12893 -4772
rect 12859 -4806 12893 -4796
rect 12951 -4796 12985 -4772
rect 12951 -4806 12985 -4796
rect 13043 -4796 13077 -4772
rect 13043 -4806 13077 -4796
rect 13135 -4796 13169 -4772
rect 13135 -4806 13169 -4796
rect 13227 -4796 13261 -4772
rect 13227 -4806 13261 -4796
rect 13319 -4796 13353 -4772
rect 13319 -4806 13353 -4796
rect 13411 -4796 13445 -4772
rect 13411 -4806 13445 -4796
rect 13503 -4796 13537 -4772
rect 13503 -4806 13537 -4796
rect 13595 -4796 13629 -4772
rect 13595 -4806 13629 -4796
rect 13687 -4796 13721 -4772
rect 13687 -4806 13721 -4796
rect 13779 -4796 13813 -4772
rect 13779 -4806 13813 -4796
rect 13871 -4796 13905 -4772
rect 13871 -4806 13905 -4796
rect 13963 -4796 13997 -4772
rect 13963 -4806 13997 -4796
rect 14055 -4796 14089 -4772
rect 14055 -4806 14089 -4796
rect 14147 -4796 14181 -4772
rect 14147 -4806 14181 -4796
rect 14239 -4796 14273 -4772
rect 14239 -4806 14273 -4796
rect 14331 -4796 14365 -4772
rect 14331 -4806 14365 -4796
rect 14423 -4796 14457 -4772
rect 14423 -4806 14457 -4796
rect 14515 -4796 14549 -4772
rect 14515 -4806 14549 -4796
rect 14607 -4796 14641 -4772
rect 14607 -4806 14641 -4796
rect 14699 -4796 14733 -4772
rect 14699 -4806 14733 -4796
rect 14791 -4796 14825 -4772
rect 14791 -4806 14825 -4796
rect 14883 -4796 14917 -4772
rect 14883 -4806 14917 -4796
rect 14975 -4796 15009 -4772
rect 14975 -4806 15009 -4796
rect 15067 -4796 15101 -4772
rect 15067 -4806 15101 -4796
rect 15159 -4796 15193 -4772
rect 15159 -4806 15193 -4796
rect 15251 -4796 15285 -4772
rect 15251 -4806 15285 -4796
rect 15343 -4796 15377 -4772
rect 15343 -4806 15377 -4796
rect 15435 -4796 15469 -4772
rect 15435 -4806 15469 -4796
rect 15527 -4796 15561 -4772
rect 15527 -4806 15561 -4796
rect 15619 -4796 15653 -4772
rect 15619 -4806 15653 -4796
rect 15711 -4796 15745 -4772
rect 15711 -4806 15745 -4796
rect 15803 -4796 15837 -4772
rect 15803 -4806 15837 -4796
rect 15895 -4796 15929 -4772
rect 15895 -4806 15929 -4796
rect 15987 -4796 16021 -4772
rect 15987 -4806 16021 -4796
rect 16079 -4796 16113 -4772
rect 16079 -4806 16113 -4796
rect 16171 -4796 16205 -4772
rect 16171 -4806 16205 -4796
rect 16263 -4796 16297 -4772
rect 16263 -4806 16297 -4796
rect 16355 -4796 16389 -4772
rect 16355 -4806 16389 -4796
rect 16447 -4796 16481 -4772
rect 16447 -4806 16481 -4796
rect 16539 -4796 16573 -4772
rect 16539 -4806 16573 -4796
rect 16631 -4796 16665 -4772
rect 16631 -4806 16665 -4796
rect 16723 -4796 16757 -4772
rect 16723 -4806 16757 -4796
rect 16815 -4796 16849 -4772
rect 16815 -4806 16849 -4796
rect 16907 -4796 16941 -4772
rect 16907 -4806 16941 -4796
rect 16999 -4796 17033 -4772
rect 16999 -4806 17033 -4796
rect 17091 -4796 17125 -4772
rect 17091 -4806 17125 -4796
rect 17183 -4796 17217 -4772
rect 17183 -4806 17217 -4796
rect 17275 -4796 17309 -4772
rect 17275 -4806 17309 -4796
rect 17367 -4796 17401 -4772
rect 17367 -4806 17401 -4796
rect 17459 -4796 17493 -4772
rect 17459 -4806 17493 -4796
rect 17551 -4796 17585 -4772
rect 17551 -4806 17585 -4796
rect 17643 -4796 17677 -4772
rect 17643 -4806 17677 -4796
rect 17735 -4796 17769 -4772
rect 17735 -4806 17769 -4796
rect 17827 -4796 17861 -4772
rect 17827 -4806 17861 -4796
rect 17919 -4796 17953 -4772
rect 17919 -4806 17953 -4796
rect 18011 -4796 18045 -4772
rect 18011 -4806 18045 -4796
rect 18103 -4796 18137 -4772
rect 18103 -4806 18137 -4796
rect 18195 -4796 18229 -4772
rect 18195 -4806 18229 -4796
rect 18287 -4796 18321 -4772
rect 18287 -4806 18321 -4796
rect 18379 -4796 18413 -4772
rect 18379 -4806 18413 -4796
rect 18471 -4796 18505 -4772
rect 18471 -4806 18505 -4796
rect 18563 -4796 18597 -4772
rect 18563 -4806 18597 -4796
rect 18655 -4796 18689 -4772
rect 18655 -4806 18689 -4796
rect 18747 -4796 18781 -4772
rect 18747 -4806 18781 -4796
rect 18839 -4796 18873 -4772
rect 18839 -4806 18873 -4796
rect 18931 -4796 18965 -4772
rect 18931 -4806 18965 -4796
rect 19023 -4796 19057 -4772
rect 19023 -4806 19057 -4796
rect 19115 -4796 19149 -4772
rect 19115 -4806 19149 -4796
rect 19207 -4796 19241 -4772
rect 19207 -4806 19241 -4796
rect 19299 -4796 19333 -4772
rect 19299 -4806 19333 -4796
rect 19391 -4796 19425 -4772
rect 19391 -4806 19425 -4796
rect 19483 -4796 19517 -4772
rect 19483 -4806 19517 -4796
rect 19575 -4796 19609 -4772
rect 19575 -4806 19609 -4796
rect 19667 -4796 19701 -4772
rect 19667 -4806 19701 -4796
rect 19759 -4796 19793 -4772
rect 19759 -4806 19793 -4796
rect 19851 -4796 19885 -4772
rect 19851 -4806 19885 -4796
rect 19943 -4796 19977 -4772
rect 19943 -4806 19977 -4796
rect 20035 -4796 20069 -4772
rect 20035 -4806 20069 -4796
rect 20127 -4796 20161 -4772
rect 20127 -4806 20161 -4796
rect 20219 -4796 20253 -4772
rect 20219 -4806 20253 -4796
rect 20311 -4796 20345 -4772
rect 20311 -4806 20345 -4796
rect 20403 -4796 20437 -4772
rect 20403 -4806 20437 -4796
rect 20495 -4796 20529 -4772
rect 20495 -4806 20529 -4796
rect 20587 -4796 20621 -4772
rect 20587 -4806 20621 -4796
rect 20679 -4796 20713 -4772
rect 20679 -4806 20713 -4796
rect 20771 -4796 20805 -4772
rect 20771 -4806 20805 -4796
rect 20863 -4796 20897 -4772
rect 20863 -4806 20897 -4796
rect 20955 -4796 20989 -4772
rect 20955 -4806 20989 -4796
rect 21047 -4796 21081 -4772
rect 21047 -4806 21081 -4796
rect 21139 -4796 21173 -4772
rect 21139 -4806 21173 -4796
rect 21231 -4796 21265 -4772
rect 21231 -4806 21265 -4796
rect 21323 -4796 21357 -4772
rect 21323 -4806 21357 -4796
rect 21415 -4796 21449 -4772
rect 21415 -4806 21449 -4796
rect 21507 -4796 21541 -4772
rect 21507 -4806 21541 -4796
rect 21599 -4796 21633 -4772
rect 21599 -4806 21633 -4796
rect 21691 -4796 21725 -4772
rect 21691 -4806 21725 -4796
rect 21783 -4796 21817 -4772
rect 21783 -4806 21817 -4796
rect 21875 -4796 21909 -4772
rect 21875 -4806 21909 -4796
rect 21967 -4796 22001 -4772
rect 21967 -4806 22001 -4796
rect 22059 -4796 22093 -4772
rect 22059 -4806 22093 -4796
rect 22151 -4796 22185 -4772
rect 22151 -4806 22185 -4796
rect 22243 -4796 22277 -4772
rect 22243 -4806 22277 -4796
rect 22335 -4796 22369 -4772
rect 22335 -4806 22369 -4796
rect 22427 -4796 22461 -4772
rect 22427 -4806 22461 -4796
rect 22519 -4796 22553 -4772
rect 22519 -4806 22553 -4796
rect 22611 -4796 22645 -4772
rect 22611 -4806 22645 -4796
rect 22703 -4796 22737 -4772
rect 22703 -4806 22737 -4796
rect 22795 -4796 22829 -4772
rect 22795 -4806 22829 -4796
rect 22887 -4796 22921 -4772
rect 22887 -4806 22921 -4796
rect 22979 -4796 23013 -4772
rect 22979 -4806 23013 -4796
rect 23071 -4796 23105 -4772
rect 23071 -4806 23105 -4796
rect 23163 -4796 23197 -4772
rect 23163 -4806 23197 -4796
rect 23255 -4796 23289 -4772
rect 23255 -4806 23289 -4796
rect 23347 -4796 23381 -4772
rect 23347 -4806 23381 -4796
rect 23439 -4796 23473 -4772
rect 23439 -4806 23473 -4796
rect 23531 -4796 23565 -4772
rect 23531 -4806 23565 -4796
rect 23623 -4796 23657 -4772
rect 23623 -4806 23657 -4796
rect 23715 -4796 23749 -4772
rect 23715 -4806 23749 -4796
rect 23807 -4796 23841 -4772
rect 23807 -4806 23841 -4796
rect 23899 -4796 23933 -4772
rect 23899 -4806 23933 -4796
rect 23991 -4796 24025 -4772
rect 23991 -4806 24025 -4796
rect 24083 -4796 24117 -4772
rect 24083 -4806 24117 -4796
rect 24175 -4796 24209 -4772
rect 24175 -4806 24209 -4796
rect 24267 -4796 24301 -4772
rect 24267 -4806 24301 -4796
rect 24359 -4796 24393 -4772
rect 24359 -4806 24393 -4796
rect 24451 -4796 24485 -4772
rect 24451 -4806 24485 -4796
rect 24543 -4796 24577 -4772
rect 24543 -4806 24577 -4796
rect 24635 -4796 24669 -4772
rect 24635 -4806 24669 -4796
rect 24727 -4796 24761 -4772
rect 24727 -4806 24761 -4796
rect 24819 -4796 24853 -4772
rect 24819 -4806 24853 -4796
rect 24911 -4796 24945 -4772
rect 24911 -4806 24945 -4796
rect 25003 -4796 25037 -4772
rect 25003 -4806 25037 -4796
rect 25095 -4796 25129 -4772
rect 25095 -4806 25129 -4796
rect 25187 -4796 25221 -4772
rect 25187 -4806 25221 -4796
rect 25279 -4796 25313 -4772
rect 25279 -4806 25313 -4796
rect 25371 -4796 25405 -4772
rect 25371 -4806 25405 -4796
rect 25463 -4796 25497 -4772
rect 25463 -4806 25497 -4796
rect 25555 -4796 25589 -4772
rect 25555 -4806 25589 -4796
rect 25647 -4796 25681 -4772
rect 25647 -4806 25681 -4796
rect 25739 -4796 25773 -4772
rect 25739 -4806 25773 -4796
rect 25831 -4796 25865 -4772
rect 25831 -4806 25865 -4796
rect 25923 -4796 25957 -4772
rect 25923 -4806 25957 -4796
rect 26015 -4796 26049 -4772
rect 26015 -4806 26049 -4796
rect 26107 -4796 26141 -4772
rect 26107 -4806 26141 -4796
rect 26199 -4796 26233 -4772
rect 26199 -4806 26233 -4796
rect 26291 -4796 26325 -4772
rect 26291 -4806 26325 -4796
rect 26383 -4796 26417 -4772
rect 26383 -4806 26417 -4796
rect 26475 -4796 26509 -4772
rect 26475 -4806 26509 -4796
rect 26567 -4796 26601 -4772
rect 26567 -4806 26601 -4796
rect 26659 -4796 26693 -4772
rect 26659 -4806 26693 -4796
rect 26751 -4796 26785 -4772
rect 26751 -4806 26785 -4796
rect 26843 -4796 26877 -4772
rect 26843 -4806 26877 -4796
rect 26935 -4796 26969 -4772
rect 26935 -4806 26969 -4796
rect 27027 -4796 27061 -4772
rect 27027 -4806 27061 -4796
rect 27119 -4796 27153 -4772
rect 27119 -4806 27153 -4796
rect 27211 -4796 27245 -4772
rect 27211 -4806 27245 -4796
rect 27303 -4796 27337 -4772
rect 27303 -4806 27337 -4796
rect 27395 -4796 27429 -4772
rect 27395 -4806 27429 -4796
rect 27487 -4796 27521 -4772
rect 27487 -4806 27521 -4796
rect 27579 -4796 27613 -4772
rect 27579 -4806 27613 -4796
rect 27671 -4796 27705 -4772
rect 27671 -4806 27705 -4796
rect 27763 -4796 27797 -4772
rect 27763 -4806 27797 -4796
rect 27855 -4796 27889 -4772
rect 27855 -4806 27889 -4796
rect 27947 -4796 27981 -4772
rect 27947 -4806 27981 -4796
rect 28039 -4796 28073 -4772
rect 28039 -4806 28073 -4796
rect 28131 -4796 28165 -4772
rect 28131 -4806 28165 -4796
rect 28223 -4796 28257 -4772
rect 28223 -4806 28257 -4796
rect 28315 -4796 28349 -4772
rect 28315 -4806 28349 -4796
rect 28407 -4796 28441 -4772
rect 28407 -4806 28441 -4796
rect 28499 -4796 28533 -4772
rect 28499 -4806 28533 -4796
rect 28591 -4796 28625 -4772
rect 28591 -4806 28625 -4796
rect 28683 -4796 28717 -4772
rect 28683 -4806 28717 -4796
rect 28775 -4796 28809 -4772
rect 28775 -4806 28809 -4796
rect 28867 -4796 28901 -4772
rect 28867 -4806 28901 -4796
rect 28959 -4796 28993 -4772
rect 28959 -4806 28993 -4796
rect 29051 -4796 29085 -4772
rect 29051 -4806 29085 -4796
rect 29143 -4796 29177 -4772
rect 29143 -4806 29177 -4796
rect 29235 -4796 29269 -4772
rect 29235 -4806 29269 -4796
rect 29327 -4796 29361 -4772
rect 29327 -4806 29361 -4796
rect 29419 -4796 29453 -4772
rect 29419 -4806 29453 -4796
rect 29511 -4796 29545 -4772
rect 29511 -4806 29545 -4796
rect 29603 -4796 29637 -4772
rect 29603 -4806 29637 -4796
rect 29695 -4796 29729 -4772
rect 29695 -4806 29729 -4796
rect 29787 -4796 29821 -4772
rect 29787 -4806 29821 -4796
rect 29879 -4796 29913 -4772
rect 29879 -4806 29913 -4796
rect 29971 -4796 30005 -4772
rect 29971 -4806 30005 -4796
rect 30063 -4796 30097 -4772
rect 30063 -4806 30097 -4796
rect 30155 -4796 30189 -4772
rect 30155 -4806 30189 -4796
rect 30247 -4796 30281 -4772
rect 30247 -4806 30281 -4796
rect 30339 -4796 30373 -4772
rect 30339 -4806 30373 -4796
rect 30431 -4796 30465 -4772
rect 30431 -4806 30465 -4796
rect 30523 -4796 30557 -4772
rect 30523 -4806 30557 -4796
rect 30615 -4796 30649 -4772
rect 30615 -4806 30649 -4796
rect 30707 -4796 30741 -4772
rect 30707 -4806 30741 -4796
rect 30799 -4796 30833 -4772
rect 30799 -4806 30833 -4796
rect 30891 -4796 30925 -4772
rect 30891 -4806 30925 -4796
rect 30983 -4796 31017 -4772
rect 30983 -4806 31017 -4796
rect 31075 -4796 31109 -4772
rect 31075 -4806 31109 -4796
rect 31167 -4796 31201 -4772
rect 31167 -4806 31201 -4796
rect 31259 -4796 31293 -4772
rect 31259 -4806 31293 -4796
rect 31351 -4796 31385 -4772
rect 31351 -4806 31385 -4796
rect 31443 -4796 31477 -4772
rect 31443 -4806 31477 -4796
rect 31535 -4796 31569 -4772
rect 31535 -4806 31569 -4796
rect 31627 -4796 31661 -4772
rect 31627 -4806 31661 -4796
rect 31719 -4796 31753 -4772
rect 31719 -4806 31753 -4796
rect 31811 -4796 31845 -4772
rect 31811 -4806 31845 -4796
rect 31903 -4796 31937 -4772
rect 31903 -4806 31937 -4796
rect 31995 -4796 32029 -4772
rect 31995 -4806 32029 -4796
rect 32087 -4796 32121 -4772
rect 32087 -4806 32121 -4796
rect 32179 -4796 32213 -4772
rect 32179 -4806 32213 -4796
rect 32271 -4796 32305 -4772
rect 32271 -4806 32305 -4796
rect 32363 -4796 32397 -4772
rect 32363 -4806 32397 -4796
rect 32455 -4796 32489 -4772
rect 32455 -4806 32489 -4796
rect 32547 -4796 32581 -4772
rect 32547 -4806 32581 -4796
rect 32639 -4796 32673 -4772
rect 32639 -4806 32673 -4796
rect 32731 -4796 32765 -4772
rect 32731 -4806 32765 -4796
rect 32823 -4796 32857 -4772
rect 32823 -4806 32857 -4796
rect 32915 -4796 32949 -4772
rect 32915 -4806 32949 -4796
rect 33007 -4796 33041 -4772
rect 33007 -4806 33041 -4796
rect 33099 -4796 33133 -4772
rect 33099 -4806 33133 -4796
rect 4254 -7545 4290 -7518
rect 4254 -25711 4255 -7545
rect 4255 -25711 4289 -7545
rect 4289 -25711 4290 -7545
rect 4369 -9011 4403 -7635
rect 7798 -7545 7834 -7519
rect 4369 -10521 4403 -9145
rect 4369 -12031 4403 -10655
rect 4369 -13541 4403 -12165
rect 4369 -15051 4403 -13675
rect 4369 -16561 4403 -15185
rect 4369 -18071 4403 -16695
rect 4369 -19581 4403 -18205
rect 4369 -21091 4403 -19715
rect 4369 -22601 4403 -21225
rect 4369 -24111 4403 -22735
rect 4369 -25621 4403 -24245
rect 4254 -25771 4290 -25711
rect 6027 -9011 6061 -7635
rect 6027 -10521 6061 -9145
rect 6027 -12031 6061 -10655
rect 6027 -13541 6061 -12165
rect 6027 -15051 6061 -13675
rect 6027 -16561 6061 -15185
rect 6027 -18071 6061 -16695
rect 6027 -19581 6061 -18205
rect 6027 -21091 6061 -19715
rect 6027 -22601 6061 -21225
rect 6027 -24111 6061 -22735
rect 6027 -25621 6061 -24245
rect 7685 -9011 7719 -7635
rect 7685 -10521 7719 -9145
rect 7685 -12031 7719 -10655
rect 7685 -13541 7719 -12165
rect 7685 -15051 7719 -13675
rect 7685 -16561 7719 -15185
rect 7685 -18071 7719 -16695
rect 7685 -19581 7719 -18205
rect 7685 -21091 7719 -19715
rect 7685 -22601 7719 -21225
rect 7685 -24111 7719 -22735
rect 7685 -25621 7719 -24245
rect 7798 -25711 7799 -7545
rect 7799 -25711 7833 -7545
rect 7833 -25711 7834 -7545
rect 10176 -7628 10210 -7594
rect 10176 -7956 10210 -7922
rect 13064 -7629 13098 -7595
rect 13322 -7629 13356 -7595
rect 13064 -7957 13098 -7923
rect 13580 -7629 13614 -7595
rect 13838 -7629 13872 -7595
rect 14096 -7629 14130 -7595
rect 13322 -7957 13356 -7923
rect 13580 -7957 13614 -7923
rect 13838 -7957 13872 -7923
rect 14096 -7957 14130 -7923
rect 9036 -8675 9209 -8657
rect 9036 -8937 9055 -8675
rect 9055 -8937 9192 -8675
rect 9192 -8937 9209 -8675
rect 10093 -8568 10173 -8567
rect 10093 -8602 10173 -8568
rect 10093 -8628 10173 -8602
rect 10094 -8806 10174 -8788
rect 10094 -8840 10174 -8806
rect 10094 -8849 10174 -8840
rect 9036 -8959 9209 -8937
rect 12767 -8602 12865 -8571
rect 12767 -8654 12865 -8602
rect 12767 -8806 12865 -8766
rect 12767 -8840 12865 -8806
rect 12767 -8849 12865 -8840
rect 17875 -7544 17910 -7518
rect 15419 -8601 15517 -8571
rect 15419 -8654 15517 -8601
rect 15419 -8805 15517 -8766
rect 15419 -8839 15517 -8805
rect 15419 -8849 15517 -8839
rect 16436 -8694 16651 -8670
rect 12755 -9445 12850 -9366
rect 15428 -9445 15523 -9366
rect 16436 -8956 16474 -8694
rect 16474 -8956 16611 -8694
rect 16611 -8956 16651 -8694
rect 16436 -8989 16651 -8956
rect 16664 -9431 16832 -9253
rect 9242 -9598 9276 -9564
rect 9500 -9598 9534 -9564
rect 9758 -9598 9792 -9564
rect 10016 -9598 10050 -9564
rect 10274 -9598 10308 -9564
rect 10532 -9598 10566 -9564
rect 10790 -9598 10824 -9564
rect 11048 -9598 11082 -9564
rect 9242 -9908 9276 -9874
rect 9242 -10016 9276 -9982
rect 9500 -9908 9534 -9874
rect 9500 -10016 9534 -9982
rect 9242 -10326 9276 -10292
rect 9242 -10434 9276 -10400
rect 9758 -9908 9792 -9874
rect 9758 -10016 9792 -9982
rect 9500 -10326 9534 -10292
rect 9500 -10434 9534 -10400
rect 9242 -10744 9276 -10710
rect 9242 -10852 9276 -10818
rect 10016 -9908 10050 -9874
rect 10016 -10016 10050 -9982
rect 9758 -10326 9792 -10292
rect 9758 -10434 9792 -10400
rect 9500 -10744 9534 -10710
rect 9500 -10852 9534 -10818
rect 9242 -11162 9276 -11128
rect 9242 -11270 9276 -11236
rect 10274 -9908 10308 -9874
rect 10274 -10016 10308 -9982
rect 10016 -10326 10050 -10292
rect 10016 -10434 10050 -10400
rect 9758 -10744 9792 -10710
rect 9758 -10852 9792 -10818
rect 9500 -11162 9534 -11128
rect 9500 -11270 9534 -11236
rect 9242 -11580 9276 -11546
rect 9242 -11688 9276 -11654
rect 10532 -9908 10566 -9874
rect 10532 -10016 10566 -9982
rect 10274 -10326 10308 -10292
rect 10274 -10434 10308 -10400
rect 10016 -10744 10050 -10710
rect 10016 -10852 10050 -10818
rect 9758 -11162 9792 -11128
rect 9758 -11270 9792 -11236
rect 9500 -11580 9534 -11546
rect 9500 -11688 9534 -11654
rect 9242 -11998 9276 -11964
rect 9242 -12106 9276 -12072
rect 10790 -9908 10824 -9874
rect 10790 -10016 10824 -9982
rect 10532 -10326 10566 -10292
rect 10532 -10434 10566 -10400
rect 10274 -10744 10308 -10710
rect 10274 -10852 10308 -10818
rect 10016 -11162 10050 -11128
rect 10016 -11270 10050 -11236
rect 9758 -11580 9792 -11546
rect 9758 -11688 9792 -11654
rect 9500 -11998 9534 -11964
rect 9500 -12106 9534 -12072
rect 9242 -12416 9276 -12382
rect 11912 -9598 11946 -9564
rect 12170 -9598 12204 -9564
rect 12428 -9598 12462 -9564
rect 12686 -9598 12720 -9564
rect 12944 -9598 12978 -9564
rect 13202 -9598 13236 -9564
rect 13460 -9598 13494 -9564
rect 13718 -9598 13752 -9564
rect 11048 -9908 11082 -9874
rect 11048 -10016 11082 -9982
rect 10790 -10326 10824 -10292
rect 10790 -10434 10824 -10400
rect 10532 -10744 10566 -10710
rect 10532 -10852 10566 -10818
rect 10274 -11162 10308 -11128
rect 10274 -11270 10308 -11236
rect 10016 -11580 10050 -11546
rect 10016 -11688 10050 -11654
rect 9758 -11998 9792 -11964
rect 9758 -12106 9792 -12072
rect 9500 -12416 9534 -12382
rect 11048 -10326 11082 -10292
rect 11048 -10434 11082 -10400
rect 10790 -10744 10824 -10710
rect 10790 -10852 10824 -10818
rect 10532 -11162 10566 -11128
rect 10532 -11270 10566 -11236
rect 10274 -11580 10308 -11546
rect 10274 -11688 10308 -11654
rect 10016 -11998 10050 -11964
rect 10016 -12106 10050 -12072
rect 9758 -12416 9792 -12382
rect 11048 -10744 11082 -10710
rect 11048 -10852 11082 -10818
rect 10790 -11162 10824 -11128
rect 10790 -11270 10824 -11236
rect 10532 -11580 10566 -11546
rect 10532 -11688 10566 -11654
rect 10274 -11998 10308 -11964
rect 10274 -12106 10308 -12072
rect 10016 -12416 10050 -12382
rect 11048 -11162 11082 -11128
rect 11048 -11270 11082 -11236
rect 10790 -11580 10824 -11546
rect 10790 -11688 10824 -11654
rect 10532 -11998 10566 -11964
rect 10532 -12106 10566 -12072
rect 10274 -12416 10308 -12382
rect 11048 -11580 11082 -11546
rect 11048 -11688 11082 -11654
rect 10790 -11998 10824 -11964
rect 10790 -12106 10824 -12072
rect 10532 -12416 10566 -12382
rect 11048 -11998 11082 -11964
rect 11048 -12106 11082 -12072
rect 10790 -12416 10824 -12382
rect 11048 -12416 11082 -12382
rect 11912 -9908 11946 -9874
rect 11912 -10016 11946 -9982
rect 12170 -9908 12204 -9874
rect 12170 -10016 12204 -9982
rect 11912 -10326 11946 -10292
rect 11912 -10434 11946 -10400
rect 12428 -9908 12462 -9874
rect 12428 -10016 12462 -9982
rect 12170 -10326 12204 -10292
rect 12170 -10434 12204 -10400
rect 11912 -10744 11946 -10710
rect 11912 -10852 11946 -10818
rect 12686 -9908 12720 -9874
rect 12686 -10016 12720 -9982
rect 12428 -10326 12462 -10292
rect 12428 -10434 12462 -10400
rect 12170 -10744 12204 -10710
rect 12170 -10852 12204 -10818
rect 11912 -11162 11946 -11128
rect 11912 -11270 11946 -11236
rect 12944 -9908 12978 -9874
rect 12944 -10016 12978 -9982
rect 12686 -10326 12720 -10292
rect 12686 -10434 12720 -10400
rect 12428 -10744 12462 -10710
rect 12428 -10852 12462 -10818
rect 12170 -11162 12204 -11128
rect 12170 -11270 12204 -11236
rect 11912 -11580 11946 -11546
rect 11912 -11688 11946 -11654
rect 13202 -9908 13236 -9874
rect 13202 -10016 13236 -9982
rect 12944 -10326 12978 -10292
rect 12944 -10434 12978 -10400
rect 12686 -10744 12720 -10710
rect 12686 -10852 12720 -10818
rect 12428 -11162 12462 -11128
rect 12428 -11270 12462 -11236
rect 12170 -11580 12204 -11546
rect 12170 -11688 12204 -11654
rect 11912 -11998 11946 -11964
rect 11912 -12106 11946 -12072
rect 13460 -9908 13494 -9874
rect 13460 -10016 13494 -9982
rect 13202 -10326 13236 -10292
rect 13202 -10434 13236 -10400
rect 12944 -10744 12978 -10710
rect 12944 -10852 12978 -10818
rect 12686 -11162 12720 -11128
rect 12686 -11270 12720 -11236
rect 12428 -11580 12462 -11546
rect 12428 -11688 12462 -11654
rect 12170 -11998 12204 -11964
rect 12170 -12106 12204 -12072
rect 11912 -12416 11946 -12382
rect 14575 -9597 14609 -9563
rect 14833 -9597 14867 -9563
rect 15091 -9597 15125 -9563
rect 15349 -9597 15383 -9563
rect 15607 -9597 15641 -9563
rect 15865 -9597 15899 -9563
rect 16123 -9597 16157 -9563
rect 16381 -9597 16415 -9563
rect 13718 -9908 13752 -9874
rect 13718 -10016 13752 -9982
rect 13460 -10326 13494 -10292
rect 13460 -10434 13494 -10400
rect 13202 -10744 13236 -10710
rect 13202 -10852 13236 -10818
rect 12944 -11162 12978 -11128
rect 12944 -11270 12978 -11236
rect 12686 -11580 12720 -11546
rect 12686 -11688 12720 -11654
rect 12428 -11998 12462 -11964
rect 12428 -12106 12462 -12072
rect 12170 -12416 12204 -12382
rect 13718 -10326 13752 -10292
rect 13718 -10434 13752 -10400
rect 13460 -10744 13494 -10710
rect 13460 -10852 13494 -10818
rect 13202 -11162 13236 -11128
rect 13202 -11270 13236 -11236
rect 12944 -11580 12978 -11546
rect 12944 -11688 12978 -11654
rect 12686 -11998 12720 -11964
rect 12686 -12106 12720 -12072
rect 12428 -12416 12462 -12382
rect 13718 -10744 13752 -10710
rect 13718 -10852 13752 -10818
rect 13460 -11162 13494 -11128
rect 13460 -11270 13494 -11236
rect 13202 -11580 13236 -11546
rect 13202 -11688 13236 -11654
rect 12944 -11998 12978 -11964
rect 12944 -12106 12978 -12072
rect 12686 -12416 12720 -12382
rect 13718 -11162 13752 -11128
rect 13718 -11270 13752 -11236
rect 13460 -11580 13494 -11546
rect 13460 -11688 13494 -11654
rect 13202 -11998 13236 -11964
rect 13202 -12106 13236 -12072
rect 12944 -12416 12978 -12382
rect 13718 -11580 13752 -11546
rect 13718 -11688 13752 -11654
rect 13460 -11998 13494 -11964
rect 13460 -12106 13494 -12072
rect 13202 -12416 13236 -12382
rect 13718 -11998 13752 -11964
rect 13718 -12106 13752 -12072
rect 13460 -12416 13494 -12382
rect 13718 -12416 13752 -12382
rect 14575 -9907 14609 -9873
rect 14575 -10015 14609 -9981
rect 14833 -9907 14867 -9873
rect 14833 -10015 14867 -9981
rect 14575 -10325 14609 -10291
rect 14575 -10433 14609 -10399
rect 15091 -9907 15125 -9873
rect 15091 -10015 15125 -9981
rect 14833 -10325 14867 -10291
rect 14833 -10433 14867 -10399
rect 14575 -10743 14609 -10709
rect 14575 -10851 14609 -10817
rect 15349 -9907 15383 -9873
rect 15349 -10015 15383 -9981
rect 15091 -10325 15125 -10291
rect 15091 -10433 15125 -10399
rect 14833 -10743 14867 -10709
rect 14833 -10851 14867 -10817
rect 14575 -11161 14609 -11127
rect 14575 -11269 14609 -11235
rect 15607 -9907 15641 -9873
rect 15607 -10015 15641 -9981
rect 15349 -10325 15383 -10291
rect 15349 -10433 15383 -10399
rect 15091 -10743 15125 -10709
rect 15091 -10851 15125 -10817
rect 14833 -11161 14867 -11127
rect 14833 -11269 14867 -11235
rect 14575 -11579 14609 -11545
rect 14575 -11687 14609 -11653
rect 15865 -9907 15899 -9873
rect 15865 -10015 15899 -9981
rect 15607 -10325 15641 -10291
rect 15607 -10433 15641 -10399
rect 15349 -10743 15383 -10709
rect 15349 -10851 15383 -10817
rect 15091 -11161 15125 -11127
rect 15091 -11269 15125 -11235
rect 14833 -11579 14867 -11545
rect 14833 -11687 14867 -11653
rect 14575 -11997 14609 -11963
rect 14575 -12105 14609 -12071
rect 16123 -9907 16157 -9873
rect 16123 -10015 16157 -9981
rect 15865 -10325 15899 -10291
rect 15865 -10433 15899 -10399
rect 15607 -10743 15641 -10709
rect 15607 -10851 15641 -10817
rect 15349 -11161 15383 -11127
rect 15349 -11269 15383 -11235
rect 15091 -11579 15125 -11545
rect 15091 -11687 15125 -11653
rect 14833 -11997 14867 -11963
rect 14833 -12105 14867 -12071
rect 14575 -12415 14609 -12381
rect 16381 -9907 16415 -9873
rect 16381 -10015 16415 -9981
rect 16123 -10325 16157 -10291
rect 16123 -10433 16157 -10399
rect 15865 -10743 15899 -10709
rect 15865 -10851 15899 -10817
rect 15607 -11161 15641 -11127
rect 15607 -11269 15641 -11235
rect 15349 -11579 15383 -11545
rect 15349 -11687 15383 -11653
rect 15091 -11997 15125 -11963
rect 15091 -12105 15125 -12071
rect 14833 -12415 14867 -12381
rect 16381 -10325 16415 -10291
rect 16381 -10433 16415 -10399
rect 16123 -10743 16157 -10709
rect 16123 -10851 16157 -10817
rect 15865 -11161 15899 -11127
rect 15865 -11269 15899 -11235
rect 15607 -11579 15641 -11545
rect 15607 -11687 15641 -11653
rect 15349 -11997 15383 -11963
rect 15349 -12105 15383 -12071
rect 15091 -12415 15125 -12381
rect 16381 -10743 16415 -10709
rect 16381 -10851 16415 -10817
rect 16123 -11161 16157 -11127
rect 16123 -11269 16157 -11235
rect 15865 -11579 15899 -11545
rect 15865 -11687 15899 -11653
rect 15607 -11997 15641 -11963
rect 15607 -12105 15641 -12071
rect 15349 -12415 15383 -12381
rect 16381 -11161 16415 -11127
rect 16381 -11269 16415 -11235
rect 16123 -11579 16157 -11545
rect 16123 -11687 16157 -11653
rect 15865 -11997 15899 -11963
rect 15865 -12105 15899 -12071
rect 15607 -12415 15641 -12381
rect 16381 -11579 16415 -11545
rect 16381 -11687 16415 -11653
rect 16123 -11997 16157 -11963
rect 16123 -12105 16157 -12071
rect 15865 -12415 15899 -12381
rect 16381 -11997 16415 -11963
rect 16381 -12105 16415 -12071
rect 16123 -12415 16157 -12381
rect 16381 -12415 16415 -12381
rect 10137 -12758 10142 -12724
rect 10142 -12758 10176 -12724
rect 10176 -12758 10187 -12724
rect 10137 -12764 10187 -12758
rect 12807 -12758 12812 -12724
rect 12812 -12758 12846 -12724
rect 12846 -12758 12857 -12724
rect 12807 -12764 12857 -12758
rect 10140 -13034 10178 -13031
rect 10140 -13068 10142 -13034
rect 10142 -13068 10176 -13034
rect 10176 -13068 10178 -13034
rect 10140 -13071 10178 -13068
rect 15470 -12757 15475 -12723
rect 15475 -12757 15509 -12723
rect 15509 -12757 15520 -12723
rect 15470 -12763 15520 -12757
rect 12810 -13034 12848 -13031
rect 12810 -13068 12812 -13034
rect 12812 -13068 12846 -13034
rect 12846 -13068 12848 -13034
rect 12810 -13071 12848 -13068
rect 15472 -13033 15510 -13031
rect 15472 -13067 15475 -13033
rect 15475 -13067 15509 -13033
rect 15509 -13067 15510 -13033
rect 15472 -13071 15510 -13067
rect 9970 -13267 10076 -13161
rect 12634 -13267 12740 -13161
rect 15296 -13267 15402 -13161
rect 8991 -14241 9174 -14220
rect 8991 -14503 9014 -14241
rect 9014 -14503 9151 -14241
rect 9151 -14503 9174 -14241
rect 10093 -14250 10173 -14249
rect 10093 -14284 10173 -14250
rect 10093 -14310 10173 -14284
rect 10092 -14488 10172 -14470
rect 8991 -14525 9174 -14503
rect 10092 -14522 10172 -14488
rect 10092 -14531 10172 -14522
rect 12748 -14284 12846 -14253
rect 12748 -14336 12846 -14284
rect 15423 -14283 15521 -14253
rect 15423 -14336 15521 -14283
rect 12748 -14488 12846 -14448
rect 12748 -14522 12846 -14488
rect 12748 -14531 12846 -14522
rect 8856 -15171 9014 -15007
rect 15423 -14487 15521 -14448
rect 15423 -14521 15521 -14487
rect 15423 -14531 15521 -14521
rect 11562 -15191 11680 -15057
rect 9242 -15315 9276 -15281
rect 9500 -15315 9534 -15281
rect 9758 -15315 9792 -15281
rect 10016 -15315 10050 -15281
rect 10274 -15315 10308 -15281
rect 10532 -15315 10566 -15281
rect 10790 -15315 10824 -15281
rect 11048 -15315 11082 -15281
rect 9242 -15625 9276 -15591
rect 9242 -15733 9276 -15699
rect 9500 -15625 9534 -15591
rect 9500 -15733 9534 -15699
rect 9242 -16043 9276 -16009
rect 9242 -16151 9276 -16117
rect 9758 -15625 9792 -15591
rect 9758 -15733 9792 -15699
rect 9500 -16043 9534 -16009
rect 9500 -16151 9534 -16117
rect 9242 -16461 9276 -16427
rect 9242 -16569 9276 -16535
rect 10016 -15625 10050 -15591
rect 10016 -15733 10050 -15699
rect 9758 -16043 9792 -16009
rect 9758 -16151 9792 -16117
rect 9500 -16461 9534 -16427
rect 9500 -16569 9534 -16535
rect 9242 -16879 9276 -16845
rect 9242 -16987 9276 -16953
rect 10274 -15625 10308 -15591
rect 10274 -15733 10308 -15699
rect 10016 -16043 10050 -16009
rect 10016 -16151 10050 -16117
rect 9758 -16461 9792 -16427
rect 9758 -16569 9792 -16535
rect 9500 -16879 9534 -16845
rect 9500 -16987 9534 -16953
rect 9242 -17297 9276 -17263
rect 9242 -17405 9276 -17371
rect 10532 -15625 10566 -15591
rect 10532 -15733 10566 -15699
rect 10274 -16043 10308 -16009
rect 10274 -16151 10308 -16117
rect 10016 -16461 10050 -16427
rect 10016 -16569 10050 -16535
rect 9758 -16879 9792 -16845
rect 9758 -16987 9792 -16953
rect 9500 -17297 9534 -17263
rect 9500 -17405 9534 -17371
rect 9242 -17715 9276 -17681
rect 9242 -17823 9276 -17789
rect 14168 -15191 14280 -15067
rect 11912 -15315 11946 -15281
rect 12170 -15315 12204 -15281
rect 12428 -15315 12462 -15281
rect 12686 -15315 12720 -15281
rect 12944 -15315 12978 -15281
rect 13202 -15315 13236 -15281
rect 13460 -15315 13494 -15281
rect 13718 -15315 13752 -15281
rect 10790 -15625 10824 -15591
rect 10790 -15733 10824 -15699
rect 10532 -16043 10566 -16009
rect 10532 -16151 10566 -16117
rect 10274 -16461 10308 -16427
rect 10274 -16569 10308 -16535
rect 10016 -16879 10050 -16845
rect 10016 -16987 10050 -16953
rect 9758 -17297 9792 -17263
rect 9758 -17405 9792 -17371
rect 9500 -17715 9534 -17681
rect 9500 -17823 9534 -17789
rect 9242 -18133 9276 -18099
rect 11048 -15625 11082 -15591
rect 11048 -15733 11082 -15699
rect 10790 -16043 10824 -16009
rect 10790 -16151 10824 -16117
rect 10532 -16461 10566 -16427
rect 10532 -16569 10566 -16535
rect 10274 -16879 10308 -16845
rect 10274 -16987 10308 -16953
rect 10016 -17297 10050 -17263
rect 10016 -17405 10050 -17371
rect 9758 -17715 9792 -17681
rect 9758 -17823 9792 -17789
rect 9500 -18133 9534 -18099
rect 11048 -16043 11082 -16009
rect 11048 -16151 11082 -16117
rect 10790 -16461 10824 -16427
rect 10790 -16569 10824 -16535
rect 10532 -16879 10566 -16845
rect 10532 -16987 10566 -16953
rect 10274 -17297 10308 -17263
rect 10274 -17405 10308 -17371
rect 10016 -17715 10050 -17681
rect 10016 -17823 10050 -17789
rect 9758 -18133 9792 -18099
rect 11048 -16461 11082 -16427
rect 11048 -16569 11082 -16535
rect 10790 -16879 10824 -16845
rect 10790 -16987 10824 -16953
rect 10532 -17297 10566 -17263
rect 10532 -17405 10566 -17371
rect 10274 -17715 10308 -17681
rect 10274 -17823 10308 -17789
rect 10016 -18133 10050 -18099
rect 11048 -16879 11082 -16845
rect 11048 -16987 11082 -16953
rect 10790 -17297 10824 -17263
rect 10790 -17405 10824 -17371
rect 10532 -17715 10566 -17681
rect 10532 -17823 10566 -17789
rect 10274 -18133 10308 -18099
rect 11048 -17297 11082 -17263
rect 11048 -17405 11082 -17371
rect 10790 -17715 10824 -17681
rect 10790 -17823 10824 -17789
rect 10532 -18133 10566 -18099
rect 11048 -17715 11082 -17681
rect 11048 -17823 11082 -17789
rect 10790 -18133 10824 -18099
rect 11912 -15625 11946 -15591
rect 11912 -15733 11946 -15699
rect 12170 -15625 12204 -15591
rect 12170 -15733 12204 -15699
rect 11912 -16043 11946 -16009
rect 11912 -16151 11946 -16117
rect 12428 -15625 12462 -15591
rect 12428 -15733 12462 -15699
rect 12170 -16043 12204 -16009
rect 12170 -16151 12204 -16117
rect 11912 -16461 11946 -16427
rect 11912 -16569 11946 -16535
rect 12686 -15625 12720 -15591
rect 12686 -15733 12720 -15699
rect 12428 -16043 12462 -16009
rect 12428 -16151 12462 -16117
rect 12170 -16461 12204 -16427
rect 12170 -16569 12204 -16535
rect 11912 -16879 11946 -16845
rect 11912 -16987 11946 -16953
rect 12944 -15625 12978 -15591
rect 12944 -15733 12978 -15699
rect 12686 -16043 12720 -16009
rect 12686 -16151 12720 -16117
rect 12428 -16461 12462 -16427
rect 12428 -16569 12462 -16535
rect 12170 -16879 12204 -16845
rect 12170 -16987 12204 -16953
rect 11912 -17297 11946 -17263
rect 11912 -17405 11946 -17371
rect 13202 -15625 13236 -15591
rect 13202 -15733 13236 -15699
rect 12944 -16043 12978 -16009
rect 12944 -16151 12978 -16117
rect 12686 -16461 12720 -16427
rect 12686 -16569 12720 -16535
rect 12428 -16879 12462 -16845
rect 12428 -16987 12462 -16953
rect 12170 -17297 12204 -17263
rect 12170 -17405 12204 -17371
rect 11912 -17715 11946 -17681
rect 11912 -17823 11946 -17789
rect 11048 -18133 11082 -18099
rect 14575 -15314 14609 -15280
rect 14833 -15314 14867 -15280
rect 15091 -15314 15125 -15280
rect 15349 -15314 15383 -15280
rect 15607 -15314 15641 -15280
rect 15865 -15314 15899 -15280
rect 16123 -15314 16157 -15280
rect 16381 -15314 16415 -15280
rect 13460 -15625 13494 -15591
rect 13460 -15733 13494 -15699
rect 13202 -16043 13236 -16009
rect 13202 -16151 13236 -16117
rect 12944 -16461 12978 -16427
rect 12944 -16569 12978 -16535
rect 12686 -16879 12720 -16845
rect 12686 -16987 12720 -16953
rect 12428 -17297 12462 -17263
rect 12428 -17405 12462 -17371
rect 12170 -17715 12204 -17681
rect 12170 -17823 12204 -17789
rect 11912 -18133 11946 -18099
rect 13718 -15625 13752 -15591
rect 13718 -15733 13752 -15699
rect 13460 -16043 13494 -16009
rect 13460 -16151 13494 -16117
rect 13202 -16461 13236 -16427
rect 13202 -16569 13236 -16535
rect 12944 -16879 12978 -16845
rect 12944 -16987 12978 -16953
rect 12686 -17297 12720 -17263
rect 12686 -17405 12720 -17371
rect 12428 -17715 12462 -17681
rect 12428 -17823 12462 -17789
rect 12170 -18133 12204 -18099
rect 13718 -16043 13752 -16009
rect 13718 -16151 13752 -16117
rect 13460 -16461 13494 -16427
rect 13460 -16569 13494 -16535
rect 13202 -16879 13236 -16845
rect 13202 -16987 13236 -16953
rect 12944 -17297 12978 -17263
rect 12944 -17405 12978 -17371
rect 12686 -17715 12720 -17681
rect 12686 -17823 12720 -17789
rect 12428 -18133 12462 -18099
rect 13718 -16461 13752 -16427
rect 13718 -16569 13752 -16535
rect 13460 -16879 13494 -16845
rect 13460 -16987 13494 -16953
rect 13202 -17297 13236 -17263
rect 13202 -17405 13236 -17371
rect 12944 -17715 12978 -17681
rect 12944 -17823 12978 -17789
rect 12686 -18133 12720 -18099
rect 13718 -16879 13752 -16845
rect 13718 -16987 13752 -16953
rect 13460 -17297 13494 -17263
rect 13460 -17405 13494 -17371
rect 13202 -17715 13236 -17681
rect 13202 -17823 13236 -17789
rect 12944 -18133 12978 -18099
rect 13718 -17297 13752 -17263
rect 13718 -17405 13752 -17371
rect 13460 -17715 13494 -17681
rect 13460 -17823 13494 -17789
rect 13202 -18133 13236 -18099
rect 13718 -17715 13752 -17681
rect 13718 -17823 13752 -17789
rect 13460 -18133 13494 -18099
rect 14575 -15624 14609 -15590
rect 14575 -15732 14609 -15698
rect 14833 -15624 14867 -15590
rect 14833 -15732 14867 -15698
rect 14575 -16042 14609 -16008
rect 14575 -16150 14609 -16116
rect 15091 -15624 15125 -15590
rect 15091 -15732 15125 -15698
rect 14833 -16042 14867 -16008
rect 14833 -16150 14867 -16116
rect 14575 -16460 14609 -16426
rect 14575 -16568 14609 -16534
rect 15349 -15624 15383 -15590
rect 15349 -15732 15383 -15698
rect 15091 -16042 15125 -16008
rect 15091 -16150 15125 -16116
rect 14833 -16460 14867 -16426
rect 14833 -16568 14867 -16534
rect 14575 -16878 14609 -16844
rect 14575 -16986 14609 -16952
rect 15607 -15624 15641 -15590
rect 15607 -15732 15641 -15698
rect 15349 -16042 15383 -16008
rect 15349 -16150 15383 -16116
rect 15091 -16460 15125 -16426
rect 15091 -16568 15125 -16534
rect 14833 -16878 14867 -16844
rect 14833 -16986 14867 -16952
rect 14575 -17296 14609 -17262
rect 14575 -17404 14609 -17370
rect 15865 -15624 15899 -15590
rect 15865 -15732 15899 -15698
rect 15607 -16042 15641 -16008
rect 15607 -16150 15641 -16116
rect 15349 -16460 15383 -16426
rect 15349 -16568 15383 -16534
rect 15091 -16878 15125 -16844
rect 15091 -16986 15125 -16952
rect 14833 -17296 14867 -17262
rect 14833 -17404 14867 -17370
rect 14575 -17714 14609 -17680
rect 14575 -17822 14609 -17788
rect 13718 -18133 13752 -18099
rect 16123 -15624 16157 -15590
rect 16123 -15732 16157 -15698
rect 15865 -16042 15899 -16008
rect 15865 -16150 15899 -16116
rect 15607 -16460 15641 -16426
rect 15607 -16568 15641 -16534
rect 15349 -16878 15383 -16844
rect 15349 -16986 15383 -16952
rect 15091 -17296 15125 -17262
rect 15091 -17404 15125 -17370
rect 14833 -17714 14867 -17680
rect 14833 -17822 14867 -17788
rect 14575 -18132 14609 -18098
rect 16381 -15624 16415 -15590
rect 16381 -15732 16415 -15698
rect 16123 -16042 16157 -16008
rect 16123 -16150 16157 -16116
rect 15865 -16460 15899 -16426
rect 15865 -16568 15899 -16534
rect 15607 -16878 15641 -16844
rect 15607 -16986 15641 -16952
rect 15349 -17296 15383 -17262
rect 15349 -17404 15383 -17370
rect 15091 -17714 15125 -17680
rect 15091 -17822 15125 -17788
rect 14833 -18132 14867 -18098
rect 16381 -16042 16415 -16008
rect 16381 -16150 16415 -16116
rect 16123 -16460 16157 -16426
rect 16123 -16568 16157 -16534
rect 15865 -16878 15899 -16844
rect 15865 -16986 15899 -16952
rect 15607 -17296 15641 -17262
rect 15607 -17404 15641 -17370
rect 15349 -17714 15383 -17680
rect 15349 -17822 15383 -17788
rect 15091 -18132 15125 -18098
rect 16381 -16460 16415 -16426
rect 16381 -16568 16415 -16534
rect 16123 -16878 16157 -16844
rect 16123 -16986 16157 -16952
rect 15865 -17296 15899 -17262
rect 15865 -17404 15899 -17370
rect 15607 -17714 15641 -17680
rect 15607 -17822 15641 -17788
rect 15349 -18132 15383 -18098
rect 16381 -16878 16415 -16844
rect 16381 -16986 16415 -16952
rect 16123 -17296 16157 -17262
rect 16123 -17404 16157 -17370
rect 15865 -17714 15899 -17680
rect 15865 -17822 15899 -17788
rect 15607 -18132 15641 -18098
rect 16381 -17296 16415 -17262
rect 16381 -17404 16415 -17370
rect 16123 -17714 16157 -17680
rect 16123 -17822 16157 -17788
rect 15865 -18132 15899 -18098
rect 16381 -17714 16415 -17680
rect 16381 -17822 16415 -17788
rect 16123 -18132 16157 -18098
rect 16381 -18132 16415 -18098
rect 10137 -18475 10142 -18441
rect 10142 -18475 10176 -18441
rect 10176 -18475 10187 -18441
rect 10137 -18481 10187 -18475
rect 12807 -18475 12812 -18441
rect 12812 -18475 12846 -18441
rect 12846 -18475 12857 -18441
rect 12807 -18481 12857 -18475
rect 10140 -18751 10180 -18749
rect 10140 -18785 10142 -18751
rect 10142 -18785 10176 -18751
rect 10176 -18785 10180 -18751
rect 10140 -18787 10180 -18785
rect 15470 -18474 15475 -18440
rect 15475 -18474 15509 -18440
rect 15509 -18474 15520 -18440
rect 15470 -18480 15520 -18474
rect 12810 -18751 12850 -18749
rect 12810 -18785 12812 -18751
rect 12812 -18785 12846 -18751
rect 12846 -18785 12850 -18751
rect 12810 -18787 12850 -18785
rect 15470 -18750 15512 -18747
rect 15470 -18784 15475 -18750
rect 15475 -18784 15509 -18750
rect 15509 -18784 15512 -18750
rect 15470 -18789 15512 -18784
rect 9964 -18885 10070 -18880
rect 9964 -18979 9972 -18885
rect 9972 -18979 10064 -18885
rect 10064 -18979 10070 -18885
rect 12640 -18979 12732 -18885
rect 15306 -18979 15398 -18885
rect 9964 -18986 10070 -18979
rect 8970 -20124 9113 -20123
rect 8970 -20385 8973 -20124
rect 8973 -20385 9109 -20124
rect 9109 -20385 9113 -20124
rect 8970 -20387 9113 -20385
rect 10093 -20175 10173 -20174
rect 10093 -20209 10173 -20175
rect 10093 -20235 10173 -20209
rect 10094 -20413 10174 -20395
rect 10094 -20447 10174 -20413
rect 10094 -20456 10174 -20447
rect 12767 -20209 12865 -20178
rect 12767 -20261 12865 -20209
rect 12767 -20413 12865 -20373
rect 12767 -20447 12865 -20413
rect 12767 -20456 12865 -20447
rect 16698 -19575 16732 -19541
rect 17088 -19577 17122 -19543
rect 16247 -19579 16449 -19577
rect 16247 -19892 16248 -19579
rect 16248 -19892 16449 -19579
rect 16887 -19751 16958 -19747
rect 16887 -19813 16900 -19751
rect 16900 -19813 16956 -19751
rect 16956 -19813 16958 -19751
rect 16887 -19819 16958 -19813
rect 16698 -20039 16732 -20005
rect 17088 -20041 17122 -20007
rect 15419 -20208 15517 -20178
rect 15419 -20261 15517 -20208
rect 16848 -20219 16902 -20181
rect 17236 -20227 17284 -20183
rect 15419 -20412 15517 -20373
rect 15419 -20446 15517 -20412
rect 15419 -20456 15517 -20446
rect 16702 -20371 16736 -20337
rect 17092 -20371 17126 -20337
rect 16523 -20487 16526 -20415
rect 16526 -20487 16570 -20415
rect 16570 -20487 16579 -20415
rect 16523 -20488 16579 -20487
rect 16915 -20487 16916 -20415
rect 16916 -20487 16960 -20415
rect 16960 -20487 16961 -20415
rect 16915 -20488 16961 -20487
rect 16702 -20565 16736 -20531
rect 17092 -20565 17126 -20531
rect 12755 -21066 12850 -20987
rect 15428 -21066 15523 -20987
rect 16542 -21031 16792 -20741
rect 17164 -21033 17414 -20743
rect 9242 -21219 9276 -21185
rect 9500 -21219 9534 -21185
rect 9758 -21219 9792 -21185
rect 10016 -21219 10050 -21185
rect 10274 -21219 10308 -21185
rect 10532 -21219 10566 -21185
rect 10790 -21219 10824 -21185
rect 11048 -21219 11082 -21185
rect 9242 -21529 9276 -21495
rect 9242 -21637 9276 -21603
rect 9500 -21529 9534 -21495
rect 9500 -21637 9534 -21603
rect 9242 -21947 9276 -21913
rect 9242 -22055 9276 -22021
rect 9758 -21529 9792 -21495
rect 9758 -21637 9792 -21603
rect 9500 -21947 9534 -21913
rect 9500 -22055 9534 -22021
rect 9242 -22365 9276 -22331
rect 9242 -22473 9276 -22439
rect 10016 -21529 10050 -21495
rect 10016 -21637 10050 -21603
rect 9758 -21947 9792 -21913
rect 9758 -22055 9792 -22021
rect 9500 -22365 9534 -22331
rect 9500 -22473 9534 -22439
rect 9242 -22783 9276 -22749
rect 9242 -22891 9276 -22857
rect 10274 -21529 10308 -21495
rect 10274 -21637 10308 -21603
rect 10016 -21947 10050 -21913
rect 10016 -22055 10050 -22021
rect 9758 -22365 9792 -22331
rect 9758 -22473 9792 -22439
rect 9500 -22783 9534 -22749
rect 9500 -22891 9534 -22857
rect 9242 -23201 9276 -23167
rect 9242 -23309 9276 -23275
rect 10532 -21529 10566 -21495
rect 10532 -21637 10566 -21603
rect 10274 -21947 10308 -21913
rect 10274 -22055 10308 -22021
rect 10016 -22365 10050 -22331
rect 10016 -22473 10050 -22439
rect 9758 -22783 9792 -22749
rect 9758 -22891 9792 -22857
rect 9500 -23201 9534 -23167
rect 9500 -23309 9534 -23275
rect 9242 -23619 9276 -23585
rect 9242 -23727 9276 -23693
rect 10790 -21529 10824 -21495
rect 10790 -21637 10824 -21603
rect 10532 -21947 10566 -21913
rect 10532 -22055 10566 -22021
rect 10274 -22365 10308 -22331
rect 10274 -22473 10308 -22439
rect 10016 -22783 10050 -22749
rect 10016 -22891 10050 -22857
rect 9758 -23201 9792 -23167
rect 9758 -23309 9792 -23275
rect 9500 -23619 9534 -23585
rect 9500 -23727 9534 -23693
rect 9242 -24037 9276 -24003
rect 11912 -21219 11946 -21185
rect 12170 -21219 12204 -21185
rect 12428 -21219 12462 -21185
rect 12686 -21219 12720 -21185
rect 12944 -21219 12978 -21185
rect 13202 -21219 13236 -21185
rect 13460 -21219 13494 -21185
rect 13718 -21219 13752 -21185
rect 11048 -21529 11082 -21495
rect 11048 -21637 11082 -21603
rect 10790 -21947 10824 -21913
rect 10790 -22055 10824 -22021
rect 10532 -22365 10566 -22331
rect 10532 -22473 10566 -22439
rect 10274 -22783 10308 -22749
rect 10274 -22891 10308 -22857
rect 10016 -23201 10050 -23167
rect 10016 -23309 10050 -23275
rect 9758 -23619 9792 -23585
rect 9758 -23727 9792 -23693
rect 9500 -24037 9534 -24003
rect 11048 -21947 11082 -21913
rect 11048 -22055 11082 -22021
rect 10790 -22365 10824 -22331
rect 10790 -22473 10824 -22439
rect 10532 -22783 10566 -22749
rect 10532 -22891 10566 -22857
rect 10274 -23201 10308 -23167
rect 10274 -23309 10308 -23275
rect 10016 -23619 10050 -23585
rect 10016 -23727 10050 -23693
rect 9758 -24037 9792 -24003
rect 11048 -22365 11082 -22331
rect 11048 -22473 11082 -22439
rect 10790 -22783 10824 -22749
rect 10790 -22891 10824 -22857
rect 10532 -23201 10566 -23167
rect 10532 -23309 10566 -23275
rect 10274 -23619 10308 -23585
rect 10274 -23727 10308 -23693
rect 10016 -24037 10050 -24003
rect 11048 -22783 11082 -22749
rect 11048 -22891 11082 -22857
rect 10790 -23201 10824 -23167
rect 10790 -23309 10824 -23275
rect 10532 -23619 10566 -23585
rect 10532 -23727 10566 -23693
rect 10274 -24037 10308 -24003
rect 11048 -23201 11082 -23167
rect 11048 -23309 11082 -23275
rect 10790 -23619 10824 -23585
rect 10790 -23727 10824 -23693
rect 10532 -24037 10566 -24003
rect 11048 -23619 11082 -23585
rect 11048 -23727 11082 -23693
rect 10790 -24037 10824 -24003
rect 11048 -24037 11082 -24003
rect 11912 -21529 11946 -21495
rect 11912 -21637 11946 -21603
rect 12170 -21529 12204 -21495
rect 12170 -21637 12204 -21603
rect 11912 -21947 11946 -21913
rect 11912 -22055 11946 -22021
rect 12428 -21529 12462 -21495
rect 12428 -21637 12462 -21603
rect 12170 -21947 12204 -21913
rect 12170 -22055 12204 -22021
rect 11912 -22365 11946 -22331
rect 11912 -22473 11946 -22439
rect 12686 -21529 12720 -21495
rect 12686 -21637 12720 -21603
rect 12428 -21947 12462 -21913
rect 12428 -22055 12462 -22021
rect 12170 -22365 12204 -22331
rect 12170 -22473 12204 -22439
rect 11912 -22783 11946 -22749
rect 11912 -22891 11946 -22857
rect 12944 -21529 12978 -21495
rect 12944 -21637 12978 -21603
rect 12686 -21947 12720 -21913
rect 12686 -22055 12720 -22021
rect 12428 -22365 12462 -22331
rect 12428 -22473 12462 -22439
rect 12170 -22783 12204 -22749
rect 12170 -22891 12204 -22857
rect 11912 -23201 11946 -23167
rect 11912 -23309 11946 -23275
rect 13202 -21529 13236 -21495
rect 13202 -21637 13236 -21603
rect 12944 -21947 12978 -21913
rect 12944 -22055 12978 -22021
rect 12686 -22365 12720 -22331
rect 12686 -22473 12720 -22439
rect 12428 -22783 12462 -22749
rect 12428 -22891 12462 -22857
rect 12170 -23201 12204 -23167
rect 12170 -23309 12204 -23275
rect 11912 -23619 11946 -23585
rect 11912 -23727 11946 -23693
rect 13460 -21529 13494 -21495
rect 13460 -21637 13494 -21603
rect 13202 -21947 13236 -21913
rect 13202 -22055 13236 -22021
rect 12944 -22365 12978 -22331
rect 12944 -22473 12978 -22439
rect 12686 -22783 12720 -22749
rect 12686 -22891 12720 -22857
rect 12428 -23201 12462 -23167
rect 12428 -23309 12462 -23275
rect 12170 -23619 12204 -23585
rect 12170 -23727 12204 -23693
rect 11912 -24037 11946 -24003
rect 14575 -21218 14609 -21184
rect 14833 -21218 14867 -21184
rect 15091 -21218 15125 -21184
rect 15349 -21218 15383 -21184
rect 15607 -21218 15641 -21184
rect 15865 -21218 15899 -21184
rect 16123 -21218 16157 -21184
rect 16381 -21218 16415 -21184
rect 13718 -21529 13752 -21495
rect 13718 -21637 13752 -21603
rect 13460 -21947 13494 -21913
rect 13460 -22055 13494 -22021
rect 13202 -22365 13236 -22331
rect 13202 -22473 13236 -22439
rect 12944 -22783 12978 -22749
rect 12944 -22891 12978 -22857
rect 12686 -23201 12720 -23167
rect 12686 -23309 12720 -23275
rect 12428 -23619 12462 -23585
rect 12428 -23727 12462 -23693
rect 12170 -24037 12204 -24003
rect 13718 -21947 13752 -21913
rect 13718 -22055 13752 -22021
rect 13460 -22365 13494 -22331
rect 13460 -22473 13494 -22439
rect 13202 -22783 13236 -22749
rect 13202 -22891 13236 -22857
rect 12944 -23201 12978 -23167
rect 12944 -23309 12978 -23275
rect 12686 -23619 12720 -23585
rect 12686 -23727 12720 -23693
rect 12428 -24037 12462 -24003
rect 13718 -22365 13752 -22331
rect 13718 -22473 13752 -22439
rect 13460 -22783 13494 -22749
rect 13460 -22891 13494 -22857
rect 13202 -23201 13236 -23167
rect 13202 -23309 13236 -23275
rect 12944 -23619 12978 -23585
rect 12944 -23727 12978 -23693
rect 12686 -24037 12720 -24003
rect 13718 -22783 13752 -22749
rect 13718 -22891 13752 -22857
rect 13460 -23201 13494 -23167
rect 13460 -23309 13494 -23275
rect 13202 -23619 13236 -23585
rect 13202 -23727 13236 -23693
rect 12944 -24037 12978 -24003
rect 13718 -23201 13752 -23167
rect 13718 -23309 13752 -23275
rect 13460 -23619 13494 -23585
rect 13460 -23727 13494 -23693
rect 13202 -24037 13236 -24003
rect 13718 -23619 13752 -23585
rect 13718 -23727 13752 -23693
rect 13460 -24037 13494 -24003
rect 13718 -24037 13752 -24003
rect 14575 -21528 14609 -21494
rect 14575 -21636 14609 -21602
rect 14833 -21528 14867 -21494
rect 14833 -21636 14867 -21602
rect 14575 -21946 14609 -21912
rect 14575 -22054 14609 -22020
rect 15091 -21528 15125 -21494
rect 15091 -21636 15125 -21602
rect 14833 -21946 14867 -21912
rect 14833 -22054 14867 -22020
rect 14575 -22364 14609 -22330
rect 14575 -22472 14609 -22438
rect 15349 -21528 15383 -21494
rect 15349 -21636 15383 -21602
rect 15091 -21946 15125 -21912
rect 15091 -22054 15125 -22020
rect 14833 -22364 14867 -22330
rect 14833 -22472 14867 -22438
rect 14575 -22782 14609 -22748
rect 14575 -22890 14609 -22856
rect 15607 -21528 15641 -21494
rect 15607 -21636 15641 -21602
rect 15349 -21946 15383 -21912
rect 15349 -22054 15383 -22020
rect 15091 -22364 15125 -22330
rect 15091 -22472 15125 -22438
rect 14833 -22782 14867 -22748
rect 14833 -22890 14867 -22856
rect 14575 -23200 14609 -23166
rect 14575 -23308 14609 -23274
rect 15865 -21528 15899 -21494
rect 15865 -21636 15899 -21602
rect 15607 -21946 15641 -21912
rect 15607 -22054 15641 -22020
rect 15349 -22364 15383 -22330
rect 15349 -22472 15383 -22438
rect 15091 -22782 15125 -22748
rect 15091 -22890 15125 -22856
rect 14833 -23200 14867 -23166
rect 14833 -23308 14867 -23274
rect 14575 -23618 14609 -23584
rect 14575 -23726 14609 -23692
rect 16123 -21528 16157 -21494
rect 16123 -21636 16157 -21602
rect 15865 -21946 15899 -21912
rect 15865 -22054 15899 -22020
rect 15607 -22364 15641 -22330
rect 15607 -22472 15641 -22438
rect 15349 -22782 15383 -22748
rect 15349 -22890 15383 -22856
rect 15091 -23200 15125 -23166
rect 15091 -23308 15125 -23274
rect 14833 -23618 14867 -23584
rect 14833 -23726 14867 -23692
rect 14575 -24036 14609 -24002
rect 16381 -21528 16415 -21494
rect 16381 -21636 16415 -21602
rect 16123 -21946 16157 -21912
rect 16123 -22054 16157 -22020
rect 15865 -22364 15899 -22330
rect 15865 -22472 15899 -22438
rect 15607 -22782 15641 -22748
rect 15607 -22890 15641 -22856
rect 15349 -23200 15383 -23166
rect 15349 -23308 15383 -23274
rect 15091 -23618 15125 -23584
rect 15091 -23726 15125 -23692
rect 14833 -24036 14867 -24002
rect 16381 -21946 16415 -21912
rect 16381 -22054 16415 -22020
rect 16123 -22364 16157 -22330
rect 16123 -22472 16157 -22438
rect 15865 -22782 15899 -22748
rect 15865 -22890 15899 -22856
rect 15607 -23200 15641 -23166
rect 15607 -23308 15641 -23274
rect 15349 -23618 15383 -23584
rect 15349 -23726 15383 -23692
rect 15091 -24036 15125 -24002
rect 16381 -22364 16415 -22330
rect 16381 -22472 16415 -22438
rect 16123 -22782 16157 -22748
rect 16123 -22890 16157 -22856
rect 15865 -23200 15899 -23166
rect 15865 -23308 15899 -23274
rect 15607 -23618 15641 -23584
rect 15607 -23726 15641 -23692
rect 15349 -24036 15383 -24002
rect 16381 -22782 16415 -22748
rect 16381 -22890 16415 -22856
rect 16123 -23200 16157 -23166
rect 16123 -23308 16157 -23274
rect 15865 -23618 15899 -23584
rect 15865 -23726 15899 -23692
rect 15607 -24036 15641 -24002
rect 16381 -23200 16415 -23166
rect 16381 -23308 16415 -23274
rect 16123 -23618 16157 -23584
rect 16123 -23726 16157 -23692
rect 15865 -24036 15899 -24002
rect 16381 -23618 16415 -23584
rect 16381 -23726 16415 -23692
rect 16123 -24036 16157 -24002
rect 16381 -24036 16415 -24002
rect 10137 -24379 10142 -24345
rect 10142 -24379 10176 -24345
rect 10176 -24379 10187 -24345
rect 10137 -24385 10187 -24379
rect 12807 -24379 12812 -24345
rect 12812 -24379 12846 -24345
rect 12846 -24379 12857 -24345
rect 12807 -24385 12857 -24379
rect 10138 -24655 10178 -24654
rect 10138 -24689 10142 -24655
rect 10142 -24689 10176 -24655
rect 10176 -24689 10178 -24655
rect 10138 -24690 10178 -24689
rect 15470 -24378 15475 -24344
rect 15475 -24378 15509 -24344
rect 15509 -24378 15520 -24344
rect 15470 -24384 15520 -24378
rect 12808 -24655 12852 -24651
rect 12808 -24689 12812 -24655
rect 12812 -24689 12846 -24655
rect 12846 -24689 12852 -24655
rect 12808 -24694 12852 -24689
rect 15470 -24654 15514 -24650
rect 15470 -24688 15475 -24654
rect 15475 -24688 15509 -24654
rect 15509 -24688 15514 -24654
rect 15470 -24692 15514 -24688
rect 9972 -24875 10064 -24781
rect 12642 -24875 12734 -24781
rect 15308 -24875 15400 -24781
rect 7798 -25771 7834 -25711
rect 17875 -25710 17876 -7544
rect 17876 -25710 17910 -7544
rect 17990 -9010 18024 -7634
rect 21419 -7544 21454 -7518
rect 17990 -10520 18024 -9144
rect 17990 -12030 18024 -10654
rect 17990 -13540 18024 -12164
rect 17990 -15050 18024 -13674
rect 17990 -16560 18024 -15184
rect 17990 -18070 18024 -16694
rect 17990 -19580 18024 -18204
rect 17990 -21090 18024 -19714
rect 17990 -22600 18024 -21224
rect 17990 -24110 18024 -22734
rect 17990 -25620 18024 -24244
rect 17875 -25764 17910 -25710
rect 19648 -9010 19682 -7634
rect 19648 -10520 19682 -9144
rect 19648 -12030 19682 -10654
rect 19648 -13540 19682 -12164
rect 19648 -15050 19682 -13674
rect 19648 -16560 19682 -15184
rect 19648 -18070 19682 -16694
rect 19648 -19580 19682 -18204
rect 19648 -21090 19682 -19714
rect 19648 -22600 19682 -21224
rect 19648 -24110 19682 -22734
rect 19648 -25620 19682 -24244
rect 21306 -9010 21340 -7634
rect 21306 -10520 21340 -9144
rect 21306 -12030 21340 -10654
rect 21306 -13540 21340 -12164
rect 21306 -15050 21340 -13674
rect 21306 -16560 21340 -15184
rect 21306 -18070 21340 -16694
rect 21306 -19580 21340 -18204
rect 21306 -21090 21340 -19714
rect 21306 -22600 21340 -21224
rect 21306 -24110 21340 -22734
rect 21306 -25620 21340 -24244
rect 21419 -25710 21420 -7544
rect 21420 -25710 21454 -7544
rect 21419 -25764 21454 -25710
rect 4246 -25773 7834 -25771
rect 4246 -25807 4351 -25773
rect 4351 -25807 7737 -25773
rect 7737 -25807 7834 -25773
rect 4246 -25808 7834 -25807
rect 17874 -25772 21459 -25764
rect 17874 -25806 17972 -25772
rect 17972 -25806 21358 -25772
rect 21358 -25806 21459 -25772
rect 4246 -25814 7833 -25808
rect 17874 -25809 21459 -25806
<< metal1 >>
rect -19220 56190 -17382 56450
rect -19220 55462 -18978 56190
rect -17592 55462 -17382 56190
rect -19220 55220 -17382 55462
rect -15220 56190 -13382 56450
rect -15220 55462 -14978 56190
rect -13592 55462 -13382 56190
rect -15220 55220 -13382 55462
rect -11220 56190 -9382 56450
rect -11220 55462 -10978 56190
rect -9592 55462 -9382 56190
rect -11220 55220 -9382 55462
rect -7220 56190 -5382 56450
rect -7220 55462 -6978 56190
rect -5592 55462 -5382 56190
rect -7220 55220 -5382 55462
rect -3220 56190 -1382 56450
rect -3220 55462 -2978 56190
rect -1592 55462 -1382 56190
rect -3220 55220 -1382 55462
rect 780 56190 2618 56450
rect 780 55462 1022 56190
rect 2408 55462 2618 56190
rect 780 55220 2618 55462
rect 4780 56190 6618 56450
rect 4780 55462 5022 56190
rect 6408 55462 6618 56190
rect 4780 55220 6618 55462
rect 8780 56190 10618 56450
rect 8780 55462 9022 56190
rect 10408 55462 10618 56190
rect 8780 55220 10618 55462
rect 12780 56190 14618 56450
rect 12780 55462 13022 56190
rect 14408 55462 14618 56190
rect 12780 55220 14618 55462
rect 16780 56190 18618 56450
rect 16780 55462 17022 56190
rect 18408 55462 18618 56190
rect 16780 55220 18618 55462
rect 20780 56190 22618 56450
rect 20780 55462 21022 56190
rect 22408 55462 22618 56190
rect 20780 55220 22618 55462
rect 24780 56190 26618 56450
rect 24780 55462 25022 56190
rect 26408 55462 26618 56190
rect 24780 55220 26618 55462
rect 28780 56190 30618 56450
rect 28780 55462 29022 56190
rect 30408 55462 30618 56190
rect 28780 55220 30618 55462
rect 32780 56190 34618 56450
rect 32780 55462 33022 56190
rect 34408 55462 34618 56190
rect 32780 55220 34618 55462
rect 36780 56190 38618 56450
rect 36780 55462 37022 56190
rect 38408 55462 38618 56190
rect 36780 55220 38618 55462
rect -20956 54026 -19118 54286
rect -20956 53298 -20714 54026
rect -19328 53298 -19118 54026
rect -20956 53056 -19118 53298
rect 36822 52988 38660 53256
rect 36822 52260 37064 52988
rect 38450 52260 38660 52988
rect 36822 52018 38660 52260
rect -20956 50026 -19118 50286
rect -20956 49298 -20714 50026
rect -19328 49298 -19118 50026
rect -20956 49056 -19118 49298
rect -16276 49684 -15208 49696
rect -16276 49248 -16260 49684
rect -16184 49248 -15940 49684
rect -15864 49248 -15624 49684
rect -15548 49248 -15304 49684
rect -15228 49248 -15208 49684
rect -16276 49230 -15208 49248
rect 36822 48988 38660 49256
rect 36822 48260 37064 48988
rect 38450 48260 38660 48988
rect 36822 48018 38660 48260
rect -20956 46026 -19118 46286
rect -20956 45298 -20714 46026
rect -19328 45298 -19118 46026
rect -20956 45056 -19118 45298
rect 36822 44988 38660 45256
rect -16278 44522 -15210 44530
rect -16278 44090 -16256 44522
rect -16184 44090 -15940 44522
rect -15868 44090 -15620 44522
rect -15548 44090 -15304 44522
rect -15232 44090 -15210 44522
rect -16278 44064 -15210 44090
rect 36822 44260 37064 44988
rect 38450 44260 38660 44988
rect 36822 44018 38660 44260
rect -16220 42400 -16114 42416
rect -20956 42026 -19118 42286
rect -20956 41298 -20714 42026
rect -19328 41298 -19118 42026
rect -16220 41968 -16204 42400
rect -16132 41968 -16114 42400
rect -15872 42384 -15762 42700
rect -15872 42324 -15852 42384
rect -16220 41958 -16114 41968
rect -15868 41952 -15852 42324
rect -15780 41952 -15762 42384
rect -15550 42386 -15440 42720
rect -15550 42344 -15530 42386
rect -15868 41944 -15762 41952
rect -15546 41954 -15530 42344
rect -15458 41954 -15440 42386
rect -15546 41944 -15440 41954
rect -15152 42372 -15046 42382
rect -15152 41940 -15134 42372
rect -15062 41940 -15046 42372
rect -15152 41924 -15046 41940
rect -20956 41056 -19118 41298
rect 36822 40988 38660 41256
rect 36822 40260 37064 40988
rect 38450 40260 38660 40988
rect 36822 40018 38660 40260
rect -20956 38026 -19118 38286
rect -20956 37298 -20714 38026
rect -19328 37298 -19118 38026
rect -20956 37056 -19118 37298
rect -16220 37244 -16114 37256
rect -16220 36812 -16206 37244
rect -16132 36812 -16114 37244
rect -15862 37234 -15776 37238
rect -15862 37226 -15766 37234
rect -15862 37204 -15850 37226
rect -16220 36798 -16114 36812
rect -15860 36794 -15850 37204
rect -15778 36794 -15766 37226
rect -15860 36480 -15766 36794
rect -15550 37222 -15444 37238
rect -15550 36790 -15532 37222
rect -15460 36790 -15444 37222
rect -15550 36552 -15444 36790
rect -15150 37204 -15044 37218
rect -15150 36772 -15134 37204
rect -15060 36772 -15044 37204
rect -15150 36760 -15044 36772
rect 36822 36988 38660 37256
rect -11616 36624 -11334 36712
rect -11616 36552 -11578 36624
rect -15550 36508 -11578 36552
rect -15550 36502 -14890 36508
rect -15550 36498 -15444 36502
rect -16500 36472 -15766 36480
rect -17568 36420 -15766 36472
rect -14860 36458 -14818 36460
rect -14860 36428 -13648 36458
rect -14860 36426 -14378 36428
rect -17566 36060 -17486 36420
rect -16500 36418 -15778 36420
rect -20956 34026 -19118 34286
rect -17564 34082 -17486 36060
rect -17404 36002 -16494 36008
rect -15886 36002 -15794 36006
rect -17404 35958 -15794 36002
rect -17404 35940 -16292 35958
rect -16060 35940 -15794 35958
rect -17404 35938 -16494 35940
rect -17404 35922 -16768 35938
rect -15886 35922 -15794 35940
rect -20956 33298 -20714 34026
rect -19328 33298 -19118 34026
rect -20956 33056 -19118 33298
rect -17568 33956 -17486 34082
rect -17568 31438 -17494 33956
rect -17568 31398 -17490 31438
rect -20956 30026 -19118 30286
rect -20956 29298 -20714 30026
rect -19328 29298 -19118 30026
rect -20956 29056 -19118 29298
rect -17564 28858 -17490 31398
rect -17564 28754 -17484 28858
rect -17558 26286 -17484 28754
rect -20956 26026 -19118 26286
rect -20956 25298 -20714 26026
rect -19328 25298 -19118 26026
rect -20956 25056 -19118 25298
rect -17564 26174 -17484 26286
rect -17564 23602 -17490 26174
rect -17400 23738 -17294 35922
rect -16234 35908 -16122 35916
rect -16234 35476 -16214 35908
rect -16140 35476 -16122 35908
rect -16234 35456 -16122 35476
rect -15886 35490 -15876 35922
rect -15804 35490 -15794 35922
rect -15886 35474 -15794 35490
rect -15568 35994 -15472 35996
rect -14860 35994 -14818 36426
rect -13926 36338 -13648 36428
rect -13926 36162 -13876 36338
rect -13688 36162 -13648 36338
rect -11616 36390 -11578 36508
rect -11378 36390 -11334 36624
rect -11616 36310 -11334 36390
rect -13926 36072 -13648 36162
rect 36822 36260 37064 36988
rect 38450 36260 38660 36988
rect 36822 36018 38660 36260
rect -15568 35960 -14782 35994
rect -15568 35954 -15246 35960
rect -15064 35954 -14782 35960
rect -15568 35922 -15472 35954
rect -15568 35490 -15556 35922
rect -15484 35490 -15472 35922
rect -15568 35476 -15472 35490
rect -15214 35918 -15092 35932
rect -15214 35486 -15190 35918
rect -15116 35486 -15092 35918
rect -15214 35466 -15092 35486
rect 11096 34230 11874 34282
rect 11096 34134 11372 34230
rect 11636 34134 11874 34230
rect 11096 34006 11874 34134
rect -16240 30744 -16114 30768
rect -16240 30310 -16212 30744
rect -16142 30310 -16114 30744
rect -15892 30764 -15788 30774
rect -15892 30330 -15876 30764
rect -15802 30330 -15788 30764
rect -15892 30312 -15788 30330
rect -15572 30764 -15468 30778
rect -15572 30330 -15558 30764
rect -15484 30330 -15468 30764
rect -15572 30316 -15468 30330
rect -15208 30764 -15082 30784
rect -15208 30330 -15186 30764
rect -15116 30330 -15082 30764
rect -16240 30282 -16114 30310
rect -15876 30048 -15796 30312
rect -15560 30070 -15480 30316
rect -15208 30302 -15082 30330
rect -16628 29994 -15790 30048
rect -15560 30016 -14720 30070
rect -16244 29160 -15120 29204
rect -16244 29156 -15554 29160
rect -16244 28718 -16192 29156
rect -16120 28718 -15866 29156
rect -15794 28722 -15554 29156
rect -15482 29152 -15120 29160
rect -15482 28722 -15236 29152
rect -15794 28718 -15236 28722
rect -16244 28714 -15236 28718
rect -15164 28714 -15120 29152
rect -16244 28690 -15120 28714
rect 8998 28258 9706 28310
rect 8998 28064 9172 28258
rect 9526 28064 9706 28258
rect 8998 27782 9706 28064
rect 8990 27738 9706 27782
rect 8996 27582 9706 27738
rect -16254 23998 -15040 24032
rect -16254 23992 -15236 23998
rect -17400 23628 -17292 23738
rect -17554 22788 -17494 23602
rect -17558 22584 -17494 22788
rect -20956 22026 -19118 22286
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -61632 21124 -61262 21200
rect -61634 21108 -61262 21124
rect -94616 20556 -94570 20568
rect -94616 20504 -94610 20556
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -96266 13740 -95320 15274
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -96266 4182 -95320 5274
rect -94790 19180 -94610 20504
rect -94576 20504 -94570 20556
rect -92958 20556 -92912 20568
rect -92958 20504 -92952 20556
rect -94576 19180 -92952 20504
rect -92918 20504 -92912 20556
rect -91300 20556 -91254 20568
rect -91300 20504 -91294 20556
rect -92918 19180 -91294 20504
rect -91260 20504 -91254 20556
rect -89642 20556 -89596 20568
rect -89642 20504 -89636 20556
rect -91260 19180 -89636 20504
rect -89602 20504 -89596 20556
rect -87984 20556 -87938 20568
rect -87984 20504 -87978 20556
rect -89602 19180 -87978 20504
rect -87944 20504 -87938 20556
rect -86326 20556 -86280 20568
rect -86326 20504 -86320 20556
rect -87944 19180 -86320 20504
rect -86286 20504 -86280 20556
rect -84668 20556 -84622 20568
rect -84668 20504 -84662 20556
rect -86286 19180 -84662 20504
rect -84628 20504 -84622 20556
rect -83010 20556 -82964 20568
rect -83010 20504 -83004 20556
rect -84628 19180 -83004 20504
rect -82970 20504 -82964 20556
rect -81352 20556 -81306 20568
rect -81352 20504 -81346 20556
rect -82970 19180 -81346 20504
rect -81312 20504 -81306 20556
rect -79694 20556 -79648 20568
rect -79694 20504 -79688 20556
rect -81312 19180 -79688 20504
rect -79654 20504 -79648 20556
rect -78036 20556 -77990 20568
rect -78036 20504 -78030 20556
rect -79654 19180 -78030 20504
rect -77996 20504 -77990 20556
rect -76378 20556 -76332 20568
rect -76378 20504 -76372 20556
rect -77996 19180 -76372 20504
rect -76338 20504 -76332 20556
rect -74720 20556 -74674 20568
rect -74720 20504 -74714 20556
rect -76338 19180 -74714 20504
rect -74680 20504 -74674 20556
rect -73062 20556 -73016 20568
rect -73062 20504 -73056 20556
rect -74680 19180 -73056 20504
rect -73022 20504 -73016 20556
rect -71404 20556 -71358 20568
rect -71404 20504 -71398 20556
rect -73022 19180 -71398 20504
rect -71364 20504 -71358 20556
rect -69746 20556 -69700 20568
rect -69746 20504 -69740 20556
rect -71364 19180 -69740 20504
rect -69706 20504 -69700 20556
rect -68088 20556 -68042 20568
rect -68088 20504 -68082 20556
rect -69706 19180 -68082 20504
rect -68048 20504 -68042 20556
rect -66430 20556 -66384 20568
rect -66430 20504 -66424 20556
rect -68048 19180 -66424 20504
rect -66390 20504 -66384 20556
rect -64772 20556 -64726 20568
rect -64772 20504 -64766 20556
rect -66390 19180 -64766 20504
rect -64732 20504 -64726 20556
rect -63114 20556 -63068 20568
rect -63114 20504 -63108 20556
rect -64732 19180 -63108 20504
rect -63074 20504 -63068 20556
rect -61634 20556 -61266 21108
rect -61634 20504 -61450 20556
rect -63074 19180 -61450 20504
rect -61416 20504 -61266 20556
rect -59798 20556 -59752 20568
rect -59798 20504 -59792 20556
rect -61416 19180 -59792 20504
rect -59758 20504 -59752 20556
rect -58140 20556 -58094 20568
rect -58140 20504 -58134 20556
rect -59758 19180 -58134 20504
rect -58100 20504 -58094 20556
rect -56482 20556 -56436 20568
rect -56482 20504 -56476 20556
rect -58100 19180 -56476 20504
rect -56442 20504 -56436 20556
rect -54824 20556 -54778 20568
rect -54824 20504 -54818 20556
rect -56442 19180 -54818 20504
rect -54784 20504 -54778 20556
rect -53166 20556 -53120 20568
rect -53166 20504 -53160 20556
rect -54784 19180 -53160 20504
rect -53126 20504 -53120 20556
rect -51508 20556 -51462 20568
rect -51508 20504 -51502 20556
rect -53126 19180 -51502 20504
rect -51468 20504 -51462 20556
rect -49850 20556 -49804 20568
rect -49850 20504 -49844 20556
rect -51468 19180 -49844 20504
rect -49810 20504 -49804 20556
rect -48192 20556 -48146 20568
rect -48192 20504 -48186 20556
rect -49810 19180 -48186 20504
rect -48152 20504 -48146 20556
rect -46534 20556 -46488 20568
rect -46534 20504 -46528 20556
rect -48152 19180 -46528 20504
rect -46494 20504 -46488 20556
rect -44876 20556 -44830 20568
rect -44876 20504 -44870 20556
rect -46494 19180 -44870 20504
rect -44836 20504 -44830 20556
rect -43218 20556 -43172 20568
rect -43218 20504 -43212 20556
rect -44836 19180 -43212 20504
rect -43178 20504 -43172 20556
rect -41560 20556 -41514 20568
rect -41560 20504 -41554 20556
rect -43178 19180 -41554 20504
rect -41520 20504 -41514 20556
rect -39902 20556 -39856 20568
rect -39902 20504 -39896 20556
rect -41520 19180 -39896 20504
rect -39862 20504 -39856 20556
rect -38244 20556 -38198 20568
rect -38244 20504 -38238 20556
rect -39862 19180 -38238 20504
rect -38204 20504 -38198 20556
rect -36586 20556 -36540 20568
rect -36586 20504 -36580 20556
rect -38204 19180 -36580 20504
rect -36546 20504 -36540 20556
rect -34928 20556 -34882 20568
rect -34928 20504 -34922 20556
rect -36546 19180 -34922 20504
rect -34888 20504 -34882 20556
rect -33270 20556 -33224 20568
rect -33270 20504 -33264 20556
rect -34888 19180 -33264 20504
rect -33230 20504 -33224 20556
rect -31612 20556 -31566 20568
rect -31612 20504 -31606 20556
rect -33230 19180 -31606 20504
rect -31572 20504 -31566 20556
rect -29954 20556 -29908 20568
rect -29954 20504 -29948 20556
rect -31572 19180 -29948 20504
rect -29914 20504 -29908 20556
rect -28296 20556 -28250 20568
rect -28296 20504 -28290 20556
rect -29914 19180 -28290 20504
rect -28256 20504 -28250 20556
rect -28256 19180 -28180 20504
rect -94790 18920 -28180 19180
rect -94790 17544 -94610 18920
rect -94576 17544 -92952 18920
rect -92918 17544 -91294 18920
rect -91260 17544 -89636 18920
rect -89602 17544 -87978 18920
rect -87944 17544 -86320 18920
rect -86286 17544 -84662 18920
rect -84628 17544 -83004 18920
rect -82970 17544 -81346 18920
rect -81312 17544 -79688 18920
rect -79654 17544 -78030 18920
rect -77996 17544 -76372 18920
rect -76338 17544 -74714 18920
rect -74680 17544 -73056 18920
rect -73022 17544 -71398 18920
rect -71364 17544 -69740 18920
rect -69706 17544 -68082 18920
rect -68048 17544 -66424 18920
rect -66390 17544 -64766 18920
rect -64732 17544 -63108 18920
rect -63074 17544 -61450 18920
rect -61416 17544 -59792 18920
rect -59758 17544 -58134 18920
rect -58100 17544 -56476 18920
rect -56442 17544 -54818 18920
rect -54784 17544 -53160 18920
rect -53126 17544 -51502 18920
rect -51468 17544 -49844 18920
rect -49810 17544 -48186 18920
rect -48152 17544 -46528 18920
rect -46494 17544 -44870 18920
rect -44836 17544 -43212 18920
rect -43178 17544 -41554 18920
rect -41520 17544 -39896 18920
rect -39862 17544 -38238 18920
rect -38204 17544 -36580 18920
rect -36546 17544 -34922 18920
rect -34888 17544 -33264 18920
rect -33230 17544 -31606 18920
rect -31572 17544 -29948 18920
rect -29914 17544 -28290 18920
rect -28256 17544 -28180 18920
rect -94790 17174 -28180 17544
rect -94790 15798 -94608 17174
rect -94574 15798 -92950 17174
rect -92916 15798 -91292 17174
rect -91258 15798 -89634 17174
rect -89600 15798 -87976 17174
rect -87942 15798 -86318 17174
rect -86284 15798 -84660 17174
rect -84626 15798 -83002 17174
rect -82968 15798 -81344 17174
rect -81310 15798 -79686 17174
rect -79652 15798 -78028 17174
rect -77994 15798 -76370 17174
rect -76336 15798 -74712 17174
rect -74678 15798 -73054 17174
rect -73020 15798 -71396 17174
rect -71362 15798 -69738 17174
rect -69704 15798 -68080 17174
rect -68046 15798 -66422 17174
rect -66388 15798 -64764 17174
rect -64730 15798 -63106 17174
rect -63072 15798 -61448 17174
rect -61414 15798 -59790 17174
rect -59756 15798 -58132 17174
rect -58098 15798 -56474 17174
rect -56440 15798 -54816 17174
rect -54782 15798 -53158 17174
rect -53124 15798 -51500 17174
rect -51466 15798 -49842 17174
rect -49808 15798 -48184 17174
rect -48150 15798 -46526 17174
rect -46492 15798 -44868 17174
rect -44834 15798 -43210 17174
rect -43176 15798 -41552 17174
rect -41518 15798 -39894 17174
rect -39860 15798 -38236 17174
rect -38202 15798 -36578 17174
rect -36544 15798 -34920 17174
rect -34886 15798 -33262 17174
rect -33228 15798 -31604 17174
rect -31570 15798 -29946 17174
rect -29912 15798 -28288 17174
rect -28254 15798 -28180 17174
rect -94790 15538 -28180 15798
rect -94790 14162 -94608 15538
rect -94574 14162 -92950 15538
rect -92916 14162 -91292 15538
rect -91258 14162 -89634 15538
rect -89600 14162 -87976 15538
rect -87942 14162 -86318 15538
rect -86284 14162 -84660 15538
rect -84626 14162 -83002 15538
rect -82968 14162 -81344 15538
rect -81310 14162 -79686 15538
rect -79652 14162 -78028 15538
rect -77994 14162 -76370 15538
rect -76336 14162 -74712 15538
rect -74678 14162 -73054 15538
rect -73020 14162 -71396 15538
rect -71362 14162 -69738 15538
rect -69704 14162 -68080 15538
rect -68046 14162 -66422 15538
rect -66388 14162 -64764 15538
rect -64730 14162 -63106 15538
rect -63072 14162 -61448 15538
rect -61414 14162 -59790 15538
rect -59756 14162 -58132 15538
rect -58098 14162 -56474 15538
rect -56440 14162 -54816 15538
rect -54782 14162 -53158 15538
rect -53124 14162 -51500 15538
rect -51466 14162 -49842 15538
rect -49808 14162 -48184 15538
rect -48150 14162 -46526 15538
rect -46492 14162 -44868 15538
rect -44834 14162 -43210 15538
rect -43176 14162 -41552 15538
rect -41518 14162 -39894 15538
rect -39860 14162 -38236 15538
rect -38202 14162 -36578 15538
rect -36544 14162 -34920 15538
rect -34886 14162 -33262 15538
rect -33228 14162 -31604 15538
rect -31570 14162 -29946 15538
rect -29912 14162 -28288 15538
rect -28254 14162 -28180 15538
rect -94790 13902 -28180 14162
rect -94790 12526 -94608 13902
rect -94574 12526 -92950 13902
rect -92916 12526 -91292 13902
rect -91258 12526 -89634 13902
rect -89600 12526 -87976 13902
rect -87942 12526 -86318 13902
rect -86284 12526 -84660 13902
rect -84626 12526 -83002 13902
rect -82968 12526 -81344 13902
rect -81310 12526 -79686 13902
rect -79652 12526 -78028 13902
rect -77994 12526 -76370 13902
rect -76336 12526 -74712 13902
rect -74678 12526 -73054 13902
rect -73020 12526 -71396 13902
rect -71362 12526 -69738 13902
rect -69704 12526 -68080 13902
rect -68046 12526 -66422 13902
rect -66388 12526 -64764 13902
rect -64730 12526 -63106 13902
rect -63072 12526 -61448 13902
rect -61414 12526 -59790 13902
rect -59756 12526 -58132 13902
rect -58098 12526 -56474 13902
rect -56440 12526 -54816 13902
rect -54782 12526 -53158 13902
rect -53124 12526 -51500 13902
rect -51466 12526 -49842 13902
rect -49808 12526 -48184 13902
rect -48150 12526 -46526 13902
rect -46492 12526 -44868 13902
rect -44834 12526 -43210 13902
rect -43176 12526 -41552 13902
rect -41518 12526 -39894 13902
rect -39860 12526 -38236 13902
rect -38202 12526 -36578 13902
rect -36544 12526 -34920 13902
rect -34886 12526 -33262 13902
rect -33228 12526 -31604 13902
rect -31570 12526 -29946 13902
rect -29912 12526 -28288 13902
rect -28254 12526 -28180 13902
rect -94790 12266 -28180 12526
rect -94790 10890 -94608 12266
rect -94574 10890 -92950 12266
rect -92916 10890 -91292 12266
rect -91258 10890 -89634 12266
rect -89600 10890 -87976 12266
rect -87942 10890 -86318 12266
rect -86284 10890 -84660 12266
rect -84626 10890 -83002 12266
rect -82968 10890 -81344 12266
rect -81310 10890 -79686 12266
rect -79652 10890 -78028 12266
rect -77994 10890 -76370 12266
rect -76336 10890 -74712 12266
rect -74678 10890 -73054 12266
rect -73020 10890 -71396 12266
rect -71362 10890 -69738 12266
rect -69704 10890 -68080 12266
rect -68046 10890 -66422 12266
rect -66388 10890 -64764 12266
rect -64730 10890 -63106 12266
rect -63072 10890 -61448 12266
rect -61414 10890 -59790 12266
rect -59756 10890 -58132 12266
rect -58098 10890 -56474 12266
rect -56440 10890 -54816 12266
rect -54782 10890 -53158 12266
rect -53124 10890 -51500 12266
rect -51466 10890 -49842 12266
rect -49808 10890 -48184 12266
rect -48150 10890 -46526 12266
rect -46492 10890 -44868 12266
rect -44834 10890 -43210 12266
rect -43176 10890 -41552 12266
rect -41518 10890 -39894 12266
rect -39860 10890 -38236 12266
rect -38202 10890 -36578 12266
rect -36544 10890 -34920 12266
rect -34886 10890 -33262 12266
rect -33228 10890 -31604 12266
rect -31570 10890 -29946 12266
rect -29912 10890 -28288 12266
rect -28254 10890 -28180 12266
rect -94790 10628 -28180 10890
rect -94790 9252 -94608 10628
rect -94574 9252 -92950 10628
rect -92916 9252 -91292 10628
rect -91258 9252 -89634 10628
rect -89600 9252 -87976 10628
rect -87942 9252 -86318 10628
rect -86284 9252 -84660 10628
rect -84626 9252 -83002 10628
rect -82968 9252 -81344 10628
rect -81310 9252 -79686 10628
rect -79652 9252 -78028 10628
rect -77994 9252 -76370 10628
rect -76336 9252 -74712 10628
rect -74678 9252 -73054 10628
rect -73020 9252 -71396 10628
rect -71362 9252 -69738 10628
rect -69704 9252 -68080 10628
rect -68046 9252 -66422 10628
rect -66388 9252 -64764 10628
rect -64730 9252 -63106 10628
rect -63072 9252 -61448 10628
rect -61414 9252 -59790 10628
rect -59756 9252 -58132 10628
rect -58098 9252 -56474 10628
rect -56440 9252 -54816 10628
rect -54782 9252 -53158 10628
rect -53124 9252 -51500 10628
rect -51466 9252 -49842 10628
rect -49808 9252 -48184 10628
rect -48150 9252 -46526 10628
rect -46492 9252 -44868 10628
rect -44834 9252 -43210 10628
rect -43176 9252 -41552 10628
rect -41518 9252 -39894 10628
rect -39860 9252 -38236 10628
rect -38202 9252 -36578 10628
rect -36544 9252 -34920 10628
rect -34886 9252 -33262 10628
rect -33228 9252 -31604 10628
rect -31570 9252 -29946 10628
rect -29912 9252 -28288 10628
rect -28254 9252 -28180 10628
rect -94790 8992 -28180 9252
rect -94790 7616 -94608 8992
rect -94574 7616 -92950 8992
rect -92916 7616 -91292 8992
rect -91258 7616 -89634 8992
rect -89600 7616 -87976 8992
rect -87942 7616 -86318 8992
rect -86284 7616 -84660 8992
rect -84626 7616 -83002 8992
rect -82968 7616 -81344 8992
rect -81310 7616 -79686 8992
rect -79652 7616 -78028 8992
rect -77994 7616 -76370 8992
rect -76336 7616 -74712 8992
rect -74678 7616 -73054 8992
rect -73020 7616 -71396 8992
rect -71362 7616 -69738 8992
rect -69704 7616 -68080 8992
rect -68046 7616 -66422 8992
rect -66388 7616 -64764 8992
rect -64730 7616 -63106 8992
rect -63072 7616 -61448 8992
rect -61414 7616 -59790 8992
rect -59756 7616 -58132 8992
rect -58098 7616 -56474 8992
rect -56440 7616 -54816 8992
rect -54782 7616 -53158 8992
rect -53124 7616 -51500 8992
rect -51466 7616 -49842 8992
rect -49808 7616 -48184 8992
rect -48150 7616 -46526 8992
rect -46492 7616 -44868 8992
rect -44834 7616 -43210 8992
rect -43176 7616 -41552 8992
rect -41518 7616 -39894 8992
rect -39860 7616 -38236 8992
rect -38202 7616 -36578 8992
rect -36544 7616 -34920 8992
rect -34886 7616 -33262 8992
rect -33228 7616 -31604 8992
rect -31570 7616 -29946 8992
rect -29912 7616 -28288 8992
rect -28254 7616 -28180 8992
rect -94790 7356 -28180 7616
rect -94790 5980 -94608 7356
rect -94574 5980 -92950 7356
rect -92916 5980 -91292 7356
rect -91258 5980 -89634 7356
rect -89600 5980 -87976 7356
rect -87942 5980 -86318 7356
rect -86284 5980 -84660 7356
rect -84626 5980 -83002 7356
rect -82968 5980 -81344 7356
rect -81310 5980 -79686 7356
rect -79652 5980 -78028 7356
rect -77994 5980 -76370 7356
rect -76336 5980 -74712 7356
rect -74678 5980 -73054 7356
rect -73020 5980 -71396 7356
rect -71362 5980 -69738 7356
rect -69704 5980 -68080 7356
rect -68046 5980 -66422 7356
rect -66388 5980 -64764 7356
rect -64730 5980 -63106 7356
rect -63072 5980 -61448 7356
rect -61414 5980 -59790 7356
rect -59756 5980 -58132 7356
rect -58098 5980 -56474 7356
rect -56440 5980 -54816 7356
rect -54782 5980 -53158 7356
rect -53124 5980 -51500 7356
rect -51466 5980 -49842 7356
rect -49808 5980 -48184 7356
rect -48150 5980 -46526 7356
rect -46492 5980 -44868 7356
rect -44834 5980 -43210 7356
rect -43176 5980 -41552 7356
rect -41518 5980 -39894 7356
rect -39860 5980 -38236 7356
rect -38202 5980 -36578 7356
rect -36544 5980 -34920 7356
rect -34886 5980 -33262 7356
rect -33228 5980 -31604 7356
rect -31570 5980 -29946 7356
rect -29912 5980 -28288 7356
rect -28254 5980 -28180 7356
rect -94790 5720 -28180 5980
rect -94790 4428 -94608 5720
rect -94614 4344 -94608 4428
rect -94574 4428 -92950 5720
rect -94574 4344 -94568 4428
rect -94614 4332 -94568 4344
rect -92956 4344 -92950 4428
rect -92916 4428 -91292 5720
rect -92916 4344 -92910 4428
rect -92956 4332 -92910 4344
rect -91298 4344 -91292 4428
rect -91258 4428 -89634 5720
rect -91258 4344 -91252 4428
rect -91298 4332 -91252 4344
rect -89640 4344 -89634 4428
rect -89600 4428 -87976 5720
rect -89600 4344 -89594 4428
rect -89640 4332 -89594 4344
rect -87982 4344 -87976 4428
rect -87942 4428 -86318 5720
rect -87942 4344 -87936 4428
rect -87982 4332 -87936 4344
rect -86324 4344 -86318 4428
rect -86284 4428 -84660 5720
rect -86284 4344 -86278 4428
rect -86324 4332 -86278 4344
rect -84666 4344 -84660 4428
rect -84626 4428 -83002 5720
rect -84626 4344 -84620 4428
rect -84666 4332 -84620 4344
rect -83008 4344 -83002 4428
rect -82968 4428 -81344 5720
rect -82968 4344 -82962 4428
rect -83008 4332 -82962 4344
rect -81350 4344 -81344 4428
rect -81310 4428 -79686 5720
rect -81310 4344 -81304 4428
rect -81350 4332 -81304 4344
rect -79692 4344 -79686 4428
rect -79652 4428 -78028 5720
rect -79652 4344 -79646 4428
rect -79692 4332 -79646 4344
rect -78034 4344 -78028 4428
rect -77994 4428 -76370 5720
rect -77994 4344 -77988 4428
rect -78034 4332 -77988 4344
rect -76376 4344 -76370 4428
rect -76336 4428 -74712 5720
rect -76336 4344 -76330 4428
rect -76376 4332 -76330 4344
rect -74718 4344 -74712 4428
rect -74678 4428 -73054 5720
rect -74678 4344 -74672 4428
rect -74718 4332 -74672 4344
rect -73060 4344 -73054 4428
rect -73020 4428 -71396 5720
rect -73020 4344 -73014 4428
rect -73060 4332 -73014 4344
rect -71402 4344 -71396 4428
rect -71362 4428 -69738 5720
rect -71362 4344 -71356 4428
rect -71402 4332 -71356 4344
rect -69744 4344 -69738 4428
rect -69704 4428 -68080 5720
rect -69704 4344 -69698 4428
rect -69744 4332 -69698 4344
rect -68086 4344 -68080 4428
rect -68046 4428 -66422 5720
rect -68046 4344 -68040 4428
rect -68086 4332 -68040 4344
rect -66428 4344 -66422 4428
rect -66388 4428 -64764 5720
rect -66388 4344 -66382 4428
rect -66428 4332 -66382 4344
rect -64770 4344 -64764 4428
rect -64730 4428 -63106 5720
rect -64730 4344 -64724 4428
rect -64770 4332 -64724 4344
rect -63112 4344 -63106 4428
rect -63072 4428 -61448 5720
rect -63072 4344 -63066 4428
rect -63112 4332 -63066 4344
rect -61454 4344 -61448 4428
rect -61414 4428 -59790 5720
rect -61414 4344 -61408 4428
rect -61454 4332 -61408 4344
rect -59796 4344 -59790 4428
rect -59756 4428 -58132 5720
rect -59756 4344 -59750 4428
rect -59796 4332 -59750 4344
rect -58138 4344 -58132 4428
rect -58098 4428 -56474 5720
rect -58098 4344 -58092 4428
rect -58138 4332 -58092 4344
rect -56480 4344 -56474 4428
rect -56440 4428 -54816 5720
rect -56440 4344 -56434 4428
rect -56480 4332 -56434 4344
rect -54822 4344 -54816 4428
rect -54782 4428 -53158 5720
rect -54782 4344 -54776 4428
rect -54822 4332 -54776 4344
rect -53164 4344 -53158 4428
rect -53124 4428 -51500 5720
rect -53124 4344 -53118 4428
rect -53164 4332 -53118 4344
rect -51506 4344 -51500 4428
rect -51466 4428 -49842 5720
rect -51466 4344 -51460 4428
rect -51506 4332 -51460 4344
rect -49848 4344 -49842 4428
rect -49808 4428 -48184 5720
rect -49808 4344 -49802 4428
rect -49848 4332 -49802 4344
rect -48190 4344 -48184 4428
rect -48150 4428 -46526 5720
rect -48150 4344 -48144 4428
rect -48190 4332 -48144 4344
rect -46532 4344 -46526 4428
rect -46492 4428 -44868 5720
rect -46492 4344 -46486 4428
rect -46532 4332 -46486 4344
rect -44874 4344 -44868 4428
rect -44834 4428 -43210 5720
rect -44834 4344 -44828 4428
rect -44874 4332 -44828 4344
rect -43216 4344 -43210 4428
rect -43176 4428 -41552 5720
rect -43176 4344 -43170 4428
rect -43216 4332 -43170 4344
rect -41558 4344 -41552 4428
rect -41518 4428 -39894 5720
rect -41518 4344 -41512 4428
rect -41558 4332 -41512 4344
rect -39900 4344 -39894 4428
rect -39860 4428 -38236 5720
rect -39860 4344 -39854 4428
rect -39900 4332 -39854 4344
rect -38242 4344 -38236 4428
rect -38202 4428 -36578 5720
rect -38202 4344 -38196 4428
rect -38242 4332 -38196 4344
rect -36584 4344 -36578 4428
rect -36544 4428 -34920 5720
rect -36544 4344 -36538 4428
rect -36584 4332 -36538 4344
rect -34926 4344 -34920 4428
rect -34886 4428 -33262 5720
rect -34886 4344 -34880 4428
rect -34926 4332 -34880 4344
rect -33268 4344 -33262 4428
rect -33228 4428 -31604 5720
rect -33228 4344 -33222 4428
rect -33268 4332 -33222 4344
rect -31610 4344 -31604 4428
rect -31570 4428 -29946 5720
rect -31570 4344 -31564 4428
rect -31610 4332 -31564 4344
rect -29952 4344 -29946 4428
rect -29912 4428 -28288 5720
rect -29912 4344 -29906 4428
rect -29952 4332 -29906 4344
rect -28294 4344 -28288 4428
rect -28254 4428 -28180 5720
rect -27834 19740 -26806 21200
rect -20956 21298 -20714 22026
rect -19328 21298 -19118 22026
rect -20956 21056 -19118 21298
rect -17558 21090 -17498 22584
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -17562 20904 -17498 21090
rect -17562 19638 -17502 20904
rect -27834 17740 -26806 19274
rect -17568 19206 -17502 19638
rect -17568 18650 -17508 19206
rect -17386 19040 -17292 23628
rect -16254 23554 -16192 23992
rect -16120 23554 -15876 23992
rect -15804 23554 -15552 23992
rect -15480 23590 -15236 23992
rect -15164 23590 -15040 23998
rect -15480 23578 -15220 23590
rect -15182 23578 -15040 23590
rect -15480 23554 -15040 23578
rect -16254 23508 -15040 23554
rect -17400 18852 -17292 19040
rect 8996 21060 9684 27582
rect 11098 22844 11870 34006
rect 36822 32988 38660 33256
rect 36822 32260 37064 32988
rect 38450 32260 38660 32988
rect 36822 32018 38660 32260
rect 36822 28988 38660 29256
rect 36822 28260 37064 28988
rect 38450 28260 38660 28988
rect 36822 28018 38660 28260
rect 36822 24988 38660 25256
rect 36822 24260 37064 24988
rect 38450 24260 38660 24988
rect 36822 24018 38660 24260
rect 8996 20792 9218 21060
rect 9482 20792 9684 21060
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -27834 15740 -26806 17274
rect -20956 18026 -19118 18286
rect -20956 17298 -20714 18026
rect -19328 17298 -19118 18026
rect -20956 17056 -19118 17298
rect -17576 16146 -17504 18650
rect -17400 16740 -17306 18852
rect 8996 17144 9684 20792
rect 11364 20802 11870 22844
rect 36822 20988 38660 21256
rect 16440 20860 16836 20964
rect 16440 20802 16524 20860
rect 11364 20760 16524 20802
rect 11364 17144 11870 20760
rect 16440 20618 16524 20760
rect 16754 20618 16836 20860
rect 16440 20528 16836 20618
rect 36822 20260 37064 20988
rect 38450 20260 38660 20988
rect 36822 20018 38660 20260
rect 13066 18404 13490 18476
rect 13066 18134 13138 18404
rect 13424 18134 13490 18404
rect 13066 18052 13490 18134
rect -17408 16736 -14516 16740
rect 6010 16736 8902 16740
rect 11592 16736 11636 17144
rect -17408 16732 -9876 16736
rect 3218 16732 11638 16736
rect -17408 16728 -7340 16732
rect -2300 16728 11638 16732
rect -17408 16686 11638 16728
rect -17400 16684 -17306 16686
rect -15332 16682 6110 16686
rect 8746 16682 11638 16686
rect -14144 16680 -13470 16682
rect -10232 16678 3282 16682
rect -7826 16674 -2186 16678
rect 13196 16146 13358 18052
rect -17576 15954 13358 16146
rect 36822 16988 38660 17256
rect 36822 16260 37064 16988
rect 38450 16260 38660 16988
rect 36822 16018 38660 16260
rect -17576 15946 13342 15954
rect -17576 15944 -14106 15946
rect -13566 15944 13342 15946
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -27834 13740 -26806 15274
rect -18294 14908 -16456 15184
rect -18294 14180 -18052 14908
rect -16666 14180 -16456 14908
rect -18294 13938 -16456 14180
rect -14294 15084 -14106 15180
rect -13566 15084 -12456 15180
rect -14294 14908 -12456 15084
rect -14294 14180 -14052 14908
rect -12666 14180 -12456 14908
rect -14294 13938 -12456 14180
rect -10294 14908 -8456 15180
rect -10294 14180 -10052 14908
rect -8666 14180 -8456 14908
rect -10294 13938 -8456 14180
rect -6294 14908 -4456 15180
rect -6294 14180 -6052 14908
rect -4666 14180 -4456 14908
rect -6294 13938 -4456 14180
rect -2294 14908 -456 15180
rect -2294 14180 -2052 14908
rect -666 14180 -456 14908
rect -2294 13938 -456 14180
rect 1706 14908 3544 15180
rect 1706 14180 1948 14908
rect 3334 14180 3544 14908
rect 1706 13938 3544 14180
rect 5706 14908 7544 15180
rect 5706 14180 5948 14908
rect 7334 14180 7544 14908
rect 5706 13938 7544 14180
rect 9706 14908 11544 15180
rect 9706 14180 9948 14908
rect 11334 14180 11544 14908
rect 9706 13938 11544 14180
rect 13706 14908 15544 15180
rect 13706 14180 13948 14908
rect 15334 14180 15544 14908
rect 13706 13938 15544 14180
rect 17706 14908 19544 15180
rect 17706 14180 17948 14908
rect 19334 14180 19544 14908
rect 17706 13938 19544 14180
rect 21706 14908 23544 15180
rect 21706 14180 21948 14908
rect 23334 14180 23544 14908
rect 21706 13938 23544 14180
rect 25706 14908 27544 15180
rect 25706 14180 25948 14908
rect 27334 14180 27544 14908
rect 25706 13938 27544 14180
rect 29706 14908 31544 15180
rect 29706 14180 29948 14908
rect 31334 14180 31544 14908
rect 29706 13938 31544 14180
rect 33706 14908 35544 15180
rect 33706 14180 33948 14908
rect 35334 14180 35544 14908
rect 33706 13938 35544 14180
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -27834 11740 -26806 13274
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect 17792 12068 19104 12262
rect 17792 11574 18000 12068
rect 18960 11574 19104 12068
rect 17792 11354 19104 11574
rect -27834 9740 -26806 11274
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect -27834 7740 -26806 9274
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -27834 5740 -26806 7274
rect 0 10884 15826 10916
rect 18118 10884 18178 11354
rect 0 10786 20630 10884
rect 0 10748 142 10786
rect 539 10748 4423 10786
rect 4820 10748 5372 10786
rect 5769 10748 9653 10786
rect 10050 10748 10602 10786
rect 10999 10748 14883 10786
rect 15280 10748 15832 10786
rect 16229 10748 20113 10786
rect 20510 10748 20630 10786
rect 0 10466 20630 10748
rect 0 10428 142 10466
rect 539 10428 4423 10466
rect 4820 10428 5372 10466
rect 5769 10428 9653 10466
rect 10050 10428 10602 10466
rect 10999 10428 14883 10466
rect 15280 10428 15832 10466
rect 16229 10428 20113 10466
rect 20510 10428 20630 10466
rect 0 10300 20630 10428
rect 0 10146 5004 10300
rect 0 10108 142 10146
rect 539 10108 4423 10146
rect 4820 10108 5004 10146
rect 0 9826 5004 10108
rect 0 9788 142 9826
rect 539 9788 4423 9826
rect 4820 9788 5004 9826
rect 0 9506 5004 9788
rect 5354 10140 5804 10154
rect 5354 10070 5368 10140
rect 5800 10070 5804 10140
rect 5354 9822 5804 10070
rect 9644 10140 10098 10158
rect 9644 10070 9650 10140
rect 10082 10070 10098 10140
rect 9644 10052 10098 10070
rect 10552 10144 11002 10154
rect 10552 10070 10564 10144
rect 10998 10070 11002 10144
rect 5354 9752 5368 9822
rect 5800 9752 5804 9822
rect 5354 9742 5804 9752
rect 9642 9822 10098 9836
rect 9642 9752 9650 9822
rect 10082 9752 10098 9822
rect 0 9468 142 9506
rect 539 9468 4423 9506
rect 4820 9468 5004 9506
rect 0 9186 5004 9468
rect 5356 9504 5810 9524
rect 5356 9434 5368 9504
rect 5800 9434 5810 9504
rect 5356 9418 5810 9434
rect 9642 9504 10098 9752
rect 10552 9824 11002 10070
rect 10552 9750 10564 9824
rect 10998 9750 11002 9824
rect 10552 9738 11002 9750
rect 14834 10142 15292 10154
rect 14834 10072 14846 10142
rect 15274 10072 15292 10142
rect 14834 9822 15292 10072
rect 14834 9752 14848 9822
rect 15276 9752 15292 9822
rect 9642 9434 9650 9504
rect 10082 9434 10098 9504
rect 9642 9420 10098 9434
rect 10552 9510 11006 9520
rect 10552 9436 10562 9510
rect 10996 9436 11006 9510
rect 10552 9426 11006 9436
rect 14834 9506 15292 9752
rect 14834 9436 14848 9506
rect 15276 9436 15292 9506
rect 14834 9416 15292 9436
rect 15626 10146 20630 10300
rect 15626 10108 15832 10146
rect 16229 10108 20113 10146
rect 20510 10108 20630 10146
rect 15626 9826 20630 10108
rect 15626 9788 15832 9826
rect 16229 9788 20113 9826
rect 20510 9788 20630 9826
rect 15626 9506 20630 9788
rect 15626 9468 15832 9506
rect 16229 9468 20113 9506
rect 20510 9468 20630 9506
rect 0 9148 142 9186
rect 539 9148 4423 9186
rect 4820 9148 5004 9186
rect 0 8866 5004 9148
rect 0 8828 142 8866
rect 539 8828 4423 8866
rect 4820 8828 5004 8866
rect 0 8546 5004 8828
rect 5362 9186 5806 9194
rect 5362 9112 5368 9186
rect 5802 9112 5806 9186
rect 5362 8870 5806 9112
rect 5362 8796 5366 8870
rect 5800 8796 5806 8870
rect 5362 8786 5806 8796
rect 9636 9188 10092 9206
rect 9636 9116 9650 9188
rect 10082 9116 10092 9188
rect 9636 8870 10092 9116
rect 9636 8798 9650 8870
rect 10082 8798 10092 8870
rect 0 8508 142 8546
rect 539 8508 4423 8546
rect 4820 8508 5004 8546
rect 0 8226 5004 8508
rect 5360 8550 5808 8560
rect 5360 8480 5368 8550
rect 5800 8480 5808 8550
rect 5360 8468 5808 8480
rect 9636 8552 10092 8798
rect 10554 9188 11000 9200
rect 10554 9118 10564 9188
rect 10996 9118 11000 9188
rect 10554 8870 11000 9118
rect 14842 9188 15290 9198
rect 14842 9118 14846 9188
rect 15278 9118 15290 9188
rect 14842 9108 15290 9118
rect 15626 9186 20630 9468
rect 15626 9148 15832 9186
rect 16229 9148 20113 9186
rect 20510 9148 20630 9186
rect 10554 8800 10564 8870
rect 10996 8800 11000 8870
rect 10554 8788 11000 8800
rect 14842 8870 15288 8882
rect 14842 8800 14846 8870
rect 15278 8800 15288 8870
rect 9636 8478 9650 8552
rect 10082 8478 10092 8552
rect 9636 8466 10092 8478
rect 10554 8552 11002 8562
rect 10554 8482 10564 8552
rect 10996 8482 11002 8552
rect 10554 8472 11002 8482
rect 14842 8552 15288 8800
rect 14842 8482 14846 8552
rect 15278 8482 15288 8552
rect 14842 8470 15288 8482
rect 15626 8866 20630 9148
rect 15626 8828 15832 8866
rect 16229 8828 20113 8866
rect 20510 8828 20630 8866
rect 15626 8546 20630 8828
rect 15626 8508 15832 8546
rect 16229 8508 20113 8546
rect 20510 8508 20630 8546
rect 0 8188 142 8226
rect 539 8188 4423 8226
rect 4820 8188 5004 8226
rect 0 7906 5004 8188
rect 0 7868 142 7906
rect 539 7868 4423 7906
rect 4820 7868 5004 7906
rect 0 7586 5004 7868
rect 5354 8236 5804 8244
rect 5354 8234 5806 8236
rect 5354 8162 5368 8234
rect 5794 8162 5806 8234
rect 5354 7916 5806 8162
rect 5354 7844 5368 7916
rect 5794 7844 5806 7916
rect 5354 7842 5806 7844
rect 9646 8232 10092 8250
rect 9646 8160 9650 8232
rect 10082 8160 10092 8232
rect 9646 7916 10092 8160
rect 10556 8236 11010 8246
rect 10556 8162 10562 8236
rect 11000 8162 11010 8236
rect 10556 8152 11010 8162
rect 14836 8234 15290 8246
rect 14836 8164 14846 8234
rect 15278 8164 15290 8234
rect 14836 8152 15290 8164
rect 15626 8226 20630 8508
rect 15626 8188 15832 8226
rect 16229 8188 20113 8226
rect 20510 8188 20630 8226
rect 9646 7844 9650 7916
rect 10082 7844 10092 7916
rect 5354 7832 5804 7842
rect 9646 7832 10092 7844
rect 10552 7918 11006 7934
rect 10552 7848 10562 7918
rect 10998 7848 11006 7918
rect 0 7548 142 7586
rect 539 7548 4423 7586
rect 4820 7548 5004 7586
rect 0 7410 5004 7548
rect 5360 7598 5808 7610
rect 5360 7526 5368 7598
rect 5800 7526 5808 7598
rect 5360 7516 5808 7526
rect 9646 7598 10094 7608
rect 9646 7526 9652 7598
rect 10080 7526 10094 7598
rect 9646 7514 10094 7526
rect 10552 7598 11006 7848
rect 10552 7528 10562 7598
rect 10998 7528 11006 7598
rect 10552 7508 11006 7528
rect 14838 7916 15294 7930
rect 14838 7846 14846 7916
rect 15282 7846 15294 7916
rect 14838 7598 15294 7846
rect 14838 7528 14846 7598
rect 15282 7528 15294 7598
rect 14838 7512 15294 7528
rect 15626 7906 20630 8188
rect 15626 7868 15832 7906
rect 16229 7868 20113 7906
rect 20510 7868 20630 7906
rect 15626 7586 20630 7868
rect 15626 7548 15832 7586
rect 16229 7548 20113 7586
rect 20510 7548 20630 7586
rect 15626 7410 20630 7548
rect 0 7266 20630 7410
rect 0 7228 142 7266
rect 539 7228 4423 7266
rect 4820 7264 15832 7266
rect 4820 7234 10602 7264
rect 4820 7228 5406 7234
rect 0 7196 5406 7228
rect 5803 7196 9687 7234
rect 10084 7226 10602 7234
rect 10999 7226 14883 7264
rect 15280 7228 15832 7264
rect 16229 7228 20113 7266
rect 20510 7228 20630 7266
rect 15280 7226 20630 7228
rect 10084 7196 20630 7226
rect 0 6946 20630 7196
rect 0 6908 142 6946
rect 539 6908 4423 6946
rect 4820 6914 10602 6946
rect 4820 6908 5406 6914
rect 0 6876 5406 6908
rect 5803 6876 9687 6914
rect 10084 6908 10602 6914
rect 10999 6908 14883 6946
rect 15280 6908 15832 6946
rect 16229 6908 20113 6946
rect 20510 6908 20630 6946
rect 10084 6876 20630 6908
rect 0 6808 20630 6876
rect 4578 6778 20630 6808
rect 15626 6776 20630 6778
rect 3910 6604 4078 6634
rect 3910 6526 3932 6604
rect 4052 6526 4078 6604
rect 3910 6492 4078 6526
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 1280 5776 1374 6016
rect 1700 5900 1794 6016
rect 2600 5997 2932 6046
rect 3970 6036 4010 6492
rect 7292 6480 7502 6512
rect 7292 6356 7324 6480
rect 7464 6356 7502 6480
rect 10298 6452 10416 6478
rect 7292 6326 7502 6356
rect 7618 6406 7694 6426
rect 6168 6094 6682 6190
rect 2600 5963 2724 5997
rect 2808 5963 2932 5997
rect 2600 5900 2932 5963
rect 1700 5858 2932 5900
rect 3886 6000 4100 6036
rect 3886 5908 3926 6000
rect 4050 5908 4100 6000
rect 3886 5864 4100 5908
rect 5164 6009 5496 6050
rect 5164 5975 5286 6009
rect 5370 5975 5496 6009
rect 1700 5776 1794 5858
rect 1280 5678 1794 5776
rect -28254 4344 -28248 4428
rect -28294 4332 -28248 4344
rect -61022 4264 -60962 4280
rect -61022 4254 -61008 4264
rect -61196 4230 -61008 4254
rect -60974 4230 -60962 4264
rect -61196 4218 -60962 4230
rect -61196 4192 -61136 4218
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -61198 4050 -61136 4192
rect -61484 4030 -61136 4050
rect -61484 4010 -61134 4030
rect -61482 4006 -61134 4010
rect -61482 3978 -61452 4006
rect -61236 3998 -61134 4006
rect -61484 3976 -61452 3978
rect -61924 3930 -61652 3960
rect -61924 3918 -61848 3930
rect -96396 3740 -62544 3910
rect -61924 3884 -61904 3918
rect -61870 3884 -61848 3918
rect -61680 3890 -61652 3930
rect -61484 3890 -61454 3976
rect -61776 3888 -61730 3890
rect -61924 3864 -61848 3884
rect -61816 3878 -61730 3888
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -61902 3308 -61852 3864
rect -61816 3722 -61770 3878
rect -61816 3670 -61788 3722
rect -61816 3502 -61770 3670
rect -61736 3502 -61730 3878
rect -61816 3490 -61730 3502
rect -61680 3878 -61634 3890
rect -61680 3502 -61674 3878
rect -61640 3502 -61634 3878
rect -61680 3490 -61634 3502
rect -61584 3878 -61538 3890
rect -61584 3502 -61578 3878
rect -61544 3502 -61538 3878
rect -61584 3490 -61538 3502
rect -61488 3878 -61442 3890
rect -61488 3502 -61482 3878
rect -61448 3502 -61442 3878
rect -61488 3490 -61442 3502
rect -61392 3878 -61296 3890
rect -61392 3502 -61386 3878
rect -61352 3718 -61296 3878
rect -61318 3666 -61296 3718
rect -61352 3502 -61296 3666
rect -61392 3492 -61296 3502
rect -61392 3490 -61316 3492
rect -61780 3366 -61744 3490
rect -61584 3368 -61548 3490
rect -61780 3336 -61614 3366
rect -61584 3340 -61390 3368
rect -61584 3338 -61498 3340
rect -61584 3336 -61538 3338
rect -61902 3280 -61710 3308
rect -96396 2966 -62544 3274
rect -61738 3246 -61710 3280
rect -61642 3246 -61614 3336
rect -61426 3246 -61390 3340
rect -61824 3242 -61778 3246
rect -61858 3234 -61778 3242
rect -61858 3184 -61818 3234
rect -61858 3088 -61844 3184
rect -61858 3058 -61818 3088
rect -61784 3058 -61778 3234
rect -61858 3050 -61778 3058
rect -61824 3046 -61778 3050
rect -61738 3234 -61682 3246
rect -61738 3058 -61722 3234
rect -61688 3058 -61682 3234
rect -61738 3046 -61682 3058
rect -61642 3234 -61586 3246
rect -61642 3058 -61626 3234
rect -61592 3058 -61586 3234
rect -61642 3050 -61586 3058
rect -61632 3046 -61586 3050
rect -61536 3234 -61490 3246
rect -61536 3058 -61530 3234
rect -61496 3060 -61490 3234
rect -61440 3242 -61390 3246
rect -61440 3234 -61358 3242
rect -61496 3058 -61484 3060
rect -61536 3046 -61484 3058
rect -61440 3058 -61434 3234
rect -61400 3184 -61358 3234
rect -61374 3098 -61358 3184
rect -61400 3058 -61358 3098
rect -61440 3052 -61358 3058
rect -61440 3046 -61394 3052
rect -61524 2974 -61484 3046
rect -61196 2978 -61134 3998
rect -27834 3846 -26806 5274
rect 2600 5660 2932 5858
rect 1192 5240 1780 5242
rect 1192 5206 2256 5240
rect 1192 5202 1780 5206
rect 1192 5040 1246 5202
rect 1730 5200 1780 5202
rect 970 5026 1114 5040
rect 1160 5038 1246 5040
rect 970 4880 1074 5026
rect 970 4816 988 4880
rect 1048 4816 1074 4880
rect 970 4650 1074 4816
rect 1108 4650 1114 5026
rect 970 4638 1114 4650
rect 1156 5026 1246 5038
rect 1302 5138 1670 5172
rect 1302 5036 1334 5138
rect 1620 5136 1670 5138
rect 1630 5040 1670 5136
rect 1156 4650 1162 5026
rect 1196 4650 1246 5026
rect 1156 4640 1246 4650
rect 1300 5024 1346 5036
rect 1300 4648 1306 5024
rect 1340 4648 1346 5024
rect 1156 4638 1210 4640
rect 1058 4532 1102 4638
rect 1300 4636 1346 4648
rect 1384 5024 1456 5036
rect 1384 4862 1394 5024
rect 1428 4862 1456 5024
rect 1384 4798 1386 4862
rect 1450 4798 1456 4862
rect 1384 4648 1394 4798
rect 1428 4648 1456 4798
rect 1384 4636 1456 4648
rect 1484 5022 1574 5040
rect 1630 5034 1692 5040
rect 1740 5036 1780 5200
rect 1836 5036 1912 5038
rect 1740 5034 1792 5036
rect 1616 5032 1692 5034
rect 1484 4974 1534 5022
rect 1568 4974 1574 5022
rect 1484 4904 1492 4974
rect 1570 4904 1574 4974
rect 1484 4646 1534 4904
rect 1568 4646 1574 4904
rect 1608 5022 1692 5032
rect 1608 4870 1622 5022
rect 1616 4802 1622 4870
rect 1306 4536 1334 4636
rect 1484 4634 1574 4646
rect 1608 4764 1622 4802
rect 1656 4764 1692 5022
rect 1608 4698 1616 4764
rect 1688 4698 1692 4764
rect 1608 4646 1622 4698
rect 1656 4646 1692 4698
rect 1608 4636 1692 4646
rect 1746 5024 1792 5034
rect 1746 4648 1752 5024
rect 1786 4648 1792 5024
rect 1746 4636 1792 4648
rect 1834 5024 1912 5036
rect 1834 4978 1840 5024
rect 1874 4978 1912 5024
rect 1834 4912 1836 4978
rect 1908 4912 1912 4978
rect 1834 4648 1840 4912
rect 1874 4648 1912 4912
rect 1834 4636 1912 4648
rect 1058 4504 1246 4532
rect 1306 4508 1462 4536
rect 1218 4400 1246 4504
rect 1426 4404 1462 4508
rect 1520 4534 1558 4634
rect 1608 4632 1684 4636
rect 1520 4506 1678 4534
rect 1426 4402 1510 4404
rect 1642 4402 1678 4506
rect 1746 4532 1780 4636
rect 1746 4504 1906 4532
rect 1308 4400 1354 4402
rect 1092 4390 1138 4400
rect 1054 4388 1138 4390
rect 1054 4324 1098 4388
rect 1054 4266 1068 4324
rect 1054 4212 1098 4266
rect 1132 4212 1138 4388
rect 1054 4202 1138 4212
rect 1092 4200 1138 4202
rect 1180 4390 1354 4400
rect 1180 4388 1314 4390
rect 1180 4212 1186 4388
rect 1220 4214 1314 4388
rect 1348 4214 1354 4390
rect 1220 4212 1354 4214
rect 1180 4202 1354 4212
rect 1396 4400 1572 4402
rect 1614 4400 1748 4402
rect 1866 4400 1906 4504
rect 1396 4390 1574 4400
rect 1396 4214 1402 4390
rect 1436 4214 1532 4390
rect 1566 4214 1574 4390
rect 1396 4206 1574 4214
rect 1614 4390 1794 4400
rect 1614 4214 1620 4390
rect 1654 4388 1794 4390
rect 1654 4214 1754 4388
rect 1614 4212 1754 4214
rect 1788 4212 1794 4388
rect 1396 4204 1572 4206
rect 1396 4202 1442 4204
rect 1508 4202 1572 4204
rect 1614 4204 1794 4212
rect 1614 4202 1660 4204
rect 1180 4200 1340 4202
rect 1508 4200 1548 4202
rect 1748 4200 1794 4204
rect 1836 4388 1914 4400
rect 1836 4212 1842 4388
rect 1876 4322 1914 4388
rect 1902 4264 1914 4322
rect 1876 4212 1914 4264
rect 1836 4206 1914 4212
rect 1836 4200 1882 4206
rect 1420 4172 1472 4174
rect 2220 4172 2256 5206
rect 2600 5172 2620 5660
rect 2654 5172 2878 5660
rect 2912 5172 2932 5660
rect 2600 5048 2932 5172
rect 5164 5672 5496 5975
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 6168 5756 6682 5854
rect 5164 5184 5182 5672
rect 5216 5184 5440 5672
rect 5474 5184 5496 5672
rect 5164 5048 5496 5184
rect 6378 5220 6966 5260
rect 6378 5058 6432 5220
rect 6916 5218 6966 5220
rect 2600 5000 5496 5048
rect 2600 4874 2932 5000
rect 5164 4878 5496 5000
rect 6156 5044 6300 5058
rect 6346 5056 6432 5058
rect 6156 4898 6260 5044
rect 6156 4834 6174 4898
rect 6234 4834 6260 4898
rect 6156 4668 6260 4834
rect 6294 4668 6300 5044
rect 6156 4656 6300 4668
rect 6342 5044 6432 5056
rect 6488 5156 6856 5190
rect 6488 5054 6520 5156
rect 6806 5154 6856 5156
rect 6816 5058 6856 5154
rect 6342 4668 6348 5044
rect 6382 4668 6432 5044
rect 6342 4658 6432 4668
rect 6486 5042 6532 5054
rect 6486 4666 6492 5042
rect 6526 4666 6532 5042
rect 6342 4656 6396 4658
rect 6244 4550 6288 4656
rect 6486 4654 6532 4666
rect 6570 5042 6642 5054
rect 6570 4880 6580 5042
rect 6614 4880 6642 5042
rect 6570 4816 6572 4880
rect 6636 4816 6642 4880
rect 6570 4666 6580 4816
rect 6614 4666 6642 4816
rect 6570 4654 6642 4666
rect 6670 5040 6760 5058
rect 6816 5052 6878 5058
rect 6926 5054 6966 5218
rect 7022 5054 7098 5056
rect 6926 5052 6978 5054
rect 6802 5050 6878 5052
rect 6670 4992 6720 5040
rect 6754 4992 6760 5040
rect 6670 4922 6678 4992
rect 6756 4922 6760 4992
rect 6670 4664 6720 4922
rect 6754 4664 6760 4922
rect 6794 5040 6878 5050
rect 6794 4888 6808 5040
rect 6802 4820 6808 4888
rect 6492 4554 6520 4654
rect 6670 4652 6760 4664
rect 6794 4782 6808 4820
rect 6842 4782 6878 5040
rect 6794 4716 6802 4782
rect 6874 4716 6878 4782
rect 6794 4664 6808 4716
rect 6842 4664 6878 4716
rect 6794 4654 6878 4664
rect 6932 5042 6978 5052
rect 6932 4666 6938 5042
rect 6972 4666 6978 5042
rect 6932 4654 6978 4666
rect 7020 5042 7098 5054
rect 7020 4996 7026 5042
rect 7060 4996 7098 5042
rect 7020 4930 7022 4996
rect 7094 4990 7098 4996
rect 7360 4994 7400 6326
rect 7618 6306 7630 6406
rect 7682 6306 7694 6406
rect 7618 6286 7694 6306
rect 7794 6402 7880 6426
rect 7794 6318 7810 6402
rect 7862 6318 7880 6402
rect 7794 6294 7880 6318
rect 8522 6424 8622 6444
rect 8522 6326 8534 6424
rect 8612 6326 8622 6424
rect 8522 6294 8622 6326
rect 10298 6320 10312 6452
rect 10400 6320 10416 6452
rect 10298 6300 10416 6320
rect 14776 6236 14874 6254
rect 12764 6192 12872 6204
rect 7894 6118 8126 6142
rect 7894 6066 7918 6118
rect 8094 6106 8126 6118
rect 9882 6106 10080 6130
rect 8094 6098 10080 6106
rect 8094 6066 9902 6098
rect 7894 6046 8126 6066
rect 7440 6022 7580 6040
rect 7440 5936 7456 6022
rect 7564 5994 7580 6022
rect 9220 6012 9406 6038
rect 9220 5994 9246 6012
rect 7564 5946 9246 5994
rect 7564 5944 7982 5946
rect 7564 5936 7580 5944
rect 7440 5916 7580 5936
rect 9220 5928 9246 5946
rect 9378 5928 9406 6012
rect 9882 5988 9902 6066
rect 10058 5988 10080 6098
rect 12764 6106 12778 6192
rect 12860 6106 12872 6192
rect 12764 6088 12872 6106
rect 14196 6174 14294 6180
rect 14196 6120 14218 6174
rect 14278 6120 14294 6174
rect 14776 6176 14794 6236
rect 14856 6176 14874 6236
rect 14196 6104 14294 6120
rect 14466 6114 14518 6166
rect 14776 6158 14874 6176
rect 9882 5952 10080 5988
rect 9220 5900 9406 5928
rect 10438 5864 10554 5904
rect 11480 5882 11994 5978
rect 8832 5858 10554 5864
rect 10704 5858 10810 5878
rect 8832 5818 10810 5858
rect 8832 5814 10554 5818
rect 8834 5746 8872 5814
rect 8652 5743 8872 5746
rect 8648 5737 8872 5743
rect 8648 5703 8660 5737
rect 8744 5703 8872 5737
rect 10438 5712 10554 5814
rect 10704 5808 10810 5818
rect 8648 5697 8872 5703
rect 8652 5696 8872 5697
rect 10430 5711 10908 5712
rect 10430 5677 10454 5711
rect 10538 5677 10908 5711
rect 10430 5664 10908 5677
rect 11480 5642 11574 5882
rect 11900 5642 11994 5882
rect 11480 5544 11994 5642
rect 13780 5609 14168 5642
rect 13780 5575 13934 5609
rect 14018 5575 14168 5609
rect 14468 5604 14516 6114
rect 14800 5932 14840 6158
rect 16222 6124 16480 6142
rect 16222 6060 16254 6124
rect 16448 6106 16480 6124
rect 16448 6068 18262 6106
rect 16448 6060 16480 6068
rect 16222 6042 16480 6060
rect 16332 6004 16502 6010
rect 16332 5954 16344 6004
rect 16478 5954 16502 6004
rect 16332 5946 16502 5954
rect 14760 5886 14874 5932
rect 14760 5784 14782 5886
rect 14842 5784 14874 5886
rect 14760 5732 14874 5784
rect 15370 5621 15758 5670
rect 11726 5488 11766 5544
rect 13780 5488 14168 5575
rect 14356 5596 15156 5604
rect 14356 5594 14950 5596
rect 14356 5556 14378 5594
rect 14562 5558 14950 5594
rect 15134 5558 15156 5596
rect 14562 5556 15156 5558
rect 14356 5544 15156 5556
rect 15370 5587 15522 5621
rect 15606 5587 15758 5621
rect 11726 5460 14168 5488
rect 11734 5452 14168 5460
rect 9002 5424 9085 5444
rect 9661 5426 9743 5446
rect 9661 5424 10287 5426
rect 8810 5412 8862 5418
rect 8550 5400 8596 5412
rect 7360 4990 7878 4994
rect 7094 4950 7878 4990
rect 7094 4946 7400 4950
rect 7094 4930 7098 4946
rect 7020 4666 7026 4930
rect 7060 4666 7098 4930
rect 7020 4654 7098 4666
rect 6244 4522 6432 4550
rect 6492 4526 6648 4554
rect 6404 4418 6432 4522
rect 6612 4422 6648 4526
rect 6706 4552 6744 4652
rect 6794 4650 6870 4654
rect 6706 4524 6864 4552
rect 6612 4420 6696 4422
rect 6828 4420 6864 4524
rect 6932 4550 6966 4654
rect 7834 4560 7874 4950
rect 8550 4912 8556 5400
rect 8590 4912 8596 5400
rect 8550 4900 8596 4912
rect 8808 5400 8862 5412
rect 8808 4912 8814 5400
rect 8848 4912 8862 5400
rect 9002 5408 9629 5424
rect 9002 5316 9022 5408
rect 8808 4900 8862 4912
rect 7834 4554 8170 4560
rect 8810 4554 8862 4900
rect 9003 4894 9022 5316
rect 9080 5386 9629 5408
rect 9080 4898 9551 5386
rect 9585 4898 9629 5386
rect 9080 4894 9629 4898
rect 9003 4866 9629 4894
rect 9661 4900 9691 5424
rect 9731 5388 10287 5424
rect 9731 4900 10209 5388
rect 10243 4900 10287 5388
rect 9661 4868 10287 4900
rect 10344 5374 10390 5386
rect 10344 4886 10350 5374
rect 10384 4886 10390 5374
rect 10344 4874 10390 4886
rect 10602 5374 10648 5386
rect 10602 4886 10608 5374
rect 10642 4886 10648 5374
rect 10934 5292 11110 5324
rect 10934 5216 10964 5292
rect 11074 5264 11110 5292
rect 13780 5272 14168 5452
rect 11554 5264 12142 5272
rect 11074 5232 12142 5264
rect 11074 5222 11608 5232
rect 12092 5230 12142 5232
rect 11074 5216 11110 5222
rect 10934 5174 11110 5216
rect 11554 5070 11608 5222
rect 10602 4874 10648 4886
rect 11332 5056 11476 5070
rect 11522 5068 11608 5070
rect 11332 4910 11436 5056
rect 11332 4846 11350 4910
rect 11410 4846 11436 4910
rect 11332 4680 11436 4846
rect 11470 4680 11476 5056
rect 11332 4668 11476 4680
rect 11518 5056 11608 5068
rect 11664 5168 12032 5202
rect 11664 5066 11696 5168
rect 11982 5166 12032 5168
rect 11992 5070 12032 5166
rect 11518 4680 11524 5056
rect 11558 4680 11608 5056
rect 11518 4670 11608 4680
rect 11662 5054 11708 5066
rect 11662 4678 11668 5054
rect 11702 4678 11708 5054
rect 11518 4668 11572 4670
rect 6932 4522 7092 4550
rect 7052 4488 7092 4522
rect 7834 4520 8862 4554
rect 7840 4516 8862 4520
rect 8020 4514 8862 4516
rect 9216 4558 9418 4584
rect 7448 4488 7500 4490
rect 7052 4442 7500 4488
rect 6494 4418 6540 4420
rect 6278 4408 6324 4418
rect 6240 4406 6324 4408
rect 6240 4342 6284 4406
rect 3630 4246 3894 4288
rect 3630 4172 3668 4246
rect 1396 4168 1750 4172
rect 1396 4130 1426 4168
rect 1466 4164 1750 4168
rect 1466 4130 1704 4164
rect 1738 4130 1750 4164
rect 1396 4126 1750 4130
rect 2220 4126 3668 4172
rect 1420 4124 1472 4126
rect 1694 4120 1750 4126
rect 3630 4070 3668 4126
rect 3862 4070 3894 4246
rect 6240 4284 6254 4342
rect 6240 4230 6284 4284
rect 6318 4230 6324 4406
rect 6240 4220 6324 4230
rect 6278 4218 6324 4220
rect 6366 4408 6540 4418
rect 6366 4406 6500 4408
rect 6366 4230 6372 4406
rect 6406 4232 6500 4406
rect 6534 4232 6540 4408
rect 6406 4230 6540 4232
rect 6366 4220 6540 4230
rect 6582 4418 6758 4420
rect 6800 4418 6934 4420
rect 7052 4418 7100 4442
rect 6582 4408 6760 4418
rect 6582 4232 6588 4408
rect 6622 4232 6718 4408
rect 6752 4232 6760 4408
rect 6582 4224 6760 4232
rect 6800 4408 6980 4418
rect 6800 4232 6806 4408
rect 6840 4406 6980 4408
rect 6840 4232 6940 4406
rect 6800 4230 6940 4232
rect 6974 4230 6980 4406
rect 6582 4222 6758 4224
rect 6582 4220 6628 4222
rect 6694 4220 6758 4222
rect 6800 4222 6980 4230
rect 6800 4220 6846 4222
rect 6366 4218 6526 4220
rect 6694 4218 6734 4220
rect 6934 4218 6980 4222
rect 7022 4406 7100 4418
rect 7022 4230 7028 4406
rect 7062 4340 7100 4406
rect 7088 4282 7100 4340
rect 7448 4324 7500 4442
rect 7924 4462 8082 4474
rect 7924 4408 7950 4462
rect 8056 4450 8082 4462
rect 9216 4470 9248 4558
rect 9382 4470 9418 4558
rect 11180 4576 11296 4590
rect 11180 4506 11198 4576
rect 11274 4564 11296 4576
rect 11420 4564 11464 4668
rect 11662 4666 11708 4678
rect 11746 5054 11818 5066
rect 11746 4892 11756 5054
rect 11790 4892 11818 5054
rect 11746 4828 11748 4892
rect 11812 4828 11818 4892
rect 11746 4678 11756 4828
rect 11790 4678 11818 4828
rect 11746 4666 11818 4678
rect 11846 5052 11936 5070
rect 11992 5064 12054 5070
rect 12102 5066 12142 5230
rect 12198 5066 12274 5068
rect 12102 5064 12154 5066
rect 11978 5062 12054 5064
rect 11846 5004 11896 5052
rect 11930 5004 11936 5052
rect 11846 4934 11854 5004
rect 11932 4934 11936 5004
rect 11846 4676 11896 4934
rect 11930 4676 11936 4934
rect 11970 5052 12054 5062
rect 11970 4900 11984 5052
rect 11978 4832 11984 4900
rect 11274 4562 11464 4564
rect 11668 4566 11696 4666
rect 11846 4664 11936 4676
rect 11970 4794 11984 4832
rect 12018 4794 12054 5052
rect 11970 4728 11978 4794
rect 12050 4728 12054 4794
rect 11970 4676 11984 4728
rect 12018 4676 12054 4728
rect 11970 4666 12054 4676
rect 12108 5054 12154 5064
rect 12108 4678 12114 5054
rect 12148 4678 12154 5054
rect 12108 4666 12154 4678
rect 12196 5054 12274 5066
rect 12196 5008 12202 5054
rect 12236 5052 12274 5054
rect 12236 5008 12630 5052
rect 12196 4942 12198 5008
rect 12270 5006 12630 5008
rect 12270 4942 12274 5006
rect 12196 4678 12202 4942
rect 12236 4678 12274 4942
rect 12196 4666 12274 4678
rect 11274 4534 11608 4562
rect 11668 4538 11824 4566
rect 11274 4530 11452 4534
rect 11274 4506 11296 4530
rect 11180 4488 11296 4506
rect 9216 4450 9418 4470
rect 8056 4440 9418 4450
rect 8056 4418 9334 4440
rect 11580 4430 11608 4534
rect 11788 4434 11824 4538
rect 11882 4564 11920 4664
rect 11970 4662 12046 4666
rect 11882 4536 12040 4564
rect 11788 4432 11872 4434
rect 12004 4432 12040 4536
rect 12108 4562 12142 4666
rect 12108 4534 12268 4562
rect 11670 4430 11716 4432
rect 11454 4420 11500 4430
rect 11416 4418 11500 4420
rect 8056 4408 8082 4418
rect 7924 4394 8082 4408
rect 10188 4366 10252 4382
rect 10188 4324 10200 4366
rect 7446 4298 10200 4324
rect 10244 4298 10252 4366
rect 7446 4288 10252 4298
rect 11416 4354 11460 4418
rect 11416 4296 11430 4354
rect 7062 4230 7100 4282
rect 10188 4280 10252 4288
rect 10488 4264 10756 4296
rect 10488 4230 10514 4264
rect 7022 4224 7100 4230
rect 7984 4228 10514 4230
rect 7022 4218 7068 4224
rect 3630 4038 3894 4070
rect 5820 4026 5960 4062
rect 4636 3966 4900 4004
rect 2190 3880 2310 3902
rect -60278 3740 -26756 3846
rect 2190 3812 2210 3880
rect 2286 3866 2310 3880
rect 4636 3866 4682 3966
rect 2286 3820 4682 3866
rect 2286 3812 2310 3820
rect 2190 3786 2310 3812
rect 4636 3790 4682 3820
rect 4876 3790 4900 3966
rect 5820 3958 5854 4026
rect 5916 4014 5960 4026
rect 6432 4014 6472 4218
rect 6606 4190 6658 4192
rect 6582 4186 6936 4190
rect 6582 4148 6612 4186
rect 6652 4182 6936 4186
rect 6652 4148 6890 4182
rect 6924 4148 6936 4182
rect 6582 4144 6936 4148
rect 6606 4142 6658 4144
rect 6880 4138 6936 4144
rect 7970 4180 10514 4228
rect 5916 3994 6476 4014
rect 7970 3994 8024 4180
rect 10488 4142 10514 4180
rect 10716 4142 10756 4264
rect 11416 4242 11460 4296
rect 11494 4242 11500 4418
rect 11416 4232 11500 4242
rect 11454 4230 11500 4232
rect 11542 4420 11716 4430
rect 11542 4418 11676 4420
rect 11542 4242 11548 4418
rect 11582 4244 11676 4418
rect 11710 4244 11716 4420
rect 11582 4242 11716 4244
rect 11542 4232 11716 4242
rect 11758 4430 11934 4432
rect 11976 4430 12110 4432
rect 12228 4430 12268 4534
rect 11758 4420 11936 4430
rect 11758 4244 11764 4420
rect 11798 4244 11894 4420
rect 11928 4244 11936 4420
rect 11758 4236 11936 4244
rect 11976 4420 12156 4430
rect 11976 4244 11982 4420
rect 12016 4418 12156 4420
rect 12016 4244 12116 4418
rect 11976 4242 12116 4244
rect 12150 4242 12156 4418
rect 11758 4234 11934 4236
rect 11758 4232 11804 4234
rect 11870 4232 11934 4234
rect 11976 4234 12156 4242
rect 11976 4232 12022 4234
rect 11542 4230 11702 4232
rect 11870 4230 11910 4232
rect 12110 4230 12156 4234
rect 12198 4418 12276 4430
rect 12198 4242 12204 4418
rect 12238 4352 12276 4418
rect 12264 4294 12276 4352
rect 12238 4242 12276 4294
rect 12198 4236 12276 4242
rect 12198 4230 12244 4236
rect 11782 4202 11834 4204
rect 11758 4198 12112 4202
rect 11758 4160 11788 4198
rect 11828 4194 12112 4198
rect 11828 4160 12066 4194
rect 12100 4160 12112 4194
rect 11758 4156 12112 4160
rect 11782 4154 11834 4156
rect 12056 4150 12112 4156
rect 10488 4106 10756 4142
rect 5916 3958 8024 3994
rect 5820 3956 8024 3958
rect 10490 3976 10748 4002
rect 5820 3934 5960 3956
rect 6384 3952 8010 3956
rect 6432 3950 6472 3952
rect 10490 3844 10514 3976
rect 10720 3844 10748 3976
rect 4636 3754 4900 3790
rect 8487 3765 9634 3831
rect 10490 3830 10748 3844
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect 8487 3664 8505 3765
rect 8605 3664 9634 3765
rect 8487 3599 9634 3664
rect 9728 3820 10748 3830
rect 9728 3599 10648 3820
rect 10712 3768 10888 3786
rect 10712 3716 10738 3768
rect 10862 3716 10888 3768
rect 10712 3698 10888 3716
rect -60278 3224 -26756 3274
rect 8744 3590 9634 3599
rect 8744 3574 9554 3590
rect 8744 3382 9028 3574
rect 9088 3398 9554 3574
rect 9614 3398 9634 3590
rect 9088 3382 9634 3398
rect 8744 3034 9634 3382
rect 8744 3028 9556 3034
rect -61200 2976 -61132 2978
rect -61234 2974 -61132 2976
rect -61524 2928 -61132 2974
rect -61234 2924 -61132 2928
rect -61234 2922 -61194 2924
rect 5572 2920 5628 2924
rect -61896 2878 -61292 2894
rect -61896 2826 -61864 2878
rect -61806 2826 -61464 2878
rect -61406 2826 -61292 2878
rect -61896 2812 -61292 2826
rect 4036 2876 5628 2920
rect 2604 2604 2936 2638
rect 4036 2628 4082 2876
rect 5572 2874 5628 2876
rect 8744 2836 9032 3028
rect 9092 2842 9556 3028
rect 9612 2842 9634 3034
rect 9092 2836 9634 2842
rect 8744 2744 9634 2836
rect 9758 3590 10648 3599
rect 9758 3574 10568 3590
rect 9758 3382 10042 3574
rect 10102 3398 10568 3574
rect 10628 3398 10648 3590
rect 10102 3382 10648 3398
rect 9758 3034 10648 3382
rect 9758 3028 10570 3034
rect 9758 2836 10046 3028
rect 10106 2842 10570 3028
rect 10626 2842 10648 3034
rect 10106 2836 10648 2842
rect 9758 2744 10648 2836
rect 2604 2570 2730 2604
rect 2814 2570 2936 2604
rect 2604 2476 2936 2570
rect 3334 2606 4740 2628
rect 3334 2572 3356 2606
rect 3740 2572 4328 2606
rect 4712 2572 4740 2606
rect 3334 2556 4740 2572
rect 5154 2604 5486 2630
rect 5154 2570 5264 2604
rect 5348 2570 5486 2604
rect 9588 2600 9772 2628
rect 2604 2388 2626 2476
rect 2660 2388 2884 2476
rect 2918 2388 2936 2476
rect 2604 2298 2936 2388
rect 3088 2490 4122 2508
rect 3088 2478 4134 2490
rect 3088 2390 3102 2478
rect 3136 2390 4074 2478
rect 4108 2390 4134 2478
rect 3088 2368 4134 2390
rect 2736 2250 2786 2298
rect 4056 2250 4134 2368
rect 5154 2476 5486 2570
rect 8524 2568 8882 2580
rect 8524 2528 8538 2568
rect 8580 2528 8882 2568
rect 8524 2516 8882 2528
rect 5154 2388 5160 2476
rect 5194 2388 5418 2476
rect 5452 2388 5486 2476
rect 5154 2290 5486 2388
rect 5268 2250 5318 2290
rect 2730 2214 5318 2250
rect 2730 2198 5312 2214
rect 3990 1892 4032 2198
rect 8836 1982 8882 2516
rect 9588 2464 9616 2600
rect 9736 2578 9772 2600
rect 10714 2598 10860 2608
rect 10714 2578 10728 2598
rect 9736 2536 10728 2578
rect 10846 2536 10860 2598
rect 9736 2532 10860 2536
rect 9736 2464 9772 2532
rect 10714 2524 10860 2532
rect 10916 2544 11106 2574
rect 9588 2430 9772 2464
rect 10916 2452 10952 2544
rect 11072 2518 11106 2544
rect 12588 2518 12630 5006
rect 13780 4784 13830 5272
rect 13864 4784 14088 5272
rect 14122 4966 14168 5272
rect 15370 5284 15758 5587
rect 15370 4966 15418 5284
rect 14122 4930 15418 4966
rect 14122 4784 14168 4930
rect 13780 4462 14168 4784
rect 15370 4796 15418 4930
rect 15452 4796 15676 5284
rect 15710 4796 15758 5284
rect 15370 4490 15758 4796
rect 16462 4364 16498 5946
rect 16916 5824 17430 5920
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect 16638 5108 16776 5134
rect 16638 5008 16664 5108
rect 16746 5062 16776 5108
rect 17210 5062 17798 5064
rect 16746 5024 17798 5062
rect 16746 5008 16776 5024
rect 16638 4978 16776 5008
rect 17210 4862 17264 5024
rect 17748 5022 17798 5024
rect 16988 4848 17132 4862
rect 17178 4860 17264 4862
rect 16988 4702 17092 4848
rect 16988 4638 17006 4702
rect 17066 4638 17092 4702
rect 16988 4472 17092 4638
rect 17126 4472 17132 4848
rect 16988 4460 17132 4472
rect 17174 4848 17264 4860
rect 17320 4960 17688 4994
rect 17320 4858 17352 4960
rect 17638 4958 17688 4960
rect 17648 4862 17688 4958
rect 17174 4472 17180 4848
rect 17214 4472 17264 4848
rect 17174 4462 17264 4472
rect 17318 4846 17364 4858
rect 17318 4470 17324 4846
rect 17358 4470 17364 4846
rect 17174 4460 17228 4462
rect 17076 4364 17120 4460
rect 17318 4458 17364 4470
rect 17402 4846 17474 4858
rect 17402 4684 17412 4846
rect 17446 4684 17474 4846
rect 17402 4620 17404 4684
rect 17468 4620 17474 4684
rect 17402 4470 17412 4620
rect 17446 4470 17474 4620
rect 17402 4458 17474 4470
rect 17502 4844 17592 4862
rect 17648 4856 17710 4862
rect 17758 4858 17798 5022
rect 17854 4858 17930 4860
rect 17758 4856 17810 4858
rect 17634 4854 17710 4856
rect 17502 4796 17552 4844
rect 17586 4796 17592 4844
rect 17502 4726 17510 4796
rect 17588 4726 17592 4796
rect 17502 4468 17552 4726
rect 17586 4468 17592 4726
rect 17626 4844 17710 4854
rect 17626 4692 17640 4844
rect 17634 4624 17640 4692
rect 16462 4354 17120 4364
rect 17324 4358 17352 4458
rect 17502 4456 17592 4468
rect 17626 4586 17640 4624
rect 17674 4586 17710 4844
rect 17626 4520 17634 4586
rect 17706 4520 17710 4586
rect 17626 4468 17640 4520
rect 17674 4468 17710 4520
rect 17626 4458 17710 4468
rect 17764 4846 17810 4856
rect 17764 4470 17770 4846
rect 17804 4470 17810 4846
rect 17764 4458 17810 4470
rect 17852 4846 17930 4858
rect 18214 4846 18252 6068
rect 17852 4800 17858 4846
rect 17892 4808 18252 4846
rect 17892 4800 17930 4808
rect 17852 4734 17854 4800
rect 17926 4734 17930 4800
rect 18214 4796 18252 4808
rect 17852 4470 17858 4734
rect 17892 4470 17930 4734
rect 17852 4458 17930 4470
rect 16462 4328 17264 4354
rect 17324 4330 17480 4358
rect 17076 4326 17264 4328
rect 17236 4222 17264 4326
rect 17444 4226 17480 4330
rect 17538 4356 17576 4456
rect 17626 4454 17702 4458
rect 17538 4328 17696 4356
rect 17444 4224 17528 4226
rect 17660 4224 17696 4328
rect 17764 4354 17798 4458
rect 17764 4326 17924 4354
rect 17326 4222 17372 4224
rect 17110 4212 17156 4222
rect 17072 4210 17156 4212
rect 17072 4146 17116 4210
rect 17072 4088 17086 4146
rect 17072 4034 17116 4088
rect 17150 4034 17156 4210
rect 17072 4024 17156 4034
rect 17110 4022 17156 4024
rect 17198 4212 17372 4222
rect 17198 4210 17332 4212
rect 17198 4034 17204 4210
rect 17238 4036 17332 4210
rect 17366 4036 17372 4212
rect 17238 4034 17372 4036
rect 17198 4024 17372 4034
rect 17414 4222 17590 4224
rect 17632 4222 17766 4224
rect 17884 4222 17924 4326
rect 17414 4212 17592 4222
rect 17414 4036 17420 4212
rect 17454 4036 17550 4212
rect 17584 4036 17592 4212
rect 17414 4028 17592 4036
rect 17632 4212 17812 4222
rect 17632 4036 17638 4212
rect 17672 4210 17812 4212
rect 17672 4036 17772 4210
rect 17632 4034 17772 4036
rect 17806 4034 17812 4210
rect 17414 4026 17590 4028
rect 17414 4024 17460 4026
rect 17526 4024 17590 4026
rect 17632 4026 17812 4034
rect 17632 4024 17678 4026
rect 17198 4022 17358 4024
rect 17526 4022 17566 4024
rect 17766 4022 17812 4026
rect 17854 4210 17932 4222
rect 17854 4034 17860 4210
rect 17894 4144 17932 4210
rect 17920 4086 17932 4144
rect 17894 4034 17932 4086
rect 17854 4028 17932 4034
rect 17854 4022 17900 4028
rect 17438 3994 17490 3996
rect 17414 3990 17768 3994
rect 17414 3952 17444 3990
rect 17484 3986 17768 3990
rect 17484 3952 17722 3986
rect 17756 3952 17768 3986
rect 17414 3948 17768 3952
rect 17438 3946 17490 3948
rect 17712 3942 17768 3948
rect 26112 3638 26592 3676
rect 12850 3506 13108 3516
rect 12850 3414 12876 3506
rect 13064 3476 13108 3506
rect 13064 3432 15128 3476
rect 13064 3414 13108 3432
rect 12850 3402 13108 3414
rect 12668 3376 12776 3396
rect 12668 3272 12686 3376
rect 12746 3368 12776 3376
rect 12746 3364 13322 3368
rect 12746 3322 14142 3364
rect 12746 3314 13322 3322
rect 12746 3272 12776 3314
rect 12668 3262 12776 3272
rect 13260 3186 13672 3260
rect 13260 3152 13422 3186
rect 13506 3152 13672 3186
rect 11072 2476 12642 2518
rect 11072 2452 11106 2476
rect 10916 2434 11106 2452
rect 13260 2408 13672 3152
rect 14104 3096 14142 3322
rect 12272 2228 12500 2270
rect 12272 2096 12308 2228
rect 12452 2096 12500 2228
rect 12272 2064 12500 2096
rect 8834 1980 9258 1982
rect 8834 1960 10296 1980
rect 8834 1920 9248 1960
rect 9446 1958 10296 1960
rect 9446 1920 9859 1958
rect 10063 1920 10296 1958
rect 8834 1918 10296 1920
rect 9106 1914 10296 1918
rect 9228 1908 10296 1914
rect 3316 1698 4628 1892
rect 3316 1204 3524 1698
rect 4484 1204 4628 1698
rect 3316 984 4628 1204
rect 10738 1514 12050 1708
rect 10738 1020 10946 1514
rect 11906 1020 12050 1514
rect 10738 800 12050 1020
rect 13260 1020 13318 2408
rect 13352 1020 13576 2408
rect 13610 1020 13672 2408
rect 13934 3070 14142 3096
rect 15086 3074 15128 3432
rect 26112 3246 26138 3638
rect 26538 3246 26592 3638
rect 14938 3070 15128 3074
rect 15850 3136 16262 3226
rect 26112 3216 26592 3246
rect 26206 3204 26522 3216
rect 15850 3102 16020 3136
rect 16104 3102 16262 3136
rect 13934 3052 14590 3070
rect 13934 3018 13972 3052
rect 14056 3018 14230 3052
rect 14314 3018 14488 3052
rect 14572 3018 14590 3052
rect 13934 3002 14590 3018
rect 14938 3052 15592 3070
rect 14938 3018 14972 3052
rect 15056 3018 15230 3052
rect 15314 3018 15488 3052
rect 15572 3018 15592 3052
rect 14938 3002 15592 3018
rect 13934 2120 14112 3002
rect 13934 2096 14592 2120
rect 13934 2062 13972 2096
rect 14056 2062 14230 2096
rect 14314 2062 14488 2096
rect 14572 2062 14592 2096
rect 13934 2052 14592 2062
rect 14938 2116 15116 3002
rect 15850 2358 16262 3102
rect 26974 2876 27220 2908
rect 27586 2884 27832 2916
rect 26974 2806 27008 2876
rect 27178 2848 27218 2876
rect 27078 2832 27134 2844
rect 26874 2796 26932 2806
rect 26874 2478 26876 2796
rect 26928 2478 26932 2796
rect 26874 2472 26932 2478
rect 26962 2794 27022 2806
rect 26962 2482 26974 2794
rect 27008 2690 27022 2794
rect 27008 2482 27020 2690
rect 27078 2520 27082 2832
rect 27078 2508 27134 2520
rect 27168 2834 27224 2848
rect 27168 2520 27178 2834
rect 27212 2520 27224 2834
rect 27586 2814 27620 2884
rect 27790 2856 27830 2884
rect 28164 2880 28410 2912
rect 28738 2888 28984 2920
rect 29316 2888 29562 2920
rect 29894 2888 30140 2920
rect 30476 2892 30722 2924
rect 27690 2840 27746 2852
rect 27168 2506 27224 2520
rect 27486 2804 27544 2814
rect 26886 2468 26920 2472
rect 26962 2470 27020 2482
rect 14938 2096 15592 2116
rect 14938 2062 14972 2096
rect 15056 2062 15230 2096
rect 15314 2062 15488 2096
rect 15572 2062 15592 2096
rect 13934 1166 14112 2052
rect 14938 2048 15592 2062
rect 13934 1140 14594 1166
rect 13934 1106 13972 1140
rect 14056 1106 14230 1140
rect 14314 1106 14488 1140
rect 14572 1106 14594 1140
rect 13934 1098 14594 1106
rect 14938 1162 15116 2048
rect 14938 1140 15592 1162
rect 14938 1106 14972 1140
rect 15056 1106 15230 1140
rect 15314 1106 15488 1140
rect 15572 1106 15592 1140
rect 13934 1072 14112 1098
rect 14938 1094 15592 1106
rect 14938 1050 15116 1094
rect 13260 814 13672 1020
rect 15850 970 15916 2358
rect 15950 970 16174 2358
rect 16208 1610 16262 2358
rect 26678 2264 26796 2280
rect 26678 2190 26690 2264
rect 26780 2190 26796 2264
rect 26678 2176 26796 2190
rect 26874 2202 26936 2208
rect 26874 2060 26936 2068
rect 27062 2196 27124 2208
rect 27062 2072 27078 2196
rect 27112 2166 27124 2196
rect 27178 2182 27214 2506
rect 27486 2486 27488 2804
rect 27540 2486 27544 2804
rect 27486 2480 27544 2486
rect 27574 2802 27634 2814
rect 27574 2490 27586 2802
rect 27620 2698 27634 2802
rect 27620 2490 27632 2698
rect 27690 2528 27694 2840
rect 27690 2516 27746 2528
rect 27780 2842 27836 2856
rect 27780 2528 27790 2842
rect 27824 2528 27836 2842
rect 28164 2810 28198 2880
rect 28368 2852 28408 2880
rect 28268 2836 28324 2848
rect 27780 2514 27836 2528
rect 28064 2800 28122 2810
rect 27498 2476 27532 2480
rect 27574 2478 27632 2490
rect 27486 2210 27548 2216
rect 27178 2166 27220 2182
rect 27112 2128 27220 2166
rect 27112 2072 27124 2128
rect 27180 2114 27220 2128
rect 27062 2060 27124 2072
rect 27486 2068 27548 2076
rect 27674 2204 27736 2216
rect 27674 2080 27690 2204
rect 27724 2174 27736 2204
rect 27790 2186 27826 2514
rect 28064 2482 28066 2800
rect 28118 2482 28122 2800
rect 28064 2476 28122 2482
rect 28152 2798 28212 2810
rect 28152 2486 28164 2798
rect 28198 2694 28212 2798
rect 28198 2486 28210 2694
rect 28268 2524 28272 2836
rect 28268 2512 28324 2524
rect 28358 2838 28414 2852
rect 28358 2524 28368 2838
rect 28402 2524 28414 2838
rect 28738 2818 28772 2888
rect 28942 2860 28982 2888
rect 28842 2844 28898 2856
rect 28358 2510 28414 2524
rect 28638 2808 28696 2818
rect 28076 2472 28110 2476
rect 28152 2474 28210 2486
rect 28064 2206 28126 2214
rect 28266 2212 28300 2216
rect 27790 2174 27838 2186
rect 27724 2136 27838 2174
rect 27724 2080 27736 2136
rect 27798 2118 27838 2136
rect 27674 2068 27736 2080
rect 28064 2058 28126 2072
rect 28252 2200 28314 2212
rect 28252 2076 28268 2200
rect 28302 2170 28314 2200
rect 28368 2184 28404 2510
rect 28638 2490 28640 2808
rect 28692 2490 28696 2808
rect 28638 2484 28696 2490
rect 28726 2806 28786 2818
rect 28726 2494 28738 2806
rect 28772 2702 28786 2806
rect 28772 2494 28784 2702
rect 28842 2532 28846 2844
rect 28842 2520 28898 2532
rect 28932 2846 28988 2860
rect 28932 2532 28942 2846
rect 28976 2532 28988 2846
rect 29316 2818 29350 2888
rect 29520 2860 29560 2888
rect 29420 2844 29476 2856
rect 28932 2518 28988 2532
rect 29216 2808 29274 2818
rect 28650 2480 28684 2484
rect 28726 2482 28784 2494
rect 28832 2220 28876 2224
rect 28638 2214 28700 2220
rect 28368 2170 28416 2184
rect 28302 2132 28416 2170
rect 28302 2076 28314 2132
rect 28376 2116 28416 2132
rect 28252 2064 28314 2076
rect 28638 2072 28700 2080
rect 28826 2208 28888 2220
rect 28826 2084 28842 2208
rect 28876 2178 28888 2208
rect 28942 2190 28978 2518
rect 29216 2490 29218 2808
rect 29270 2490 29274 2808
rect 29216 2484 29274 2490
rect 29304 2806 29364 2818
rect 29304 2494 29316 2806
rect 29350 2702 29364 2806
rect 29350 2494 29362 2702
rect 29420 2532 29424 2844
rect 29420 2520 29476 2532
rect 29510 2846 29566 2860
rect 29510 2532 29520 2846
rect 29554 2532 29566 2846
rect 29894 2818 29928 2888
rect 30098 2860 30138 2888
rect 29998 2844 30054 2856
rect 29510 2518 29566 2532
rect 29794 2808 29852 2818
rect 29228 2480 29262 2484
rect 29304 2482 29362 2494
rect 29412 2220 29458 2224
rect 29216 2214 29278 2220
rect 28942 2178 28988 2190
rect 28876 2140 28988 2178
rect 28876 2084 28888 2140
rect 28946 2132 28988 2140
rect 28948 2122 28988 2132
rect 28826 2072 28888 2084
rect 29216 2072 29278 2080
rect 29404 2208 29466 2220
rect 29404 2084 29420 2208
rect 29454 2178 29466 2208
rect 29520 2178 29556 2518
rect 29794 2490 29796 2808
rect 29848 2490 29852 2808
rect 29794 2484 29852 2490
rect 29882 2806 29942 2818
rect 29882 2494 29894 2806
rect 29928 2702 29942 2806
rect 29928 2494 29940 2702
rect 29998 2532 30002 2844
rect 29998 2520 30054 2532
rect 30088 2846 30144 2860
rect 30088 2532 30098 2846
rect 30132 2532 30144 2846
rect 30476 2822 30510 2892
rect 30680 2864 30720 2892
rect 31052 2888 31298 2920
rect 30580 2848 30636 2860
rect 30088 2518 30144 2532
rect 30376 2812 30434 2822
rect 29806 2480 29840 2484
rect 29882 2482 29940 2494
rect 29994 2220 30026 2224
rect 29454 2140 29556 2178
rect 29794 2214 29856 2220
rect 29454 2138 29552 2140
rect 29454 2084 29466 2138
rect 29404 2072 29466 2084
rect 29794 2072 29856 2080
rect 29982 2208 30044 2220
rect 29982 2084 29998 2208
rect 30032 2178 30044 2208
rect 30098 2178 30134 2518
rect 30376 2494 30378 2812
rect 30430 2494 30434 2812
rect 30376 2488 30434 2494
rect 30464 2810 30524 2822
rect 30464 2498 30476 2810
rect 30510 2706 30524 2810
rect 30510 2498 30522 2706
rect 30580 2536 30584 2848
rect 30580 2524 30636 2536
rect 30670 2850 30726 2864
rect 30670 2536 30680 2850
rect 30714 2536 30726 2850
rect 31052 2818 31086 2888
rect 31256 2860 31296 2888
rect 31622 2884 31868 2916
rect 31156 2844 31212 2856
rect 30670 2522 30726 2536
rect 30952 2808 31010 2818
rect 30388 2484 30422 2488
rect 30464 2486 30522 2498
rect 30574 2224 30612 2228
rect 30032 2140 30134 2178
rect 30376 2218 30438 2224
rect 30032 2084 30044 2140
rect 29982 2072 30044 2084
rect 30376 2076 30438 2084
rect 30564 2212 30626 2224
rect 30564 2088 30580 2212
rect 30614 2182 30626 2212
rect 30680 2194 30716 2522
rect 30952 2490 30954 2808
rect 31006 2490 31010 2808
rect 30952 2484 31010 2490
rect 31040 2806 31100 2818
rect 31040 2494 31052 2806
rect 31086 2702 31100 2806
rect 31086 2494 31098 2702
rect 31156 2532 31160 2844
rect 31156 2520 31212 2532
rect 31246 2846 31302 2860
rect 31246 2532 31256 2846
rect 31290 2532 31302 2846
rect 31622 2814 31656 2884
rect 31826 2856 31866 2884
rect 31726 2840 31782 2852
rect 31246 2518 31302 2532
rect 31522 2804 31580 2814
rect 30964 2480 30998 2484
rect 31040 2482 31098 2494
rect 31150 2220 31188 2224
rect 30952 2214 31014 2220
rect 30680 2182 30722 2194
rect 30614 2144 30722 2182
rect 30614 2088 30626 2144
rect 30688 2136 30722 2144
rect 30564 2076 30626 2088
rect 30952 2072 31014 2080
rect 31140 2208 31202 2220
rect 31140 2084 31156 2208
rect 31190 2178 31202 2208
rect 31256 2194 31292 2518
rect 31522 2486 31524 2804
rect 31576 2486 31580 2804
rect 31522 2480 31580 2486
rect 31610 2802 31670 2814
rect 31610 2490 31622 2802
rect 31656 2698 31670 2802
rect 31656 2490 31668 2698
rect 31726 2528 31730 2840
rect 31726 2516 31782 2528
rect 31816 2842 31872 2856
rect 31816 2528 31826 2842
rect 31860 2528 31872 2842
rect 31816 2514 31872 2528
rect 31534 2476 31568 2480
rect 31610 2478 31668 2490
rect 31522 2210 31584 2216
rect 31256 2178 31296 2194
rect 31190 2140 31296 2178
rect 31190 2084 31202 2140
rect 31262 2136 31296 2140
rect 31140 2072 31202 2084
rect 31306 2074 31396 2090
rect 17370 1832 18682 2026
rect 31306 2012 31320 2074
rect 31382 2012 31396 2074
rect 31522 2068 31584 2076
rect 31710 2204 31772 2216
rect 31710 2080 31726 2204
rect 31760 2174 31772 2204
rect 31826 2194 31862 2514
rect 32364 2206 32976 2274
rect 31826 2174 31870 2194
rect 31760 2136 31870 2174
rect 31760 2080 31772 2136
rect 31710 2068 31772 2080
rect 32364 2064 32424 2206
rect 31306 1998 31396 2012
rect 32252 1974 32424 2064
rect 17370 1610 17578 1832
rect 16208 1338 17578 1610
rect 18538 1338 18682 1832
rect 32364 1746 32424 1974
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 16208 1294 18682 1338
rect 16208 970 16262 1294
rect 17370 1118 18682 1294
rect 15850 814 16262 970
rect 13260 750 16262 814
rect 28354 906 28530 908
rect 28354 904 28672 906
rect 28354 860 28822 904
rect 28354 846 28820 860
rect 13260 236 13672 750
rect 15850 202 16262 750
rect 28268 740 28326 752
rect 28268 428 28270 740
rect 28324 428 28326 740
rect 28354 740 28416 846
rect 28496 844 28820 846
rect 28554 842 28820 844
rect 28554 790 28612 842
rect 28354 728 28368 740
rect 28268 416 28326 428
rect 28356 428 28368 728
rect 28402 728 28416 740
rect 28468 778 28526 790
rect 28402 428 28414 728
rect 28468 466 28470 778
rect 28524 466 28526 778
rect 28554 778 28614 790
rect 28554 724 28568 778
rect 28468 454 28526 466
rect 28556 466 28568 724
rect 28602 466 28614 778
rect 28762 752 28820 842
rect 28268 234 28326 246
rect 28268 -78 28270 234
rect 28324 -78 28326 234
rect 28268 -90 28326 -78
rect 28356 234 28414 428
rect 28356 -78 28368 234
rect 28402 -78 28414 234
rect 28468 272 28526 284
rect 28468 -40 28470 272
rect 28524 -40 28526 272
rect 28468 -52 28526 -40
rect 28556 272 28614 466
rect 28670 738 28728 750
rect 28670 426 28672 738
rect 28726 426 28728 738
rect 28670 414 28728 426
rect 28756 738 28820 752
rect 28756 426 28770 738
rect 28804 714 28820 738
rect 28804 426 28814 714
rect 28556 -40 28568 272
rect 28602 -40 28614 272
rect 28756 292 28814 426
rect 29792 358 29854 370
rect 29792 292 29808 358
rect 28756 252 29808 292
rect 28268 -274 28326 -262
rect 28268 -586 28270 -274
rect 28324 -586 28326 -274
rect 28268 -598 28326 -586
rect 28356 -274 28414 -78
rect 28356 -586 28368 -274
rect 28402 -586 28414 -274
rect 28468 -236 28526 -224
rect 28468 -548 28470 -236
rect 28524 -548 28526 -236
rect 28468 -560 28526 -548
rect 28556 -236 28614 -40
rect 28668 234 28726 246
rect 28668 -78 28670 234
rect 28724 -78 28726 234
rect 28668 -90 28726 -78
rect 28756 234 28814 252
rect 28844 250 28898 252
rect 28756 -78 28768 234
rect 28802 -78 28814 234
rect 28556 -548 28568 -236
rect 28602 -548 28614 -236
rect 28556 -560 28614 -548
rect 28668 -274 28726 -262
rect 28356 -598 28414 -586
rect 28668 -586 28670 -274
rect 28724 -586 28726 -274
rect 28668 -598 28726 -586
rect 28756 -274 28814 -78
rect 28756 -586 28768 -274
rect 28802 -586 28814 -274
rect 29792 -266 29808 252
rect 29842 -266 29854 358
rect 29792 -278 29854 -266
rect 28756 -598 28814 -586
rect 9025 -847 10957 -804
rect 13408 -805 13447 -804
rect 9025 -859 10890 -847
rect 9025 -892 9089 -859
rect 8734 -958 10850 -892
rect 8734 -992 8763 -958
rect 8797 -992 8855 -958
rect 8889 -992 8947 -958
rect 8981 -992 9039 -958
rect 9073 -992 9131 -958
rect 9165 -992 9223 -958
rect 9257 -992 9315 -958
rect 9349 -992 9407 -958
rect 9441 -992 9499 -958
rect 9533 -992 9591 -958
rect 9625 -992 9683 -958
rect 9717 -992 9775 -958
rect 9809 -992 9867 -958
rect 9901 -992 9959 -958
rect 9993 -992 10051 -958
rect 10085 -992 10143 -958
rect 10177 -992 10235 -958
rect 10269 -992 10327 -958
rect 10361 -992 10419 -958
rect 10453 -992 10511 -958
rect 10545 -992 10603 -958
rect 10637 -992 10695 -958
rect 10729 -992 10787 -958
rect 10821 -992 10850 -958
rect 8734 -1023 10850 -992
rect 8925 -1128 8983 -1122
rect 8925 -1162 8937 -1128
rect 8971 -1131 8983 -1128
rect 9025 -1131 9089 -1023
rect 9303 -1128 9361 -1122
rect 9303 -1131 9315 -1128
rect 8971 -1159 9315 -1131
rect 8971 -1162 8983 -1159
rect 8925 -1168 8983 -1162
rect 9025 -1184 9089 -1159
rect 9303 -1162 9315 -1159
rect 9349 -1131 9361 -1128
rect 9927 -1128 9985 -1122
rect 9927 -1131 9939 -1128
rect 9349 -1159 9939 -1131
rect 9349 -1162 9361 -1159
rect 9303 -1168 9361 -1162
rect 9927 -1162 9939 -1159
rect 9973 -1162 9985 -1128
rect 9927 -1168 9985 -1162
rect 9025 -1236 9031 -1184
rect 9083 -1236 9089 -1184
rect 9025 -1239 9089 -1236
rect 10460 -1256 10546 -1234
rect 10919 -1251 10955 -847
rect 11491 -855 13447 -805
rect 11491 -892 11556 -855
rect 11200 -958 13316 -892
rect 11200 -992 11229 -958
rect 11263 -992 11321 -958
rect 11355 -992 11413 -958
rect 11447 -992 11505 -958
rect 11539 -992 11597 -958
rect 11631 -992 11689 -958
rect 11723 -992 11781 -958
rect 11815 -992 11873 -958
rect 11907 -992 11965 -958
rect 11999 -992 12057 -958
rect 12091 -992 12149 -958
rect 12183 -992 12241 -958
rect 12275 -992 12333 -958
rect 12367 -992 12425 -958
rect 12459 -992 12517 -958
rect 12551 -992 12609 -958
rect 12643 -992 12701 -958
rect 12735 -992 12793 -958
rect 12827 -992 12885 -958
rect 12919 -992 12977 -958
rect 13011 -992 13069 -958
rect 13103 -992 13161 -958
rect 13195 -992 13253 -958
rect 13287 -992 13316 -958
rect 11200 -1023 13316 -992
rect 11391 -1128 11449 -1122
rect 11391 -1162 11403 -1128
rect 11437 -1131 11449 -1128
rect 11491 -1131 11556 -1023
rect 11769 -1128 11827 -1122
rect 11769 -1131 11781 -1128
rect 11437 -1159 11781 -1131
rect 11437 -1162 11449 -1159
rect 11391 -1168 11449 -1162
rect 11491 -1183 11556 -1159
rect 11769 -1162 11781 -1159
rect 11815 -1131 11827 -1128
rect 12393 -1128 12451 -1122
rect 12393 -1131 12405 -1128
rect 11815 -1159 12405 -1131
rect 11815 -1162 11827 -1159
rect 11769 -1168 11827 -1162
rect 12393 -1162 12405 -1159
rect 12439 -1162 12451 -1128
rect 12393 -1168 12451 -1162
rect 11491 -1235 11497 -1183
rect 11549 -1235 11556 -1183
rect 11491 -1239 11556 -1235
rect 8844 -1264 8902 -1258
rect 8844 -1298 8856 -1264
rect 8890 -1267 8902 -1264
rect 9211 -1264 9269 -1258
rect 9211 -1267 9223 -1264
rect 8890 -1295 9223 -1267
rect 8890 -1298 8902 -1295
rect 8844 -1304 8902 -1298
rect 9211 -1298 9223 -1295
rect 9257 -1267 9269 -1264
rect 9927 -1264 9985 -1258
rect 9927 -1267 9939 -1264
rect 9257 -1295 9939 -1267
rect 9257 -1298 9269 -1295
rect 9211 -1304 9269 -1298
rect 9927 -1298 9939 -1295
rect 9973 -1298 9985 -1264
rect 9927 -1304 9985 -1298
rect 10143 -1269 10201 -1263
rect 10143 -1303 10155 -1269
rect 10189 -1303 10201 -1269
rect 10143 -1322 10201 -1303
rect 10460 -1308 10478 -1256
rect 10530 -1308 10546 -1256
rect 10143 -1325 10265 -1322
rect 9483 -1332 9613 -1326
rect 9483 -1366 9495 -1332
rect 9529 -1366 9567 -1332
rect 9601 -1335 9613 -1332
rect 10143 -1335 10205 -1325
rect 9601 -1363 10205 -1335
rect 9601 -1366 9613 -1363
rect 9483 -1372 9613 -1366
rect 9841 -1373 10205 -1363
rect 9841 -1471 9894 -1373
rect 10197 -1377 10205 -1373
rect 10257 -1377 10265 -1325
rect 10197 -1471 10265 -1377
rect 10460 -1377 10546 -1308
rect 10769 -1257 10955 -1251
rect 10769 -1309 10775 -1257
rect 10827 -1309 10955 -1257
rect 10769 -1315 10955 -1309
rect 11061 -1254 11282 -1248
rect 13408 -1249 13447 -855
rect 11061 -1286 11220 -1254
rect 11061 -1377 11091 -1286
rect 11140 -1306 11220 -1286
rect 11272 -1306 11282 -1254
rect 13232 -1254 13447 -1249
rect 11310 -1264 11368 -1258
rect 11310 -1298 11322 -1264
rect 11356 -1267 11368 -1264
rect 11677 -1264 11735 -1258
rect 11677 -1267 11689 -1264
rect 11356 -1295 11689 -1267
rect 11356 -1298 11368 -1295
rect 11310 -1304 11368 -1298
rect 11677 -1298 11689 -1295
rect 11723 -1267 11735 -1264
rect 12393 -1264 12451 -1258
rect 12393 -1267 12405 -1264
rect 11723 -1295 12405 -1267
rect 11723 -1298 11735 -1295
rect 11677 -1304 11735 -1298
rect 12393 -1298 12405 -1295
rect 12439 -1298 12451 -1264
rect 12393 -1304 12451 -1298
rect 12609 -1269 12667 -1263
rect 12609 -1303 12621 -1269
rect 12655 -1303 12667 -1269
rect 11140 -1313 11282 -1306
rect 12609 -1323 12667 -1303
rect 13232 -1306 13244 -1254
rect 13296 -1306 13447 -1254
rect 13232 -1313 13447 -1306
rect 11949 -1332 12079 -1326
rect 11949 -1366 11961 -1332
rect 11995 -1366 12033 -1332
rect 12067 -1335 12079 -1332
rect 12609 -1327 12738 -1323
rect 12609 -1335 12674 -1327
rect 12067 -1363 12674 -1335
rect 12067 -1366 12079 -1363
rect 11949 -1372 12079 -1366
rect 10460 -1415 11091 -1377
rect 10870 -1419 11091 -1415
rect 12664 -1379 12674 -1363
rect 12726 -1379 12738 -1327
rect 10870 -1444 10906 -1419
rect 8734 -1502 10850 -1471
rect 8734 -1536 8763 -1502
rect 8797 -1536 8855 -1502
rect 8889 -1536 8947 -1502
rect 8981 -1536 9039 -1502
rect 9073 -1536 9131 -1502
rect 9165 -1536 9223 -1502
rect 9257 -1536 9315 -1502
rect 9349 -1536 9407 -1502
rect 9441 -1536 9499 -1502
rect 9533 -1536 9591 -1502
rect 9625 -1536 9683 -1502
rect 9717 -1536 9775 -1502
rect 9809 -1536 9867 -1502
rect 9901 -1536 9959 -1502
rect 9993 -1536 10051 -1502
rect 10085 -1536 10143 -1502
rect 10177 -1536 10235 -1502
rect 10269 -1536 10327 -1502
rect 10361 -1536 10419 -1502
rect 10453 -1536 10511 -1502
rect 10545 -1536 10603 -1502
rect 10637 -1536 10695 -1502
rect 10729 -1536 10787 -1502
rect 10821 -1536 10850 -1502
rect 8734 -1567 10850 -1536
rect 8733 -1614 10850 -1567
rect 9841 -2099 9894 -1614
rect 10878 -1651 10906 -1444
rect 12664 -1432 12738 -1379
rect 12664 -1471 13663 -1432
rect 11200 -1488 13663 -1471
rect 11200 -1502 13316 -1488
rect 11200 -1536 11229 -1502
rect 11263 -1536 11321 -1502
rect 11355 -1536 11413 -1502
rect 11447 -1536 11505 -1502
rect 11539 -1536 11597 -1502
rect 11631 -1536 11689 -1502
rect 11723 -1536 11781 -1502
rect 11815 -1536 11873 -1502
rect 11907 -1536 11965 -1502
rect 11999 -1536 12057 -1502
rect 12091 -1536 12149 -1502
rect 12183 -1536 12241 -1502
rect 12275 -1536 12333 -1502
rect 12367 -1536 12425 -1502
rect 12459 -1536 12517 -1502
rect 12551 -1536 12609 -1502
rect 12643 -1536 12701 -1502
rect 12735 -1536 12793 -1502
rect 12827 -1536 12885 -1502
rect 12919 -1536 12977 -1502
rect 13011 -1536 13069 -1502
rect 13103 -1536 13161 -1502
rect 13195 -1536 13253 -1502
rect 13287 -1536 13316 -1502
rect 11200 -1567 13316 -1536
rect 11201 -1606 13317 -1567
rect 9842 -2443 9894 -2099
rect 10075 -1680 10906 -1651
rect 10075 -1684 10124 -1680
rect 10456 -1684 10906 -1680
rect 10075 -2050 10103 -1684
rect 11490 -1699 13447 -1670
rect 11490 -1729 11561 -1699
rect 10152 -1760 10428 -1729
rect 10152 -1794 10181 -1760
rect 10215 -1794 10273 -1760
rect 10307 -1794 10365 -1760
rect 10399 -1794 10428 -1760
rect 10152 -1825 10428 -1794
rect 11200 -1760 13316 -1729
rect 11200 -1794 11229 -1760
rect 11263 -1794 11321 -1760
rect 11355 -1794 11413 -1760
rect 11447 -1794 11505 -1760
rect 11539 -1794 11597 -1760
rect 11631 -1794 11689 -1760
rect 11723 -1794 11781 -1760
rect 11815 -1794 11873 -1760
rect 11907 -1794 11965 -1760
rect 11999 -1794 12057 -1760
rect 12091 -1794 12149 -1760
rect 12183 -1794 12241 -1760
rect 12275 -1794 12333 -1760
rect 12367 -1794 12425 -1760
rect 12459 -1794 12517 -1760
rect 12551 -1794 12609 -1760
rect 12643 -1794 12701 -1760
rect 12735 -1794 12793 -1760
rect 12827 -1794 12885 -1760
rect 12919 -1794 12977 -1760
rect 13011 -1794 13069 -1760
rect 13103 -1794 13161 -1760
rect 13195 -1794 13253 -1760
rect 13287 -1794 13316 -1760
rect 11200 -1825 13316 -1794
rect 11391 -1930 11449 -1924
rect 11391 -1964 11403 -1930
rect 11437 -1933 11449 -1930
rect 11490 -1933 11561 -1825
rect 11769 -1930 11827 -1924
rect 11769 -1933 11781 -1930
rect 11437 -1961 11781 -1933
rect 11437 -1964 11449 -1961
rect 11391 -1970 11449 -1964
rect 11490 -2016 11561 -1961
rect 11769 -1964 11781 -1961
rect 11815 -1933 11827 -1930
rect 12393 -1930 12451 -1924
rect 12393 -1933 12405 -1930
rect 11815 -1961 12405 -1933
rect 11815 -1964 11827 -1961
rect 11769 -1970 11827 -1964
rect 12393 -1964 12405 -1961
rect 12439 -1964 12451 -1930
rect 12393 -1970 12451 -1964
rect 10759 -2019 10907 -2018
rect 10759 -2025 11279 -2019
rect 10075 -2066 10221 -2050
rect 10075 -2086 10181 -2066
rect 10215 -2086 10221 -2066
rect 10759 -2077 11221 -2025
rect 11273 -2077 11279 -2025
rect 10759 -2082 11279 -2077
rect 10075 -2138 10166 -2086
rect 10218 -2138 10221 -2086
rect 10075 -2150 10221 -2138
rect 10258 -2083 11279 -2082
rect 11310 -2066 11368 -2060
rect 10258 -2088 10811 -2083
rect 10258 -2140 10264 -2088
rect 10316 -2140 10811 -2088
rect 11310 -2100 11322 -2066
rect 11356 -2069 11368 -2066
rect 11490 -2068 11500 -2016
rect 11552 -2068 11561 -2016
rect 11490 -2069 11561 -2068
rect 11677 -2066 11735 -2060
rect 11677 -2069 11689 -2066
rect 11356 -2097 11689 -2069
rect 11356 -2100 11368 -2097
rect 11310 -2106 11368 -2100
rect 11677 -2100 11689 -2097
rect 11723 -2069 11735 -2066
rect 12393 -2066 12451 -2060
rect 12393 -2069 12405 -2066
rect 11723 -2097 12405 -2069
rect 11723 -2100 11735 -2097
rect 11677 -2106 11735 -2100
rect 12393 -2100 12405 -2097
rect 12439 -2100 12451 -2066
rect 12393 -2106 12451 -2100
rect 12609 -2071 12667 -2065
rect 12609 -2105 12621 -2071
rect 12655 -2105 12667 -2071
rect 13402 -2086 13447 -1699
rect 12609 -2123 12667 -2105
rect 13236 -2090 13447 -2086
rect 12609 -2128 12739 -2123
rect 10258 -2146 10811 -2140
rect 11949 -2134 12079 -2128
rect 11949 -2168 11961 -2134
rect 11995 -2168 12033 -2134
rect 12067 -2137 12079 -2134
rect 12609 -2137 12674 -2128
rect 12067 -2165 12674 -2137
rect 12067 -2168 12079 -2165
rect 11949 -2174 12079 -2168
rect 12664 -2180 12674 -2165
rect 12726 -2180 12739 -2128
rect 13236 -2142 13242 -2090
rect 13294 -2142 13447 -2090
rect 13236 -2146 13447 -2142
rect 13402 -2147 13447 -2146
rect 12664 -2273 12739 -2180
rect 10152 -2304 10428 -2273
rect 10152 -2338 10181 -2304
rect 10215 -2338 10273 -2304
rect 10307 -2338 10365 -2304
rect 10399 -2338 10428 -2304
rect 10152 -2395 10428 -2338
rect 11200 -2304 13316 -2273
rect 11200 -2338 11229 -2304
rect 11263 -2338 11321 -2304
rect 11355 -2338 11413 -2304
rect 11447 -2338 11505 -2304
rect 11539 -2338 11597 -2304
rect 11631 -2338 11689 -2304
rect 11723 -2338 11781 -2304
rect 11815 -2338 11873 -2304
rect 11907 -2338 11965 -2304
rect 11999 -2338 12057 -2304
rect 12091 -2338 12149 -2304
rect 12183 -2338 12241 -2304
rect 12275 -2338 12333 -2304
rect 12367 -2338 12425 -2304
rect 12459 -2338 12517 -2304
rect 12551 -2338 12609 -2304
rect 12643 -2338 12701 -2304
rect 12735 -2338 12793 -2304
rect 12827 -2338 12885 -2304
rect 12919 -2338 12977 -2304
rect 13011 -2338 13069 -2304
rect 13103 -2338 13161 -2304
rect 13195 -2338 13253 -2304
rect 13287 -2338 13316 -2304
rect 11200 -2387 13316 -2338
rect 12664 -2443 12739 -2387
rect 13603 -2443 13663 -1488
rect 9842 -2480 13665 -2443
rect 9842 -2482 12677 -2480
rect 12738 -2481 13665 -2480
rect -9158 -4228 33162 -4197
rect -9158 -4262 -9129 -4228
rect -9095 -4262 -9037 -4228
rect -9003 -4262 -8945 -4228
rect -8911 -4262 -8853 -4228
rect -8819 -4262 -8761 -4228
rect -8727 -4262 -8669 -4228
rect -8635 -4262 -8577 -4228
rect -8543 -4262 -8485 -4228
rect -8451 -4262 -8393 -4228
rect -8359 -4262 -8301 -4228
rect -8267 -4262 -8209 -4228
rect -8175 -4262 -8117 -4228
rect -8083 -4262 -8025 -4228
rect -7991 -4262 -7933 -4228
rect -7899 -4262 -7841 -4228
rect -7807 -4262 -7749 -4228
rect -7715 -4262 -7657 -4228
rect -7623 -4262 -7565 -4228
rect -7531 -4262 -7473 -4228
rect -7439 -4262 -7381 -4228
rect -7347 -4262 -7289 -4228
rect -7255 -4262 -7197 -4228
rect -7163 -4262 -7105 -4228
rect -7071 -4262 -7013 -4228
rect -6979 -4262 -6921 -4228
rect -6887 -4262 -6829 -4228
rect -6795 -4262 -6737 -4228
rect -6703 -4262 -6645 -4228
rect -6611 -4262 -6553 -4228
rect -6519 -4262 -6461 -4228
rect -6427 -4262 -6369 -4228
rect -6335 -4262 -6277 -4228
rect -6243 -4262 -6185 -4228
rect -6151 -4262 -6093 -4228
rect -6059 -4262 -6001 -4228
rect -5967 -4262 -5909 -4228
rect -5875 -4262 -5817 -4228
rect -5783 -4262 -5725 -4228
rect -5691 -4262 -5633 -4228
rect -5599 -4262 -5541 -4228
rect -5507 -4262 -5449 -4228
rect -5415 -4262 -5357 -4228
rect -5323 -4262 -5265 -4228
rect -5231 -4262 -5173 -4228
rect -5139 -4262 -5081 -4228
rect -5047 -4262 -4989 -4228
rect -4955 -4262 -4897 -4228
rect -4863 -4262 -4805 -4228
rect -4771 -4262 -4713 -4228
rect -4679 -4262 -4621 -4228
rect -4587 -4262 -4529 -4228
rect -4495 -4262 -4437 -4228
rect -4403 -4262 -4345 -4228
rect -4311 -4262 -4253 -4228
rect -4219 -4262 -4161 -4228
rect -4127 -4262 -4069 -4228
rect -4035 -4262 -3977 -4228
rect -3943 -4262 -3885 -4228
rect -3851 -4262 -3793 -4228
rect -3759 -4262 -3701 -4228
rect -3667 -4262 -3609 -4228
rect -3575 -4262 -3517 -4228
rect -3483 -4262 -3425 -4228
rect -3391 -4262 -3333 -4228
rect -3299 -4262 -3241 -4228
rect -3207 -4262 -3149 -4228
rect -3115 -4262 -3057 -4228
rect -3023 -4262 -2965 -4228
rect -2931 -4262 -2873 -4228
rect -2839 -4262 -2781 -4228
rect -2747 -4262 -2689 -4228
rect -2655 -4262 -2597 -4228
rect -2563 -4262 -2505 -4228
rect -2471 -4262 -2413 -4228
rect -2379 -4262 -2321 -4228
rect -2287 -4262 -2229 -4228
rect -2195 -4262 -2137 -4228
rect -2103 -4262 -2045 -4228
rect -2011 -4262 -1953 -4228
rect -1919 -4262 -1861 -4228
rect -1827 -4262 -1769 -4228
rect -1735 -4262 -1677 -4228
rect -1643 -4262 -1585 -4228
rect -1551 -4262 -1493 -4228
rect -1459 -4262 -1401 -4228
rect -1367 -4262 -1309 -4228
rect -1275 -4262 -1217 -4228
rect -1183 -4262 -1125 -4228
rect -1091 -4262 -1033 -4228
rect -999 -4262 -941 -4228
rect -907 -4262 -849 -4228
rect -815 -4262 -757 -4228
rect -723 -4262 -665 -4228
rect -631 -4262 -573 -4228
rect -539 -4262 -481 -4228
rect -447 -4262 -389 -4228
rect -355 -4262 -297 -4228
rect -263 -4262 -205 -4228
rect -171 -4262 -113 -4228
rect -79 -4262 -21 -4228
rect 13 -4262 71 -4228
rect 105 -4262 163 -4228
rect 197 -4262 255 -4228
rect 289 -4262 347 -4228
rect 381 -4262 439 -4228
rect 473 -4262 531 -4228
rect 565 -4262 623 -4228
rect 657 -4262 715 -4228
rect 749 -4262 807 -4228
rect 841 -4262 899 -4228
rect 933 -4262 991 -4228
rect 1025 -4262 1083 -4228
rect 1117 -4262 1175 -4228
rect 1209 -4262 1267 -4228
rect 1301 -4262 1359 -4228
rect 1393 -4262 1451 -4228
rect 1485 -4262 1543 -4228
rect 1577 -4262 1635 -4228
rect 1669 -4262 1727 -4228
rect 1761 -4262 1819 -4228
rect 1853 -4262 1911 -4228
rect 1945 -4262 2003 -4228
rect 2037 -4262 2095 -4228
rect 2129 -4262 2187 -4228
rect 2221 -4262 2279 -4228
rect 2313 -4262 2371 -4228
rect 2405 -4262 2463 -4228
rect 2497 -4262 2555 -4228
rect 2589 -4262 2647 -4228
rect 2681 -4262 2739 -4228
rect 2773 -4262 2831 -4228
rect 2865 -4262 2923 -4228
rect 2957 -4262 3015 -4228
rect 3049 -4262 3107 -4228
rect 3141 -4262 3199 -4228
rect 3233 -4262 3291 -4228
rect 3325 -4262 3383 -4228
rect 3417 -4262 3475 -4228
rect 3509 -4262 3567 -4228
rect 3601 -4262 3659 -4228
rect 3693 -4262 3751 -4228
rect 3785 -4262 3843 -4228
rect 3877 -4262 3935 -4228
rect 3969 -4262 4027 -4228
rect 4061 -4262 4119 -4228
rect 4153 -4262 4211 -4228
rect 4245 -4262 4303 -4228
rect 4337 -4262 4395 -4228
rect 4429 -4262 4487 -4228
rect 4521 -4262 4579 -4228
rect 4613 -4262 4671 -4228
rect 4705 -4262 4763 -4228
rect 4797 -4262 4855 -4228
rect 4889 -4262 4947 -4228
rect 4981 -4262 5039 -4228
rect 5073 -4262 5131 -4228
rect 5165 -4262 5223 -4228
rect 5257 -4262 5315 -4228
rect 5349 -4262 5407 -4228
rect 5441 -4262 5499 -4228
rect 5533 -4262 5591 -4228
rect 5625 -4262 5683 -4228
rect 5717 -4262 5775 -4228
rect 5809 -4262 5867 -4228
rect 5901 -4262 5959 -4228
rect 5993 -4262 6051 -4228
rect 6085 -4262 6143 -4228
rect 6177 -4262 6235 -4228
rect 6269 -4262 6327 -4228
rect 6361 -4262 6419 -4228
rect 6453 -4262 6511 -4228
rect 6545 -4262 6603 -4228
rect 6637 -4262 6695 -4228
rect 6729 -4262 6787 -4228
rect 6821 -4262 6879 -4228
rect 6913 -4262 6971 -4228
rect 7005 -4262 7063 -4228
rect 7097 -4262 7155 -4228
rect 7189 -4262 7247 -4228
rect 7281 -4262 7339 -4228
rect 7373 -4262 7431 -4228
rect 7465 -4262 7523 -4228
rect 7557 -4262 7615 -4228
rect 7649 -4262 7707 -4228
rect 7741 -4262 7799 -4228
rect 7833 -4262 7891 -4228
rect 7925 -4262 7983 -4228
rect 8017 -4262 8075 -4228
rect 8109 -4262 8167 -4228
rect 8201 -4262 8259 -4228
rect 8293 -4262 8351 -4228
rect 8385 -4262 8443 -4228
rect 8477 -4262 8535 -4228
rect 8569 -4262 8627 -4228
rect 8661 -4262 8719 -4228
rect 8753 -4262 8811 -4228
rect 8845 -4262 8903 -4228
rect 8937 -4262 8995 -4228
rect 9029 -4262 9087 -4228
rect 9121 -4262 9179 -4228
rect 9213 -4262 9271 -4228
rect 9305 -4262 9363 -4228
rect 9397 -4262 9455 -4228
rect 9489 -4262 9547 -4228
rect 9581 -4262 9639 -4228
rect 9673 -4262 9731 -4228
rect 9765 -4262 9823 -4228
rect 9857 -4262 9915 -4228
rect 9949 -4262 10007 -4228
rect 10041 -4262 10099 -4228
rect 10133 -4262 10191 -4228
rect 10225 -4262 10283 -4228
rect 10317 -4262 10375 -4228
rect 10409 -4262 10467 -4228
rect 10501 -4262 10559 -4228
rect 10593 -4262 10651 -4228
rect 10685 -4262 10743 -4228
rect 10777 -4262 10835 -4228
rect 10869 -4262 10927 -4228
rect 10961 -4262 11019 -4228
rect 11053 -4262 11111 -4228
rect 11145 -4262 11203 -4228
rect 11237 -4262 11295 -4228
rect 11329 -4262 11387 -4228
rect 11421 -4262 11479 -4228
rect 11513 -4262 11571 -4228
rect 11605 -4262 11663 -4228
rect 11697 -4262 11755 -4228
rect 11789 -4262 11847 -4228
rect 11881 -4262 11939 -4228
rect 11973 -4262 12031 -4228
rect 12065 -4262 12123 -4228
rect 12157 -4262 12215 -4228
rect 12249 -4262 12307 -4228
rect 12341 -4262 12399 -4228
rect 12433 -4262 12491 -4228
rect 12525 -4262 12583 -4228
rect 12617 -4262 12675 -4228
rect 12709 -4262 12767 -4228
rect 12801 -4262 12859 -4228
rect 12893 -4262 12951 -4228
rect 12985 -4262 13043 -4228
rect 13077 -4262 13135 -4228
rect 13169 -4262 13227 -4228
rect 13261 -4262 13319 -4228
rect 13353 -4262 13411 -4228
rect 13445 -4262 13503 -4228
rect 13537 -4262 13595 -4228
rect 13629 -4262 13687 -4228
rect 13721 -4262 13779 -4228
rect 13813 -4262 13871 -4228
rect 13905 -4262 13963 -4228
rect 13997 -4262 14055 -4228
rect 14089 -4262 14147 -4228
rect 14181 -4262 14239 -4228
rect 14273 -4262 14331 -4228
rect 14365 -4262 14423 -4228
rect 14457 -4262 14515 -4228
rect 14549 -4262 14607 -4228
rect 14641 -4262 14699 -4228
rect 14733 -4262 14791 -4228
rect 14825 -4262 14883 -4228
rect 14917 -4262 14975 -4228
rect 15009 -4262 15067 -4228
rect 15101 -4262 15159 -4228
rect 15193 -4262 15251 -4228
rect 15285 -4262 15343 -4228
rect 15377 -4262 15435 -4228
rect 15469 -4262 15527 -4228
rect 15561 -4262 15619 -4228
rect 15653 -4262 15711 -4228
rect 15745 -4262 15803 -4228
rect 15837 -4262 15895 -4228
rect 15929 -4262 15987 -4228
rect 16021 -4262 16079 -4228
rect 16113 -4262 16171 -4228
rect 16205 -4262 16263 -4228
rect 16297 -4262 16355 -4228
rect 16389 -4262 16447 -4228
rect 16481 -4262 16539 -4228
rect 16573 -4262 16631 -4228
rect 16665 -4262 16723 -4228
rect 16757 -4262 16815 -4228
rect 16849 -4262 16907 -4228
rect 16941 -4262 16999 -4228
rect 17033 -4262 17091 -4228
rect 17125 -4262 17183 -4228
rect 17217 -4262 17275 -4228
rect 17309 -4262 17367 -4228
rect 17401 -4262 17459 -4228
rect 17493 -4262 17551 -4228
rect 17585 -4262 17643 -4228
rect 17677 -4262 17735 -4228
rect 17769 -4262 17827 -4228
rect 17861 -4262 17919 -4228
rect 17953 -4262 18011 -4228
rect 18045 -4262 18103 -4228
rect 18137 -4262 18195 -4228
rect 18229 -4262 18287 -4228
rect 18321 -4262 18379 -4228
rect 18413 -4262 18471 -4228
rect 18505 -4262 18563 -4228
rect 18597 -4262 18655 -4228
rect 18689 -4262 18747 -4228
rect 18781 -4262 18839 -4228
rect 18873 -4262 18931 -4228
rect 18965 -4262 19023 -4228
rect 19057 -4262 19115 -4228
rect 19149 -4262 19207 -4228
rect 19241 -4262 19299 -4228
rect 19333 -4262 19391 -4228
rect 19425 -4262 19483 -4228
rect 19517 -4262 19575 -4228
rect 19609 -4262 19667 -4228
rect 19701 -4262 19759 -4228
rect 19793 -4262 19851 -4228
rect 19885 -4262 19943 -4228
rect 19977 -4262 20035 -4228
rect 20069 -4262 20127 -4228
rect 20161 -4262 20219 -4228
rect 20253 -4262 20311 -4228
rect 20345 -4262 20403 -4228
rect 20437 -4262 20495 -4228
rect 20529 -4262 20587 -4228
rect 20621 -4262 20679 -4228
rect 20713 -4262 20771 -4228
rect 20805 -4262 20863 -4228
rect 20897 -4262 20955 -4228
rect 20989 -4262 21047 -4228
rect 21081 -4262 21139 -4228
rect 21173 -4262 21231 -4228
rect 21265 -4262 21323 -4228
rect 21357 -4262 21415 -4228
rect 21449 -4262 21507 -4228
rect 21541 -4262 21599 -4228
rect 21633 -4262 21691 -4228
rect 21725 -4262 21783 -4228
rect 21817 -4262 21875 -4228
rect 21909 -4262 21967 -4228
rect 22001 -4262 22059 -4228
rect 22093 -4262 22151 -4228
rect 22185 -4262 22243 -4228
rect 22277 -4262 22335 -4228
rect 22369 -4262 22427 -4228
rect 22461 -4262 22519 -4228
rect 22553 -4262 22611 -4228
rect 22645 -4262 22703 -4228
rect 22737 -4262 22795 -4228
rect 22829 -4262 22887 -4228
rect 22921 -4262 22979 -4228
rect 23013 -4262 23071 -4228
rect 23105 -4262 23163 -4228
rect 23197 -4262 23255 -4228
rect 23289 -4262 23347 -4228
rect 23381 -4262 23439 -4228
rect 23473 -4262 23531 -4228
rect 23565 -4262 23623 -4228
rect 23657 -4262 23715 -4228
rect 23749 -4262 23807 -4228
rect 23841 -4262 23899 -4228
rect 23933 -4262 23991 -4228
rect 24025 -4262 24083 -4228
rect 24117 -4262 24175 -4228
rect 24209 -4262 24267 -4228
rect 24301 -4262 24359 -4228
rect 24393 -4262 24451 -4228
rect 24485 -4262 24543 -4228
rect 24577 -4262 24635 -4228
rect 24669 -4262 24727 -4228
rect 24761 -4262 24819 -4228
rect 24853 -4262 24911 -4228
rect 24945 -4262 25003 -4228
rect 25037 -4262 25095 -4228
rect 25129 -4262 25187 -4228
rect 25221 -4262 25279 -4228
rect 25313 -4262 25371 -4228
rect 25405 -4262 25463 -4228
rect 25497 -4262 25555 -4228
rect 25589 -4262 25647 -4228
rect 25681 -4262 25739 -4228
rect 25773 -4262 25831 -4228
rect 25865 -4262 25923 -4228
rect 25957 -4262 26015 -4228
rect 26049 -4262 26107 -4228
rect 26141 -4262 26199 -4228
rect 26233 -4262 26291 -4228
rect 26325 -4262 26383 -4228
rect 26417 -4262 26475 -4228
rect 26509 -4262 26567 -4228
rect 26601 -4262 26659 -4228
rect 26693 -4262 26751 -4228
rect 26785 -4262 26843 -4228
rect 26877 -4262 26935 -4228
rect 26969 -4262 27027 -4228
rect 27061 -4262 27119 -4228
rect 27153 -4262 27211 -4228
rect 27245 -4262 27303 -4228
rect 27337 -4262 27395 -4228
rect 27429 -4262 27487 -4228
rect 27521 -4262 27579 -4228
rect 27613 -4262 27671 -4228
rect 27705 -4262 27763 -4228
rect 27797 -4262 27855 -4228
rect 27889 -4262 27947 -4228
rect 27981 -4262 28039 -4228
rect 28073 -4262 28131 -4228
rect 28165 -4262 28223 -4228
rect 28257 -4262 28315 -4228
rect 28349 -4262 28407 -4228
rect 28441 -4262 28499 -4228
rect 28533 -4262 28591 -4228
rect 28625 -4262 28683 -4228
rect 28717 -4262 28775 -4228
rect 28809 -4262 28867 -4228
rect 28901 -4262 28959 -4228
rect 28993 -4262 29051 -4228
rect 29085 -4262 29143 -4228
rect 29177 -4262 29235 -4228
rect 29269 -4262 29327 -4228
rect 29361 -4262 29419 -4228
rect 29453 -4262 29511 -4228
rect 29545 -4262 29603 -4228
rect 29637 -4262 29695 -4228
rect 29729 -4262 29787 -4228
rect 29821 -4262 29879 -4228
rect 29913 -4262 29971 -4228
rect 30005 -4262 30063 -4228
rect 30097 -4262 30155 -4228
rect 30189 -4262 30247 -4228
rect 30281 -4262 30339 -4228
rect 30373 -4262 30431 -4228
rect 30465 -4262 30523 -4228
rect 30557 -4262 30615 -4228
rect 30649 -4262 30707 -4228
rect 30741 -4262 30799 -4228
rect 30833 -4262 30891 -4228
rect 30925 -4262 30983 -4228
rect 31017 -4262 31075 -4228
rect 31109 -4262 31167 -4228
rect 31201 -4262 31259 -4228
rect 31293 -4262 31351 -4228
rect 31385 -4262 31443 -4228
rect 31477 -4262 31535 -4228
rect 31569 -4262 31627 -4228
rect 31661 -4262 31719 -4228
rect 31753 -4262 31811 -4228
rect 31845 -4262 31903 -4228
rect 31937 -4262 31995 -4228
rect 32029 -4262 32087 -4228
rect 32121 -4262 32179 -4228
rect 32213 -4262 32271 -4228
rect 32305 -4262 32363 -4228
rect 32397 -4262 32455 -4228
rect 32489 -4262 32547 -4228
rect 32581 -4262 32639 -4228
rect 32673 -4262 32731 -4228
rect 32765 -4262 32823 -4228
rect 32857 -4262 32915 -4228
rect 32949 -4262 33007 -4228
rect 33041 -4262 33099 -4228
rect 33133 -4262 33162 -4228
rect -9158 -4293 33162 -4262
rect -8967 -4398 -8909 -4392
rect -8967 -4432 -8955 -4398
rect -8921 -4401 -8909 -4398
rect -8589 -4398 -8531 -4392
rect -8589 -4401 -8577 -4398
rect -8921 -4429 -8577 -4401
rect -8921 -4432 -8909 -4429
rect -8967 -4438 -8909 -4432
rect -8589 -4432 -8577 -4429
rect -8543 -4401 -8531 -4398
rect -7965 -4398 -7907 -4392
rect -7965 -4401 -7953 -4398
rect -8543 -4429 -7953 -4401
rect -8543 -4432 -8531 -4429
rect -8589 -4438 -8531 -4432
rect -7965 -4432 -7953 -4429
rect -7919 -4432 -7907 -4398
rect -7965 -4438 -7907 -4432
rect -6851 -4398 -6793 -4392
rect -6851 -4432 -6839 -4398
rect -6805 -4401 -6793 -4398
rect -6473 -4398 -6415 -4392
rect -6473 -4401 -6461 -4398
rect -6805 -4429 -6461 -4401
rect -6805 -4432 -6793 -4429
rect -6851 -4438 -6793 -4432
rect -6473 -4432 -6461 -4429
rect -6427 -4401 -6415 -4398
rect -5849 -4398 -5791 -4392
rect -5849 -4401 -5837 -4398
rect -6427 -4429 -5837 -4401
rect -6427 -4432 -6415 -4429
rect -6473 -4438 -6415 -4432
rect -5849 -4432 -5837 -4429
rect -5803 -4432 -5791 -4398
rect -5849 -4438 -5791 -4432
rect -4735 -4398 -4677 -4392
rect -4735 -4432 -4723 -4398
rect -4689 -4401 -4677 -4398
rect -4357 -4398 -4299 -4392
rect -4357 -4401 -4345 -4398
rect -4689 -4429 -4345 -4401
rect -4689 -4432 -4677 -4429
rect -4735 -4438 -4677 -4432
rect -4357 -4432 -4345 -4429
rect -4311 -4401 -4299 -4398
rect -3733 -4398 -3675 -4392
rect -3733 -4401 -3721 -4398
rect -4311 -4429 -3721 -4401
rect -4311 -4432 -4299 -4429
rect -4357 -4438 -4299 -4432
rect -3733 -4432 -3721 -4429
rect -3687 -4432 -3675 -4398
rect -3733 -4438 -3675 -4432
rect -2619 -4398 -2561 -4392
rect -2619 -4432 -2607 -4398
rect -2573 -4401 -2561 -4398
rect -2241 -4398 -2183 -4392
rect -2241 -4401 -2229 -4398
rect -2573 -4429 -2229 -4401
rect -2573 -4432 -2561 -4429
rect -2619 -4438 -2561 -4432
rect -2241 -4432 -2229 -4429
rect -2195 -4401 -2183 -4398
rect -1617 -4398 -1559 -4392
rect -1617 -4401 -1605 -4398
rect -2195 -4429 -1605 -4401
rect -2195 -4432 -2183 -4429
rect -2241 -4438 -2183 -4432
rect -1617 -4432 -1605 -4429
rect -1571 -4432 -1559 -4398
rect -1617 -4438 -1559 -4432
rect -503 -4398 -445 -4392
rect -503 -4432 -491 -4398
rect -457 -4401 -445 -4398
rect -125 -4398 -67 -4392
rect -125 -4401 -113 -4398
rect -457 -4429 -113 -4401
rect -457 -4432 -445 -4429
rect -503 -4438 -445 -4432
rect -125 -4432 -113 -4429
rect -79 -4401 -67 -4398
rect 499 -4398 557 -4392
rect 499 -4401 511 -4398
rect -79 -4429 511 -4401
rect -79 -4432 -67 -4429
rect -125 -4438 -67 -4432
rect 499 -4432 511 -4429
rect 545 -4432 557 -4398
rect 499 -4438 557 -4432
rect 1613 -4398 1671 -4392
rect 1613 -4432 1625 -4398
rect 1659 -4401 1671 -4398
rect 1991 -4398 2049 -4392
rect 1991 -4401 2003 -4398
rect 1659 -4429 2003 -4401
rect 1659 -4432 1671 -4429
rect 1613 -4438 1671 -4432
rect 1991 -4432 2003 -4429
rect 2037 -4401 2049 -4398
rect 2615 -4398 2673 -4392
rect 2615 -4401 2627 -4398
rect 2037 -4429 2627 -4401
rect 2037 -4432 2049 -4429
rect 1991 -4438 2049 -4432
rect 2615 -4432 2627 -4429
rect 2661 -4432 2673 -4398
rect 2615 -4438 2673 -4432
rect 3729 -4398 3787 -4392
rect 3729 -4432 3741 -4398
rect 3775 -4401 3787 -4398
rect 4107 -4398 4165 -4392
rect 4107 -4401 4119 -4398
rect 3775 -4429 4119 -4401
rect 3775 -4432 3787 -4429
rect 3729 -4438 3787 -4432
rect 4107 -4432 4119 -4429
rect 4153 -4401 4165 -4398
rect 4731 -4398 4789 -4392
rect 4731 -4401 4743 -4398
rect 4153 -4429 4743 -4401
rect 4153 -4432 4165 -4429
rect 4107 -4438 4165 -4432
rect 4731 -4432 4743 -4429
rect 4777 -4432 4789 -4398
rect 4731 -4438 4789 -4432
rect 5845 -4398 5903 -4392
rect 5845 -4432 5857 -4398
rect 5891 -4401 5903 -4398
rect 6223 -4398 6281 -4392
rect 6223 -4401 6235 -4398
rect 5891 -4429 6235 -4401
rect 5891 -4432 5903 -4429
rect 5845 -4438 5903 -4432
rect 6223 -4432 6235 -4429
rect 6269 -4401 6281 -4398
rect 6847 -4398 6905 -4392
rect 6847 -4401 6859 -4398
rect 6269 -4429 6859 -4401
rect 6269 -4432 6281 -4429
rect 6223 -4438 6281 -4432
rect 6847 -4432 6859 -4429
rect 6893 -4432 6905 -4398
rect 6847 -4438 6905 -4432
rect 7961 -4398 8019 -4392
rect 7961 -4432 7973 -4398
rect 8007 -4401 8019 -4398
rect 8339 -4398 8397 -4392
rect 8339 -4401 8351 -4398
rect 8007 -4429 8351 -4401
rect 8007 -4432 8019 -4429
rect 7961 -4438 8019 -4432
rect 8339 -4432 8351 -4429
rect 8385 -4401 8397 -4398
rect 8963 -4398 9021 -4392
rect 8963 -4401 8975 -4398
rect 8385 -4429 8975 -4401
rect 8385 -4432 8397 -4429
rect 8339 -4438 8397 -4432
rect 8963 -4432 8975 -4429
rect 9009 -4432 9021 -4398
rect 8963 -4438 9021 -4432
rect 10077 -4398 10135 -4392
rect 10077 -4432 10089 -4398
rect 10123 -4401 10135 -4398
rect 10455 -4398 10513 -4392
rect 10455 -4401 10467 -4398
rect 10123 -4429 10467 -4401
rect 10123 -4432 10135 -4429
rect 10077 -4438 10135 -4432
rect 10455 -4432 10467 -4429
rect 10501 -4401 10513 -4398
rect 11079 -4398 11137 -4392
rect 11079 -4401 11091 -4398
rect 10501 -4429 11091 -4401
rect 10501 -4432 10513 -4429
rect 10455 -4438 10513 -4432
rect 11079 -4432 11091 -4429
rect 11125 -4432 11137 -4398
rect 11079 -4438 11137 -4432
rect 12193 -4398 12251 -4392
rect 12193 -4432 12205 -4398
rect 12239 -4401 12251 -4398
rect 12571 -4398 12629 -4392
rect 12571 -4401 12583 -4398
rect 12239 -4429 12583 -4401
rect 12239 -4432 12251 -4429
rect 12193 -4438 12251 -4432
rect 12571 -4432 12583 -4429
rect 12617 -4401 12629 -4398
rect 13195 -4398 13253 -4392
rect 13195 -4401 13207 -4398
rect 12617 -4429 13207 -4401
rect 12617 -4432 12629 -4429
rect 12571 -4438 12629 -4432
rect 13195 -4432 13207 -4429
rect 13241 -4432 13253 -4398
rect 13195 -4438 13253 -4432
rect 14309 -4398 14367 -4392
rect 14309 -4432 14321 -4398
rect 14355 -4401 14367 -4398
rect 14687 -4398 14745 -4392
rect 14687 -4401 14699 -4398
rect 14355 -4429 14699 -4401
rect 14355 -4432 14367 -4429
rect 14309 -4438 14367 -4432
rect 14687 -4432 14699 -4429
rect 14733 -4401 14745 -4398
rect 15311 -4398 15369 -4392
rect 15311 -4401 15323 -4398
rect 14733 -4429 15323 -4401
rect 14733 -4432 14745 -4429
rect 14687 -4438 14745 -4432
rect 15311 -4432 15323 -4429
rect 15357 -4432 15369 -4398
rect 15311 -4438 15369 -4432
rect 16425 -4398 16483 -4392
rect 16425 -4432 16437 -4398
rect 16471 -4401 16483 -4398
rect 16803 -4398 16861 -4392
rect 16803 -4401 16815 -4398
rect 16471 -4429 16815 -4401
rect 16471 -4432 16483 -4429
rect 16425 -4438 16483 -4432
rect 16803 -4432 16815 -4429
rect 16849 -4401 16861 -4398
rect 17427 -4398 17485 -4392
rect 17427 -4401 17439 -4398
rect 16849 -4429 17439 -4401
rect 16849 -4432 16861 -4429
rect 16803 -4438 16861 -4432
rect 17427 -4432 17439 -4429
rect 17473 -4432 17485 -4398
rect 17427 -4438 17485 -4432
rect 18541 -4398 18599 -4392
rect 18541 -4432 18553 -4398
rect 18587 -4401 18599 -4398
rect 18919 -4398 18977 -4392
rect 18919 -4401 18931 -4398
rect 18587 -4429 18931 -4401
rect 18587 -4432 18599 -4429
rect 18541 -4438 18599 -4432
rect 18919 -4432 18931 -4429
rect 18965 -4401 18977 -4398
rect 19543 -4398 19601 -4392
rect 19543 -4401 19555 -4398
rect 18965 -4429 19555 -4401
rect 18965 -4432 18977 -4429
rect 18919 -4438 18977 -4432
rect 19543 -4432 19555 -4429
rect 19589 -4432 19601 -4398
rect 19543 -4438 19601 -4432
rect 20657 -4398 20715 -4392
rect 20657 -4432 20669 -4398
rect 20703 -4401 20715 -4398
rect 21035 -4398 21093 -4392
rect 21035 -4401 21047 -4398
rect 20703 -4429 21047 -4401
rect 20703 -4432 20715 -4429
rect 20657 -4438 20715 -4432
rect 21035 -4432 21047 -4429
rect 21081 -4401 21093 -4398
rect 21659 -4398 21717 -4392
rect 21659 -4401 21671 -4398
rect 21081 -4429 21671 -4401
rect 21081 -4432 21093 -4429
rect 21035 -4438 21093 -4432
rect 21659 -4432 21671 -4429
rect 21705 -4432 21717 -4398
rect 21659 -4438 21717 -4432
rect 22773 -4398 22831 -4392
rect 22773 -4432 22785 -4398
rect 22819 -4401 22831 -4398
rect 23151 -4398 23209 -4392
rect 23151 -4401 23163 -4398
rect 22819 -4429 23163 -4401
rect 22819 -4432 22831 -4429
rect 22773 -4438 22831 -4432
rect 23151 -4432 23163 -4429
rect 23197 -4401 23209 -4398
rect 23775 -4398 23833 -4392
rect 23775 -4401 23787 -4398
rect 23197 -4429 23787 -4401
rect 23197 -4432 23209 -4429
rect 23151 -4438 23209 -4432
rect 23775 -4432 23787 -4429
rect 23821 -4432 23833 -4398
rect 23775 -4438 23833 -4432
rect 24889 -4398 24947 -4392
rect 24889 -4432 24901 -4398
rect 24935 -4401 24947 -4398
rect 25267 -4398 25325 -4392
rect 25267 -4401 25279 -4398
rect 24935 -4429 25279 -4401
rect 24935 -4432 24947 -4429
rect 24889 -4438 24947 -4432
rect 25267 -4432 25279 -4429
rect 25313 -4401 25325 -4398
rect 25891 -4398 25949 -4392
rect 25891 -4401 25903 -4398
rect 25313 -4429 25903 -4401
rect 25313 -4432 25325 -4429
rect 25267 -4438 25325 -4432
rect 25891 -4432 25903 -4429
rect 25937 -4432 25949 -4398
rect 25891 -4438 25949 -4432
rect 27005 -4398 27063 -4392
rect 27005 -4432 27017 -4398
rect 27051 -4401 27063 -4398
rect 27383 -4398 27441 -4392
rect 27383 -4401 27395 -4398
rect 27051 -4429 27395 -4401
rect 27051 -4432 27063 -4429
rect 27005 -4438 27063 -4432
rect 27383 -4432 27395 -4429
rect 27429 -4401 27441 -4398
rect 28007 -4398 28065 -4392
rect 28007 -4401 28019 -4398
rect 27429 -4429 28019 -4401
rect 27429 -4432 27441 -4429
rect 27383 -4438 27441 -4432
rect 28007 -4432 28019 -4429
rect 28053 -4432 28065 -4398
rect 28007 -4438 28065 -4432
rect 29121 -4398 29179 -4392
rect 29121 -4432 29133 -4398
rect 29167 -4401 29179 -4398
rect 29499 -4398 29557 -4392
rect 29499 -4401 29511 -4398
rect 29167 -4429 29511 -4401
rect 29167 -4432 29179 -4429
rect 29121 -4438 29179 -4432
rect 29499 -4432 29511 -4429
rect 29545 -4401 29557 -4398
rect 30123 -4398 30181 -4392
rect 30123 -4401 30135 -4398
rect 29545 -4429 30135 -4401
rect 29545 -4432 29557 -4429
rect 29499 -4438 29557 -4432
rect 30123 -4432 30135 -4429
rect 30169 -4432 30181 -4398
rect 30123 -4438 30181 -4432
rect 31237 -4398 31295 -4392
rect 31237 -4432 31249 -4398
rect 31283 -4401 31295 -4398
rect 31615 -4398 31673 -4392
rect 31615 -4401 31627 -4398
rect 31283 -4429 31627 -4401
rect 31283 -4432 31295 -4429
rect 31237 -4438 31295 -4432
rect 31615 -4432 31627 -4429
rect 31661 -4401 31673 -4398
rect 32239 -4398 32297 -4392
rect 32239 -4401 32251 -4398
rect 31661 -4429 32251 -4401
rect 31661 -4432 31673 -4429
rect 31615 -4438 31673 -4432
rect 32239 -4432 32251 -4429
rect 32285 -4432 32297 -4398
rect 32239 -4438 32297 -4432
rect -7749 -4495 -7629 -4489
rect -9048 -4534 -8990 -4528
rect -9048 -4568 -9036 -4534
rect -9002 -4537 -8990 -4534
rect -8681 -4534 -8623 -4528
rect -8681 -4537 -8669 -4534
rect -9002 -4565 -8669 -4537
rect -9002 -4568 -8990 -4565
rect -9048 -4574 -8990 -4568
rect -8681 -4568 -8669 -4565
rect -8635 -4537 -8623 -4534
rect -7965 -4534 -7907 -4528
rect -7965 -4537 -7953 -4534
rect -8635 -4565 -7953 -4537
rect -8635 -4568 -8623 -4565
rect -8681 -4574 -8623 -4568
rect -7965 -4568 -7953 -4565
rect -7919 -4568 -7907 -4534
rect -7965 -4574 -7907 -4568
rect -7749 -4539 -7725 -4495
rect -7749 -4573 -7737 -4539
rect -7673 -4547 -7629 -4495
rect -7703 -4573 -7629 -4547
rect -8909 -4606 -8740 -4598
rect -8909 -4658 -8858 -4606
rect -8806 -4658 -8740 -4606
rect -8409 -4602 -8279 -4596
rect -8409 -4636 -8397 -4602
rect -8363 -4636 -8325 -4602
rect -8291 -4605 -8279 -4602
rect -7749 -4602 -7629 -4573
rect -7113 -4507 -7020 -4480
rect -7113 -4559 -7089 -4507
rect -7037 -4559 -7020 -4507
rect -5633 -4495 -5513 -4489
rect -7113 -4581 -7020 -4559
rect -6932 -4534 -6874 -4528
rect -6932 -4568 -6920 -4534
rect -6886 -4537 -6874 -4534
rect -6565 -4534 -6507 -4528
rect -6565 -4537 -6553 -4534
rect -6886 -4565 -6553 -4537
rect -6886 -4568 -6874 -4565
rect -6932 -4574 -6874 -4568
rect -6565 -4568 -6553 -4565
rect -6519 -4537 -6507 -4534
rect -5849 -4534 -5791 -4528
rect -5849 -4537 -5837 -4534
rect -6519 -4565 -5837 -4537
rect -6519 -4568 -6507 -4565
rect -6565 -4574 -6507 -4568
rect -5849 -4568 -5837 -4565
rect -5803 -4568 -5791 -4534
rect -5849 -4574 -5791 -4568
rect -5633 -4539 -5609 -4495
rect -5633 -4573 -5621 -4539
rect -5557 -4547 -5513 -4495
rect -5587 -4573 -5513 -4547
rect -7749 -4605 -7677 -4602
rect -8291 -4633 -7677 -4605
rect -8291 -4636 -8279 -4633
rect -8409 -4642 -8279 -4636
rect -7689 -4636 -7677 -4633
rect -7643 -4605 -7629 -4602
rect -7643 -4636 -7631 -4605
rect -7689 -4642 -7631 -4636
rect -6793 -4606 -6624 -4598
rect -8909 -4667 -8740 -4658
rect -6793 -4658 -6742 -4606
rect -6690 -4658 -6624 -4606
rect -6293 -4602 -6163 -4596
rect -6293 -4636 -6281 -4602
rect -6247 -4636 -6209 -4602
rect -6175 -4605 -6163 -4602
rect -5633 -4602 -5513 -4573
rect -4997 -4507 -4904 -4480
rect -4997 -4559 -4973 -4507
rect -4921 -4559 -4904 -4507
rect -3517 -4495 -3397 -4489
rect -4997 -4581 -4904 -4559
rect -4816 -4534 -4758 -4528
rect -4816 -4568 -4804 -4534
rect -4770 -4537 -4758 -4534
rect -4449 -4534 -4391 -4528
rect -4449 -4537 -4437 -4534
rect -4770 -4565 -4437 -4537
rect -4770 -4568 -4758 -4565
rect -4816 -4574 -4758 -4568
rect -4449 -4568 -4437 -4565
rect -4403 -4537 -4391 -4534
rect -3733 -4534 -3675 -4528
rect -3733 -4537 -3721 -4534
rect -4403 -4565 -3721 -4537
rect -4403 -4568 -4391 -4565
rect -4449 -4574 -4391 -4568
rect -3733 -4568 -3721 -4565
rect -3687 -4568 -3675 -4534
rect -3733 -4574 -3675 -4568
rect -3517 -4539 -3493 -4495
rect -3517 -4573 -3505 -4539
rect -3441 -4547 -3397 -4495
rect -3471 -4573 -3397 -4547
rect -5633 -4605 -5561 -4602
rect -6175 -4633 -5561 -4605
rect -6175 -4636 -6163 -4633
rect -6293 -4642 -6163 -4636
rect -5573 -4636 -5561 -4633
rect -5527 -4605 -5513 -4602
rect -5527 -4636 -5515 -4605
rect -5573 -4642 -5515 -4636
rect -4677 -4606 -4508 -4598
rect -6793 -4667 -6624 -4658
rect -4677 -4658 -4626 -4606
rect -4574 -4658 -4508 -4606
rect -4177 -4602 -4047 -4596
rect -4177 -4636 -4165 -4602
rect -4131 -4636 -4093 -4602
rect -4059 -4605 -4047 -4602
rect -3517 -4602 -3397 -4573
rect -2881 -4507 -2788 -4480
rect -2881 -4559 -2857 -4507
rect -2805 -4559 -2788 -4507
rect -1401 -4495 -1281 -4489
rect -2881 -4581 -2788 -4559
rect -2700 -4534 -2642 -4528
rect -2700 -4568 -2688 -4534
rect -2654 -4537 -2642 -4534
rect -2333 -4534 -2275 -4528
rect -2333 -4537 -2321 -4534
rect -2654 -4565 -2321 -4537
rect -2654 -4568 -2642 -4565
rect -2700 -4574 -2642 -4568
rect -2333 -4568 -2321 -4565
rect -2287 -4537 -2275 -4534
rect -1617 -4534 -1559 -4528
rect -1617 -4537 -1605 -4534
rect -2287 -4565 -1605 -4537
rect -2287 -4568 -2275 -4565
rect -2333 -4574 -2275 -4568
rect -1617 -4568 -1605 -4565
rect -1571 -4568 -1559 -4534
rect -1617 -4574 -1559 -4568
rect -1401 -4539 -1377 -4495
rect -1401 -4573 -1389 -4539
rect -1325 -4547 -1281 -4495
rect -1355 -4573 -1281 -4547
rect -3517 -4605 -3445 -4602
rect -4059 -4633 -3445 -4605
rect -4059 -4636 -4047 -4633
rect -4177 -4642 -4047 -4636
rect -3457 -4636 -3445 -4633
rect -3411 -4605 -3397 -4602
rect -3411 -4636 -3399 -4605
rect -3457 -4642 -3399 -4636
rect -2561 -4606 -2392 -4598
rect -4677 -4667 -4508 -4658
rect -2561 -4658 -2510 -4606
rect -2458 -4658 -2392 -4606
rect -2061 -4602 -1931 -4596
rect -2061 -4636 -2049 -4602
rect -2015 -4636 -1977 -4602
rect -1943 -4605 -1931 -4602
rect -1401 -4602 -1281 -4573
rect -765 -4507 -672 -4480
rect -765 -4559 -741 -4507
rect -689 -4559 -672 -4507
rect 715 -4495 835 -4489
rect -765 -4581 -672 -4559
rect -584 -4534 -526 -4528
rect -584 -4568 -572 -4534
rect -538 -4537 -526 -4534
rect -217 -4534 -159 -4528
rect -217 -4537 -205 -4534
rect -538 -4565 -205 -4537
rect -538 -4568 -526 -4565
rect -584 -4574 -526 -4568
rect -217 -4568 -205 -4565
rect -171 -4537 -159 -4534
rect 499 -4534 557 -4528
rect 499 -4537 511 -4534
rect -171 -4565 511 -4537
rect -171 -4568 -159 -4565
rect -217 -4574 -159 -4568
rect 499 -4568 511 -4565
rect 545 -4568 557 -4534
rect 499 -4574 557 -4568
rect 715 -4539 739 -4495
rect 715 -4573 727 -4539
rect 791 -4547 835 -4495
rect 761 -4573 835 -4547
rect -1401 -4605 -1329 -4602
rect -1943 -4633 -1329 -4605
rect -1943 -4636 -1931 -4633
rect -2061 -4642 -1931 -4636
rect -1341 -4636 -1329 -4633
rect -1295 -4605 -1281 -4602
rect -1295 -4636 -1283 -4605
rect -1341 -4642 -1283 -4636
rect -445 -4606 -276 -4598
rect -2561 -4667 -2392 -4658
rect -445 -4658 -394 -4606
rect -342 -4658 -276 -4606
rect 55 -4602 185 -4596
rect 55 -4636 67 -4602
rect 101 -4636 139 -4602
rect 173 -4605 185 -4602
rect 715 -4602 835 -4573
rect 1351 -4507 1444 -4480
rect 1351 -4559 1375 -4507
rect 1427 -4559 1444 -4507
rect 2831 -4495 2951 -4489
rect 1351 -4581 1444 -4559
rect 1532 -4534 1590 -4528
rect 1532 -4568 1544 -4534
rect 1578 -4537 1590 -4534
rect 1899 -4534 1957 -4528
rect 1899 -4537 1911 -4534
rect 1578 -4565 1911 -4537
rect 1578 -4568 1590 -4565
rect 1532 -4574 1590 -4568
rect 1899 -4568 1911 -4565
rect 1945 -4537 1957 -4534
rect 2615 -4534 2673 -4528
rect 2615 -4537 2627 -4534
rect 1945 -4565 2627 -4537
rect 1945 -4568 1957 -4565
rect 1899 -4574 1957 -4568
rect 2615 -4568 2627 -4565
rect 2661 -4568 2673 -4534
rect 2615 -4574 2673 -4568
rect 2831 -4539 2855 -4495
rect 2831 -4573 2843 -4539
rect 2907 -4547 2951 -4495
rect 2877 -4573 2951 -4547
rect 715 -4605 787 -4602
rect 173 -4633 787 -4605
rect 173 -4636 185 -4633
rect 55 -4642 185 -4636
rect 775 -4636 787 -4633
rect 821 -4605 835 -4602
rect 821 -4636 833 -4605
rect 775 -4642 833 -4636
rect 1671 -4606 1840 -4598
rect -445 -4667 -276 -4658
rect 1671 -4658 1722 -4606
rect 1774 -4658 1840 -4606
rect 2171 -4602 2301 -4596
rect 2171 -4636 2183 -4602
rect 2217 -4636 2255 -4602
rect 2289 -4605 2301 -4602
rect 2831 -4602 2951 -4573
rect 3467 -4507 3560 -4480
rect 3467 -4559 3491 -4507
rect 3543 -4559 3560 -4507
rect 4947 -4495 5067 -4489
rect 3467 -4581 3560 -4559
rect 3648 -4534 3706 -4528
rect 3648 -4568 3660 -4534
rect 3694 -4537 3706 -4534
rect 4015 -4534 4073 -4528
rect 4015 -4537 4027 -4534
rect 3694 -4565 4027 -4537
rect 3694 -4568 3706 -4565
rect 3648 -4574 3706 -4568
rect 4015 -4568 4027 -4565
rect 4061 -4537 4073 -4534
rect 4731 -4534 4789 -4528
rect 4731 -4537 4743 -4534
rect 4061 -4565 4743 -4537
rect 4061 -4568 4073 -4565
rect 4015 -4574 4073 -4568
rect 4731 -4568 4743 -4565
rect 4777 -4568 4789 -4534
rect 4731 -4574 4789 -4568
rect 4947 -4539 4971 -4495
rect 4947 -4573 4959 -4539
rect 5023 -4547 5067 -4495
rect 4993 -4573 5067 -4547
rect 2831 -4605 2903 -4602
rect 2289 -4633 2903 -4605
rect 2289 -4636 2301 -4633
rect 2171 -4642 2301 -4636
rect 2891 -4636 2903 -4633
rect 2937 -4605 2951 -4602
rect 2937 -4636 2949 -4605
rect 2891 -4642 2949 -4636
rect 3787 -4606 3956 -4598
rect 1671 -4667 1840 -4658
rect 3787 -4658 3838 -4606
rect 3890 -4658 3956 -4606
rect 4287 -4602 4417 -4596
rect 4287 -4636 4299 -4602
rect 4333 -4636 4371 -4602
rect 4405 -4605 4417 -4602
rect 4947 -4602 5067 -4573
rect 5583 -4507 5676 -4480
rect 5583 -4559 5607 -4507
rect 5659 -4559 5676 -4507
rect 7063 -4495 7183 -4489
rect 5583 -4581 5676 -4559
rect 5764 -4534 5822 -4528
rect 5764 -4568 5776 -4534
rect 5810 -4537 5822 -4534
rect 6131 -4534 6189 -4528
rect 6131 -4537 6143 -4534
rect 5810 -4565 6143 -4537
rect 5810 -4568 5822 -4565
rect 5764 -4574 5822 -4568
rect 6131 -4568 6143 -4565
rect 6177 -4537 6189 -4534
rect 6847 -4534 6905 -4528
rect 6847 -4537 6859 -4534
rect 6177 -4565 6859 -4537
rect 6177 -4568 6189 -4565
rect 6131 -4574 6189 -4568
rect 6847 -4568 6859 -4565
rect 6893 -4568 6905 -4534
rect 6847 -4574 6905 -4568
rect 7063 -4539 7087 -4495
rect 7063 -4573 7075 -4539
rect 7139 -4547 7183 -4495
rect 7109 -4573 7183 -4547
rect 4947 -4605 5019 -4602
rect 4405 -4633 5019 -4605
rect 4405 -4636 4417 -4633
rect 4287 -4642 4417 -4636
rect 5007 -4636 5019 -4633
rect 5053 -4605 5067 -4602
rect 5053 -4636 5065 -4605
rect 5007 -4642 5065 -4636
rect 5903 -4606 6072 -4598
rect 3787 -4667 3956 -4658
rect 5903 -4658 5954 -4606
rect 6006 -4658 6072 -4606
rect 6403 -4602 6533 -4596
rect 6403 -4636 6415 -4602
rect 6449 -4636 6487 -4602
rect 6521 -4605 6533 -4602
rect 7063 -4602 7183 -4573
rect 7699 -4507 7792 -4480
rect 7699 -4559 7723 -4507
rect 7775 -4559 7792 -4507
rect 9179 -4495 9299 -4489
rect 7699 -4581 7792 -4559
rect 7880 -4534 7938 -4528
rect 7880 -4568 7892 -4534
rect 7926 -4537 7938 -4534
rect 8247 -4534 8305 -4528
rect 8247 -4537 8259 -4534
rect 7926 -4565 8259 -4537
rect 7926 -4568 7938 -4565
rect 7880 -4574 7938 -4568
rect 8247 -4568 8259 -4565
rect 8293 -4537 8305 -4534
rect 8963 -4534 9021 -4528
rect 8963 -4537 8975 -4534
rect 8293 -4565 8975 -4537
rect 8293 -4568 8305 -4565
rect 8247 -4574 8305 -4568
rect 8963 -4568 8975 -4565
rect 9009 -4568 9021 -4534
rect 8963 -4574 9021 -4568
rect 9179 -4539 9203 -4495
rect 9179 -4573 9191 -4539
rect 9255 -4547 9299 -4495
rect 9225 -4573 9299 -4547
rect 7063 -4605 7135 -4602
rect 6521 -4633 7135 -4605
rect 6521 -4636 6533 -4633
rect 6403 -4642 6533 -4636
rect 7123 -4636 7135 -4633
rect 7169 -4605 7183 -4602
rect 7169 -4636 7181 -4605
rect 7123 -4642 7181 -4636
rect 8019 -4606 8188 -4598
rect 5903 -4667 6072 -4658
rect 8019 -4658 8070 -4606
rect 8122 -4658 8188 -4606
rect 8519 -4602 8649 -4596
rect 8519 -4636 8531 -4602
rect 8565 -4636 8603 -4602
rect 8637 -4605 8649 -4602
rect 9179 -4602 9299 -4573
rect 9815 -4507 9908 -4480
rect 9815 -4559 9839 -4507
rect 9891 -4559 9908 -4507
rect 11295 -4495 11415 -4489
rect 9815 -4581 9908 -4559
rect 9996 -4534 10054 -4528
rect 9996 -4568 10008 -4534
rect 10042 -4537 10054 -4534
rect 10363 -4534 10421 -4528
rect 10363 -4537 10375 -4534
rect 10042 -4565 10375 -4537
rect 10042 -4568 10054 -4565
rect 9996 -4574 10054 -4568
rect 10363 -4568 10375 -4565
rect 10409 -4537 10421 -4534
rect 11079 -4534 11137 -4528
rect 11079 -4537 11091 -4534
rect 10409 -4565 11091 -4537
rect 10409 -4568 10421 -4565
rect 10363 -4574 10421 -4568
rect 11079 -4568 11091 -4565
rect 11125 -4568 11137 -4534
rect 11079 -4574 11137 -4568
rect 11295 -4539 11319 -4495
rect 11295 -4573 11307 -4539
rect 11371 -4547 11415 -4495
rect 11341 -4573 11415 -4547
rect 9179 -4605 9251 -4602
rect 8637 -4633 9251 -4605
rect 8637 -4636 8649 -4633
rect 8519 -4642 8649 -4636
rect 9239 -4636 9251 -4633
rect 9285 -4605 9299 -4602
rect 9285 -4636 9297 -4605
rect 9239 -4642 9297 -4636
rect 10135 -4606 10304 -4598
rect 8019 -4667 8188 -4658
rect 10135 -4658 10186 -4606
rect 10238 -4658 10304 -4606
rect 10635 -4602 10765 -4596
rect 10635 -4636 10647 -4602
rect 10681 -4636 10719 -4602
rect 10753 -4605 10765 -4602
rect 11295 -4602 11415 -4573
rect 11931 -4507 12024 -4480
rect 11931 -4559 11955 -4507
rect 12007 -4559 12024 -4507
rect 13411 -4495 13531 -4489
rect 11931 -4581 12024 -4559
rect 12112 -4534 12170 -4528
rect 12112 -4568 12124 -4534
rect 12158 -4537 12170 -4534
rect 12479 -4534 12537 -4528
rect 12479 -4537 12491 -4534
rect 12158 -4565 12491 -4537
rect 12158 -4568 12170 -4565
rect 12112 -4574 12170 -4568
rect 12479 -4568 12491 -4565
rect 12525 -4537 12537 -4534
rect 13195 -4534 13253 -4528
rect 13195 -4537 13207 -4534
rect 12525 -4565 13207 -4537
rect 12525 -4568 12537 -4565
rect 12479 -4574 12537 -4568
rect 13195 -4568 13207 -4565
rect 13241 -4568 13253 -4534
rect 13195 -4574 13253 -4568
rect 13411 -4539 13435 -4495
rect 13411 -4573 13423 -4539
rect 13487 -4547 13531 -4495
rect 13457 -4573 13531 -4547
rect 11295 -4605 11367 -4602
rect 10753 -4633 11367 -4605
rect 10753 -4636 10765 -4633
rect 10635 -4642 10765 -4636
rect 11355 -4636 11367 -4633
rect 11401 -4605 11415 -4602
rect 11401 -4636 11413 -4605
rect 11355 -4642 11413 -4636
rect 12251 -4606 12420 -4598
rect 10135 -4667 10304 -4658
rect 12251 -4658 12302 -4606
rect 12354 -4658 12420 -4606
rect 12751 -4602 12881 -4596
rect 12751 -4636 12763 -4602
rect 12797 -4636 12835 -4602
rect 12869 -4605 12881 -4602
rect 13411 -4602 13531 -4573
rect 14047 -4507 14140 -4480
rect 14047 -4559 14071 -4507
rect 14123 -4559 14140 -4507
rect 15527 -4495 15647 -4489
rect 14047 -4581 14140 -4559
rect 14228 -4534 14286 -4528
rect 14228 -4568 14240 -4534
rect 14274 -4537 14286 -4534
rect 14595 -4534 14653 -4528
rect 14595 -4537 14607 -4534
rect 14274 -4565 14607 -4537
rect 14274 -4568 14286 -4565
rect 14228 -4574 14286 -4568
rect 14595 -4568 14607 -4565
rect 14641 -4537 14653 -4534
rect 15311 -4534 15369 -4528
rect 15311 -4537 15323 -4534
rect 14641 -4565 15323 -4537
rect 14641 -4568 14653 -4565
rect 14595 -4574 14653 -4568
rect 15311 -4568 15323 -4565
rect 15357 -4568 15369 -4534
rect 15311 -4574 15369 -4568
rect 15527 -4539 15551 -4495
rect 15527 -4573 15539 -4539
rect 15603 -4547 15647 -4495
rect 15573 -4573 15647 -4547
rect 13411 -4605 13483 -4602
rect 12869 -4633 13483 -4605
rect 12869 -4636 12881 -4633
rect 12751 -4642 12881 -4636
rect 13471 -4636 13483 -4633
rect 13517 -4605 13531 -4602
rect 13517 -4636 13529 -4605
rect 13471 -4642 13529 -4636
rect 14367 -4606 14536 -4598
rect 12251 -4667 12420 -4658
rect 14367 -4658 14418 -4606
rect 14470 -4658 14536 -4606
rect 14867 -4602 14997 -4596
rect 14867 -4636 14879 -4602
rect 14913 -4636 14951 -4602
rect 14985 -4605 14997 -4602
rect 15527 -4602 15647 -4573
rect 16163 -4507 16256 -4480
rect 16163 -4559 16187 -4507
rect 16239 -4559 16256 -4507
rect 17643 -4495 17763 -4489
rect 16163 -4581 16256 -4559
rect 16344 -4534 16402 -4528
rect 16344 -4568 16356 -4534
rect 16390 -4537 16402 -4534
rect 16711 -4534 16769 -4528
rect 16711 -4537 16723 -4534
rect 16390 -4565 16723 -4537
rect 16390 -4568 16402 -4565
rect 16344 -4574 16402 -4568
rect 16711 -4568 16723 -4565
rect 16757 -4537 16769 -4534
rect 17427 -4534 17485 -4528
rect 17427 -4537 17439 -4534
rect 16757 -4565 17439 -4537
rect 16757 -4568 16769 -4565
rect 16711 -4574 16769 -4568
rect 17427 -4568 17439 -4565
rect 17473 -4568 17485 -4534
rect 17427 -4574 17485 -4568
rect 17643 -4539 17667 -4495
rect 17643 -4573 17655 -4539
rect 17719 -4547 17763 -4495
rect 17689 -4573 17763 -4547
rect 15527 -4605 15599 -4602
rect 14985 -4633 15599 -4605
rect 14985 -4636 14997 -4633
rect 14867 -4642 14997 -4636
rect 15587 -4636 15599 -4633
rect 15633 -4605 15647 -4602
rect 15633 -4636 15645 -4605
rect 15587 -4642 15645 -4636
rect 16483 -4606 16652 -4598
rect 14367 -4667 14536 -4658
rect 16483 -4658 16534 -4606
rect 16586 -4658 16652 -4606
rect 16983 -4602 17113 -4596
rect 16983 -4636 16995 -4602
rect 17029 -4636 17067 -4602
rect 17101 -4605 17113 -4602
rect 17643 -4602 17763 -4573
rect 18279 -4507 18372 -4480
rect 18279 -4559 18303 -4507
rect 18355 -4559 18372 -4507
rect 19759 -4495 19879 -4489
rect 18279 -4581 18372 -4559
rect 18460 -4534 18518 -4528
rect 18460 -4568 18472 -4534
rect 18506 -4537 18518 -4534
rect 18827 -4534 18885 -4528
rect 18827 -4537 18839 -4534
rect 18506 -4565 18839 -4537
rect 18506 -4568 18518 -4565
rect 18460 -4574 18518 -4568
rect 18827 -4568 18839 -4565
rect 18873 -4537 18885 -4534
rect 19543 -4534 19601 -4528
rect 19543 -4537 19555 -4534
rect 18873 -4565 19555 -4537
rect 18873 -4568 18885 -4565
rect 18827 -4574 18885 -4568
rect 19543 -4568 19555 -4565
rect 19589 -4568 19601 -4534
rect 19543 -4574 19601 -4568
rect 19759 -4539 19783 -4495
rect 19759 -4573 19771 -4539
rect 19835 -4547 19879 -4495
rect 19805 -4573 19879 -4547
rect 17643 -4605 17715 -4602
rect 17101 -4633 17715 -4605
rect 17101 -4636 17113 -4633
rect 16983 -4642 17113 -4636
rect 17703 -4636 17715 -4633
rect 17749 -4605 17763 -4602
rect 17749 -4636 17761 -4605
rect 17703 -4642 17761 -4636
rect 18599 -4606 18768 -4598
rect 16483 -4667 16652 -4658
rect 18599 -4658 18650 -4606
rect 18702 -4658 18768 -4606
rect 19099 -4602 19229 -4596
rect 19099 -4636 19111 -4602
rect 19145 -4636 19183 -4602
rect 19217 -4605 19229 -4602
rect 19759 -4602 19879 -4573
rect 20395 -4507 20488 -4480
rect 20395 -4559 20419 -4507
rect 20471 -4559 20488 -4507
rect 21875 -4495 21995 -4489
rect 20395 -4581 20488 -4559
rect 20576 -4534 20634 -4528
rect 20576 -4568 20588 -4534
rect 20622 -4537 20634 -4534
rect 20943 -4534 21001 -4528
rect 20943 -4537 20955 -4534
rect 20622 -4565 20955 -4537
rect 20622 -4568 20634 -4565
rect 20576 -4574 20634 -4568
rect 20943 -4568 20955 -4565
rect 20989 -4537 21001 -4534
rect 21659 -4534 21717 -4528
rect 21659 -4537 21671 -4534
rect 20989 -4565 21671 -4537
rect 20989 -4568 21001 -4565
rect 20943 -4574 21001 -4568
rect 21659 -4568 21671 -4565
rect 21705 -4568 21717 -4534
rect 21659 -4574 21717 -4568
rect 21875 -4539 21899 -4495
rect 21875 -4573 21887 -4539
rect 21951 -4547 21995 -4495
rect 21921 -4573 21995 -4547
rect 19759 -4605 19831 -4602
rect 19217 -4633 19831 -4605
rect 19217 -4636 19229 -4633
rect 19099 -4642 19229 -4636
rect 19819 -4636 19831 -4633
rect 19865 -4605 19879 -4602
rect 19865 -4636 19877 -4605
rect 19819 -4642 19877 -4636
rect 20715 -4606 20884 -4598
rect 18599 -4667 18768 -4658
rect 20715 -4658 20766 -4606
rect 20818 -4658 20884 -4606
rect 21215 -4602 21345 -4596
rect 21215 -4636 21227 -4602
rect 21261 -4636 21299 -4602
rect 21333 -4605 21345 -4602
rect 21875 -4602 21995 -4573
rect 22511 -4507 22604 -4480
rect 22511 -4559 22535 -4507
rect 22587 -4559 22604 -4507
rect 23991 -4495 24111 -4489
rect 22511 -4581 22604 -4559
rect 22692 -4534 22750 -4528
rect 22692 -4568 22704 -4534
rect 22738 -4537 22750 -4534
rect 23059 -4534 23117 -4528
rect 23059 -4537 23071 -4534
rect 22738 -4565 23071 -4537
rect 22738 -4568 22750 -4565
rect 22692 -4574 22750 -4568
rect 23059 -4568 23071 -4565
rect 23105 -4537 23117 -4534
rect 23775 -4534 23833 -4528
rect 23775 -4537 23787 -4534
rect 23105 -4565 23787 -4537
rect 23105 -4568 23117 -4565
rect 23059 -4574 23117 -4568
rect 23775 -4568 23787 -4565
rect 23821 -4568 23833 -4534
rect 23775 -4574 23833 -4568
rect 23991 -4539 24015 -4495
rect 23991 -4573 24003 -4539
rect 24067 -4547 24111 -4495
rect 24037 -4573 24111 -4547
rect 21875 -4605 21947 -4602
rect 21333 -4633 21947 -4605
rect 21333 -4636 21345 -4633
rect 21215 -4642 21345 -4636
rect 21935 -4636 21947 -4633
rect 21981 -4605 21995 -4602
rect 21981 -4636 21993 -4605
rect 21935 -4642 21993 -4636
rect 22831 -4606 23000 -4598
rect 20715 -4667 20884 -4658
rect 22831 -4658 22882 -4606
rect 22934 -4658 23000 -4606
rect 23331 -4602 23461 -4596
rect 23331 -4636 23343 -4602
rect 23377 -4636 23415 -4602
rect 23449 -4605 23461 -4602
rect 23991 -4602 24111 -4573
rect 24627 -4507 24720 -4480
rect 24627 -4559 24651 -4507
rect 24703 -4559 24720 -4507
rect 26107 -4495 26227 -4489
rect 24627 -4581 24720 -4559
rect 24808 -4534 24866 -4528
rect 24808 -4568 24820 -4534
rect 24854 -4537 24866 -4534
rect 25175 -4534 25233 -4528
rect 25175 -4537 25187 -4534
rect 24854 -4565 25187 -4537
rect 24854 -4568 24866 -4565
rect 24808 -4574 24866 -4568
rect 25175 -4568 25187 -4565
rect 25221 -4537 25233 -4534
rect 25891 -4534 25949 -4528
rect 25891 -4537 25903 -4534
rect 25221 -4565 25903 -4537
rect 25221 -4568 25233 -4565
rect 25175 -4574 25233 -4568
rect 25891 -4568 25903 -4565
rect 25937 -4568 25949 -4534
rect 25891 -4574 25949 -4568
rect 26107 -4539 26131 -4495
rect 26107 -4573 26119 -4539
rect 26183 -4547 26227 -4495
rect 26153 -4573 26227 -4547
rect 23991 -4605 24063 -4602
rect 23449 -4633 24063 -4605
rect 23449 -4636 23461 -4633
rect 23331 -4642 23461 -4636
rect 24051 -4636 24063 -4633
rect 24097 -4605 24111 -4602
rect 24097 -4636 24109 -4605
rect 24051 -4642 24109 -4636
rect 24947 -4606 25116 -4598
rect 22831 -4667 23000 -4658
rect 24947 -4658 24998 -4606
rect 25050 -4658 25116 -4606
rect 25447 -4602 25577 -4596
rect 25447 -4636 25459 -4602
rect 25493 -4636 25531 -4602
rect 25565 -4605 25577 -4602
rect 26107 -4602 26227 -4573
rect 26743 -4507 26836 -4480
rect 26743 -4559 26767 -4507
rect 26819 -4559 26836 -4507
rect 28223 -4495 28343 -4489
rect 26743 -4581 26836 -4559
rect 26924 -4534 26982 -4528
rect 26924 -4568 26936 -4534
rect 26970 -4537 26982 -4534
rect 27291 -4534 27349 -4528
rect 27291 -4537 27303 -4534
rect 26970 -4565 27303 -4537
rect 26970 -4568 26982 -4565
rect 26924 -4574 26982 -4568
rect 27291 -4568 27303 -4565
rect 27337 -4537 27349 -4534
rect 28007 -4534 28065 -4528
rect 28007 -4537 28019 -4534
rect 27337 -4565 28019 -4537
rect 27337 -4568 27349 -4565
rect 27291 -4574 27349 -4568
rect 28007 -4568 28019 -4565
rect 28053 -4568 28065 -4534
rect 28007 -4574 28065 -4568
rect 28223 -4539 28247 -4495
rect 28223 -4573 28235 -4539
rect 28299 -4547 28343 -4495
rect 28269 -4573 28343 -4547
rect 26107 -4605 26179 -4602
rect 25565 -4633 26179 -4605
rect 25565 -4636 25577 -4633
rect 25447 -4642 25577 -4636
rect 26167 -4636 26179 -4633
rect 26213 -4605 26227 -4602
rect 26213 -4636 26225 -4605
rect 26167 -4642 26225 -4636
rect 27063 -4606 27232 -4598
rect 24947 -4667 25116 -4658
rect 27063 -4658 27114 -4606
rect 27166 -4658 27232 -4606
rect 27563 -4602 27693 -4596
rect 27563 -4636 27575 -4602
rect 27609 -4636 27647 -4602
rect 27681 -4605 27693 -4602
rect 28223 -4602 28343 -4573
rect 28859 -4507 28952 -4480
rect 28859 -4559 28883 -4507
rect 28935 -4559 28952 -4507
rect 30339 -4495 30459 -4489
rect 28859 -4581 28952 -4559
rect 29040 -4534 29098 -4528
rect 29040 -4568 29052 -4534
rect 29086 -4537 29098 -4534
rect 29407 -4534 29465 -4528
rect 29407 -4537 29419 -4534
rect 29086 -4565 29419 -4537
rect 29086 -4568 29098 -4565
rect 29040 -4574 29098 -4568
rect 29407 -4568 29419 -4565
rect 29453 -4537 29465 -4534
rect 30123 -4534 30181 -4528
rect 30123 -4537 30135 -4534
rect 29453 -4565 30135 -4537
rect 29453 -4568 29465 -4565
rect 29407 -4574 29465 -4568
rect 30123 -4568 30135 -4565
rect 30169 -4568 30181 -4534
rect 30123 -4574 30181 -4568
rect 30339 -4539 30363 -4495
rect 30339 -4573 30351 -4539
rect 30415 -4547 30459 -4495
rect 30385 -4573 30459 -4547
rect 28223 -4605 28295 -4602
rect 27681 -4633 28295 -4605
rect 27681 -4636 27693 -4633
rect 27563 -4642 27693 -4636
rect 28283 -4636 28295 -4633
rect 28329 -4605 28343 -4602
rect 28329 -4636 28341 -4605
rect 28283 -4642 28341 -4636
rect 29179 -4606 29348 -4598
rect 27063 -4667 27232 -4658
rect 29179 -4658 29230 -4606
rect 29282 -4658 29348 -4606
rect 29679 -4602 29809 -4596
rect 29679 -4636 29691 -4602
rect 29725 -4636 29763 -4602
rect 29797 -4605 29809 -4602
rect 30339 -4602 30459 -4573
rect 30975 -4507 31068 -4480
rect 30975 -4559 30999 -4507
rect 31051 -4559 31068 -4507
rect 32455 -4495 32575 -4489
rect 30975 -4581 31068 -4559
rect 31156 -4534 31214 -4528
rect 31156 -4568 31168 -4534
rect 31202 -4537 31214 -4534
rect 31523 -4534 31581 -4528
rect 31523 -4537 31535 -4534
rect 31202 -4565 31535 -4537
rect 31202 -4568 31214 -4565
rect 31156 -4574 31214 -4568
rect 31523 -4568 31535 -4565
rect 31569 -4537 31581 -4534
rect 32239 -4534 32297 -4528
rect 32239 -4537 32251 -4534
rect 31569 -4565 32251 -4537
rect 31569 -4568 31581 -4565
rect 31523 -4574 31581 -4568
rect 32239 -4568 32251 -4565
rect 32285 -4568 32297 -4534
rect 32239 -4574 32297 -4568
rect 32455 -4539 32479 -4495
rect 32455 -4573 32467 -4539
rect 32531 -4547 32575 -4495
rect 32501 -4573 32575 -4547
rect 30339 -4605 30411 -4602
rect 29797 -4633 30411 -4605
rect 29797 -4636 29809 -4633
rect 29679 -4642 29809 -4636
rect 30399 -4636 30411 -4633
rect 30445 -4605 30459 -4602
rect 30445 -4636 30457 -4605
rect 30399 -4642 30457 -4636
rect 31295 -4606 31464 -4598
rect 29179 -4667 29348 -4658
rect 31295 -4658 31346 -4606
rect 31398 -4658 31464 -4606
rect 31795 -4602 31925 -4596
rect 31795 -4636 31807 -4602
rect 31841 -4636 31879 -4602
rect 31913 -4605 31925 -4602
rect 32455 -4602 32575 -4573
rect 33091 -4507 33184 -4480
rect 33091 -4559 33115 -4507
rect 33167 -4559 33184 -4507
rect 33091 -4581 33184 -4559
rect 32455 -4605 32527 -4602
rect 31913 -4633 32527 -4605
rect 31913 -4636 31925 -4633
rect 31795 -4642 31925 -4636
rect 32515 -4636 32527 -4633
rect 32561 -4605 32575 -4602
rect 32561 -4636 32573 -4605
rect 32515 -4642 32573 -4636
rect 31295 -4667 31464 -4658
rect -9158 -4772 33162 -4741
rect -9158 -4806 -9129 -4772
rect -9095 -4806 -9037 -4772
rect -9003 -4806 -8945 -4772
rect -8911 -4806 -8853 -4772
rect -8819 -4806 -8761 -4772
rect -8727 -4806 -8669 -4772
rect -8635 -4806 -8577 -4772
rect -8543 -4806 -8485 -4772
rect -8451 -4806 -8393 -4772
rect -8359 -4806 -8301 -4772
rect -8267 -4806 -8209 -4772
rect -8175 -4806 -8117 -4772
rect -8083 -4806 -8025 -4772
rect -7991 -4806 -7933 -4772
rect -7899 -4806 -7841 -4772
rect -7807 -4806 -7749 -4772
rect -7715 -4806 -7657 -4772
rect -7623 -4806 -7565 -4772
rect -7531 -4806 -7473 -4772
rect -7439 -4806 -7381 -4772
rect -7347 -4806 -7289 -4772
rect -7255 -4806 -7197 -4772
rect -7163 -4806 -7105 -4772
rect -7071 -4806 -7013 -4772
rect -6979 -4806 -6921 -4772
rect -6887 -4806 -6829 -4772
rect -6795 -4806 -6737 -4772
rect -6703 -4806 -6645 -4772
rect -6611 -4806 -6553 -4772
rect -6519 -4806 -6461 -4772
rect -6427 -4806 -6369 -4772
rect -6335 -4806 -6277 -4772
rect -6243 -4806 -6185 -4772
rect -6151 -4806 -6093 -4772
rect -6059 -4806 -6001 -4772
rect -5967 -4806 -5909 -4772
rect -5875 -4806 -5817 -4772
rect -5783 -4806 -5725 -4772
rect -5691 -4806 -5633 -4772
rect -5599 -4806 -5541 -4772
rect -5507 -4806 -5449 -4772
rect -5415 -4806 -5357 -4772
rect -5323 -4806 -5265 -4772
rect -5231 -4806 -5173 -4772
rect -5139 -4806 -5081 -4772
rect -5047 -4806 -4989 -4772
rect -4955 -4806 -4897 -4772
rect -4863 -4806 -4805 -4772
rect -4771 -4806 -4713 -4772
rect -4679 -4806 -4621 -4772
rect -4587 -4806 -4529 -4772
rect -4495 -4806 -4437 -4772
rect -4403 -4806 -4345 -4772
rect -4311 -4806 -4253 -4772
rect -4219 -4806 -4161 -4772
rect -4127 -4806 -4069 -4772
rect -4035 -4806 -3977 -4772
rect -3943 -4806 -3885 -4772
rect -3851 -4806 -3793 -4772
rect -3759 -4806 -3701 -4772
rect -3667 -4806 -3609 -4772
rect -3575 -4806 -3517 -4772
rect -3483 -4806 -3425 -4772
rect -3391 -4806 -3333 -4772
rect -3299 -4806 -3241 -4772
rect -3207 -4806 -3149 -4772
rect -3115 -4806 -3057 -4772
rect -3023 -4806 -2965 -4772
rect -2931 -4806 -2873 -4772
rect -2839 -4806 -2781 -4772
rect -2747 -4806 -2689 -4772
rect -2655 -4806 -2597 -4772
rect -2563 -4806 -2505 -4772
rect -2471 -4806 -2413 -4772
rect -2379 -4806 -2321 -4772
rect -2287 -4806 -2229 -4772
rect -2195 -4806 -2137 -4772
rect -2103 -4806 -2045 -4772
rect -2011 -4806 -1953 -4772
rect -1919 -4806 -1861 -4772
rect -1827 -4806 -1769 -4772
rect -1735 -4806 -1677 -4772
rect -1643 -4806 -1585 -4772
rect -1551 -4806 -1493 -4772
rect -1459 -4806 -1401 -4772
rect -1367 -4806 -1309 -4772
rect -1275 -4806 -1217 -4772
rect -1183 -4806 -1125 -4772
rect -1091 -4806 -1033 -4772
rect -999 -4806 -941 -4772
rect -907 -4806 -849 -4772
rect -815 -4806 -757 -4772
rect -723 -4806 -665 -4772
rect -631 -4806 -573 -4772
rect -539 -4806 -481 -4772
rect -447 -4806 -389 -4772
rect -355 -4806 -297 -4772
rect -263 -4806 -205 -4772
rect -171 -4806 -113 -4772
rect -79 -4806 -21 -4772
rect 13 -4806 71 -4772
rect 105 -4806 163 -4772
rect 197 -4806 255 -4772
rect 289 -4806 347 -4772
rect 381 -4806 439 -4772
rect 473 -4806 531 -4772
rect 565 -4806 623 -4772
rect 657 -4806 715 -4772
rect 749 -4806 807 -4772
rect 841 -4806 899 -4772
rect 933 -4806 991 -4772
rect 1025 -4806 1083 -4772
rect 1117 -4806 1175 -4772
rect 1209 -4806 1267 -4772
rect 1301 -4806 1359 -4772
rect 1393 -4806 1451 -4772
rect 1485 -4806 1543 -4772
rect 1577 -4806 1635 -4772
rect 1669 -4806 1727 -4772
rect 1761 -4806 1819 -4772
rect 1853 -4806 1911 -4772
rect 1945 -4806 2003 -4772
rect 2037 -4806 2095 -4772
rect 2129 -4806 2187 -4772
rect 2221 -4806 2279 -4772
rect 2313 -4806 2371 -4772
rect 2405 -4806 2463 -4772
rect 2497 -4806 2555 -4772
rect 2589 -4806 2647 -4772
rect 2681 -4806 2739 -4772
rect 2773 -4806 2831 -4772
rect 2865 -4806 2923 -4772
rect 2957 -4806 3015 -4772
rect 3049 -4806 3107 -4772
rect 3141 -4806 3199 -4772
rect 3233 -4806 3291 -4772
rect 3325 -4806 3383 -4772
rect 3417 -4806 3475 -4772
rect 3509 -4806 3567 -4772
rect 3601 -4806 3659 -4772
rect 3693 -4806 3751 -4772
rect 3785 -4806 3843 -4772
rect 3877 -4806 3935 -4772
rect 3969 -4806 4027 -4772
rect 4061 -4806 4119 -4772
rect 4153 -4806 4211 -4772
rect 4245 -4806 4303 -4772
rect 4337 -4806 4395 -4772
rect 4429 -4806 4487 -4772
rect 4521 -4806 4579 -4772
rect 4613 -4806 4671 -4772
rect 4705 -4806 4763 -4772
rect 4797 -4806 4855 -4772
rect 4889 -4806 4947 -4772
rect 4981 -4806 5039 -4772
rect 5073 -4806 5131 -4772
rect 5165 -4806 5223 -4772
rect 5257 -4806 5315 -4772
rect 5349 -4806 5407 -4772
rect 5441 -4806 5499 -4772
rect 5533 -4806 5591 -4772
rect 5625 -4806 5683 -4772
rect 5717 -4806 5775 -4772
rect 5809 -4806 5867 -4772
rect 5901 -4806 5959 -4772
rect 5993 -4806 6051 -4772
rect 6085 -4806 6143 -4772
rect 6177 -4806 6235 -4772
rect 6269 -4806 6327 -4772
rect 6361 -4806 6419 -4772
rect 6453 -4806 6511 -4772
rect 6545 -4806 6603 -4772
rect 6637 -4806 6695 -4772
rect 6729 -4806 6787 -4772
rect 6821 -4806 6879 -4772
rect 6913 -4806 6971 -4772
rect 7005 -4806 7063 -4772
rect 7097 -4806 7155 -4772
rect 7189 -4806 7247 -4772
rect 7281 -4806 7339 -4772
rect 7373 -4806 7431 -4772
rect 7465 -4806 7523 -4772
rect 7557 -4806 7615 -4772
rect 7649 -4806 7707 -4772
rect 7741 -4806 7799 -4772
rect 7833 -4806 7891 -4772
rect 7925 -4806 7983 -4772
rect 8017 -4806 8075 -4772
rect 8109 -4806 8167 -4772
rect 8201 -4806 8259 -4772
rect 8293 -4806 8351 -4772
rect 8385 -4806 8443 -4772
rect 8477 -4806 8535 -4772
rect 8569 -4806 8627 -4772
rect 8661 -4806 8719 -4772
rect 8753 -4806 8811 -4772
rect 8845 -4806 8903 -4772
rect 8937 -4806 8995 -4772
rect 9029 -4806 9087 -4772
rect 9121 -4806 9179 -4772
rect 9213 -4806 9271 -4772
rect 9305 -4806 9363 -4772
rect 9397 -4806 9455 -4772
rect 9489 -4806 9547 -4772
rect 9581 -4806 9639 -4772
rect 9673 -4806 9731 -4772
rect 9765 -4806 9823 -4772
rect 9857 -4806 9915 -4772
rect 9949 -4806 10007 -4772
rect 10041 -4806 10099 -4772
rect 10133 -4806 10191 -4772
rect 10225 -4806 10283 -4772
rect 10317 -4806 10375 -4772
rect 10409 -4806 10467 -4772
rect 10501 -4806 10559 -4772
rect 10593 -4806 10651 -4772
rect 10685 -4806 10743 -4772
rect 10777 -4806 10835 -4772
rect 10869 -4806 10927 -4772
rect 10961 -4806 11019 -4772
rect 11053 -4806 11111 -4772
rect 11145 -4806 11203 -4772
rect 11237 -4806 11295 -4772
rect 11329 -4806 11387 -4772
rect 11421 -4806 11479 -4772
rect 11513 -4806 11571 -4772
rect 11605 -4806 11663 -4772
rect 11697 -4806 11755 -4772
rect 11789 -4806 11847 -4772
rect 11881 -4806 11939 -4772
rect 11973 -4806 12031 -4772
rect 12065 -4806 12123 -4772
rect 12157 -4806 12215 -4772
rect 12249 -4806 12307 -4772
rect 12341 -4806 12399 -4772
rect 12433 -4806 12491 -4772
rect 12525 -4806 12583 -4772
rect 12617 -4806 12675 -4772
rect 12709 -4806 12767 -4772
rect 12801 -4806 12859 -4772
rect 12893 -4806 12951 -4772
rect 12985 -4806 13043 -4772
rect 13077 -4806 13135 -4772
rect 13169 -4806 13227 -4772
rect 13261 -4806 13319 -4772
rect 13353 -4806 13411 -4772
rect 13445 -4806 13503 -4772
rect 13537 -4806 13595 -4772
rect 13629 -4806 13687 -4772
rect 13721 -4806 13779 -4772
rect 13813 -4806 13871 -4772
rect 13905 -4806 13963 -4772
rect 13997 -4806 14055 -4772
rect 14089 -4806 14147 -4772
rect 14181 -4806 14239 -4772
rect 14273 -4806 14331 -4772
rect 14365 -4806 14423 -4772
rect 14457 -4806 14515 -4772
rect 14549 -4806 14607 -4772
rect 14641 -4806 14699 -4772
rect 14733 -4806 14791 -4772
rect 14825 -4806 14883 -4772
rect 14917 -4806 14975 -4772
rect 15009 -4806 15067 -4772
rect 15101 -4806 15159 -4772
rect 15193 -4806 15251 -4772
rect 15285 -4806 15343 -4772
rect 15377 -4806 15435 -4772
rect 15469 -4806 15527 -4772
rect 15561 -4806 15619 -4772
rect 15653 -4806 15711 -4772
rect 15745 -4806 15803 -4772
rect 15837 -4806 15895 -4772
rect 15929 -4806 15987 -4772
rect 16021 -4806 16079 -4772
rect 16113 -4806 16171 -4772
rect 16205 -4806 16263 -4772
rect 16297 -4806 16355 -4772
rect 16389 -4806 16447 -4772
rect 16481 -4806 16539 -4772
rect 16573 -4806 16631 -4772
rect 16665 -4806 16723 -4772
rect 16757 -4806 16815 -4772
rect 16849 -4806 16907 -4772
rect 16941 -4806 16999 -4772
rect 17033 -4806 17091 -4772
rect 17125 -4806 17183 -4772
rect 17217 -4806 17275 -4772
rect 17309 -4806 17367 -4772
rect 17401 -4806 17459 -4772
rect 17493 -4806 17551 -4772
rect 17585 -4806 17643 -4772
rect 17677 -4806 17735 -4772
rect 17769 -4806 17827 -4772
rect 17861 -4806 17919 -4772
rect 17953 -4806 18011 -4772
rect 18045 -4806 18103 -4772
rect 18137 -4806 18195 -4772
rect 18229 -4806 18287 -4772
rect 18321 -4806 18379 -4772
rect 18413 -4806 18471 -4772
rect 18505 -4806 18563 -4772
rect 18597 -4806 18655 -4772
rect 18689 -4806 18747 -4772
rect 18781 -4806 18839 -4772
rect 18873 -4806 18931 -4772
rect 18965 -4806 19023 -4772
rect 19057 -4806 19115 -4772
rect 19149 -4806 19207 -4772
rect 19241 -4806 19299 -4772
rect 19333 -4806 19391 -4772
rect 19425 -4806 19483 -4772
rect 19517 -4806 19575 -4772
rect 19609 -4806 19667 -4772
rect 19701 -4806 19759 -4772
rect 19793 -4806 19851 -4772
rect 19885 -4806 19943 -4772
rect 19977 -4806 20035 -4772
rect 20069 -4806 20127 -4772
rect 20161 -4806 20219 -4772
rect 20253 -4806 20311 -4772
rect 20345 -4806 20403 -4772
rect 20437 -4806 20495 -4772
rect 20529 -4806 20587 -4772
rect 20621 -4806 20679 -4772
rect 20713 -4806 20771 -4772
rect 20805 -4806 20863 -4772
rect 20897 -4806 20955 -4772
rect 20989 -4806 21047 -4772
rect 21081 -4806 21139 -4772
rect 21173 -4806 21231 -4772
rect 21265 -4806 21323 -4772
rect 21357 -4806 21415 -4772
rect 21449 -4806 21507 -4772
rect 21541 -4806 21599 -4772
rect 21633 -4806 21691 -4772
rect 21725 -4806 21783 -4772
rect 21817 -4806 21875 -4772
rect 21909 -4806 21967 -4772
rect 22001 -4806 22059 -4772
rect 22093 -4806 22151 -4772
rect 22185 -4806 22243 -4772
rect 22277 -4806 22335 -4772
rect 22369 -4806 22427 -4772
rect 22461 -4806 22519 -4772
rect 22553 -4806 22611 -4772
rect 22645 -4806 22703 -4772
rect 22737 -4806 22795 -4772
rect 22829 -4806 22887 -4772
rect 22921 -4806 22979 -4772
rect 23013 -4806 23071 -4772
rect 23105 -4806 23163 -4772
rect 23197 -4806 23255 -4772
rect 23289 -4806 23347 -4772
rect 23381 -4806 23439 -4772
rect 23473 -4806 23531 -4772
rect 23565 -4806 23623 -4772
rect 23657 -4806 23715 -4772
rect 23749 -4806 23807 -4772
rect 23841 -4806 23899 -4772
rect 23933 -4806 23991 -4772
rect 24025 -4806 24083 -4772
rect 24117 -4806 24175 -4772
rect 24209 -4806 24267 -4772
rect 24301 -4806 24359 -4772
rect 24393 -4806 24451 -4772
rect 24485 -4806 24543 -4772
rect 24577 -4806 24635 -4772
rect 24669 -4806 24727 -4772
rect 24761 -4806 24819 -4772
rect 24853 -4806 24911 -4772
rect 24945 -4806 25003 -4772
rect 25037 -4806 25095 -4772
rect 25129 -4806 25187 -4772
rect 25221 -4806 25279 -4772
rect 25313 -4806 25371 -4772
rect 25405 -4806 25463 -4772
rect 25497 -4806 25555 -4772
rect 25589 -4806 25647 -4772
rect 25681 -4806 25739 -4772
rect 25773 -4806 25831 -4772
rect 25865 -4806 25923 -4772
rect 25957 -4806 26015 -4772
rect 26049 -4806 26107 -4772
rect 26141 -4806 26199 -4772
rect 26233 -4806 26291 -4772
rect 26325 -4806 26383 -4772
rect 26417 -4806 26475 -4772
rect 26509 -4806 26567 -4772
rect 26601 -4806 26659 -4772
rect 26693 -4806 26751 -4772
rect 26785 -4806 26843 -4772
rect 26877 -4806 26935 -4772
rect 26969 -4806 27027 -4772
rect 27061 -4806 27119 -4772
rect 27153 -4806 27211 -4772
rect 27245 -4806 27303 -4772
rect 27337 -4806 27395 -4772
rect 27429 -4806 27487 -4772
rect 27521 -4806 27579 -4772
rect 27613 -4806 27671 -4772
rect 27705 -4806 27763 -4772
rect 27797 -4806 27855 -4772
rect 27889 -4806 27947 -4772
rect 27981 -4806 28039 -4772
rect 28073 -4806 28131 -4772
rect 28165 -4806 28223 -4772
rect 28257 -4806 28315 -4772
rect 28349 -4806 28407 -4772
rect 28441 -4806 28499 -4772
rect 28533 -4806 28591 -4772
rect 28625 -4806 28683 -4772
rect 28717 -4806 28775 -4772
rect 28809 -4806 28867 -4772
rect 28901 -4806 28959 -4772
rect 28993 -4806 29051 -4772
rect 29085 -4806 29143 -4772
rect 29177 -4806 29235 -4772
rect 29269 -4806 29327 -4772
rect 29361 -4806 29419 -4772
rect 29453 -4806 29511 -4772
rect 29545 -4806 29603 -4772
rect 29637 -4806 29695 -4772
rect 29729 -4806 29787 -4772
rect 29821 -4806 29879 -4772
rect 29913 -4806 29971 -4772
rect 30005 -4806 30063 -4772
rect 30097 -4806 30155 -4772
rect 30189 -4806 30247 -4772
rect 30281 -4806 30339 -4772
rect 30373 -4806 30431 -4772
rect 30465 -4806 30523 -4772
rect 30557 -4806 30615 -4772
rect 30649 -4806 30707 -4772
rect 30741 -4806 30799 -4772
rect 30833 -4806 30891 -4772
rect 30925 -4806 30983 -4772
rect 31017 -4806 31075 -4772
rect 31109 -4806 31167 -4772
rect 31201 -4806 31259 -4772
rect 31293 -4806 31351 -4772
rect 31385 -4806 31443 -4772
rect 31477 -4806 31535 -4772
rect 31569 -4806 31627 -4772
rect 31661 -4806 31719 -4772
rect 31753 -4806 31811 -4772
rect 31845 -4806 31903 -4772
rect 31937 -4806 31995 -4772
rect 32029 -4806 32087 -4772
rect 32121 -4806 32179 -4772
rect 32213 -4806 32271 -4772
rect 32305 -4806 32363 -4772
rect 32397 -4806 32455 -4772
rect 32489 -4806 32547 -4772
rect 32581 -4806 32639 -4772
rect 32673 -4806 32731 -4772
rect 32765 -4806 32823 -4772
rect 32857 -4806 32915 -4772
rect 32949 -4806 33007 -4772
rect 33041 -4806 33099 -4772
rect 33133 -4806 33162 -4772
rect -9158 -4837 33162 -4806
rect 4216 -7518 7872 -7506
rect 4216 -25771 4254 -7518
rect 4290 -7519 7872 -7518
rect 4290 -7635 7798 -7519
rect 4290 -9011 4369 -7635
rect 4403 -9011 6027 -7635
rect 6061 -9011 7685 -7635
rect 7719 -9011 7798 -7635
rect 4290 -9145 7798 -9011
rect 4290 -10521 4369 -9145
rect 4403 -10521 6027 -9145
rect 6061 -10521 7685 -9145
rect 7719 -10521 7798 -9145
rect 4290 -10655 7798 -10521
rect 4290 -12031 4369 -10655
rect 4403 -12031 6027 -10655
rect 6061 -12031 7685 -10655
rect 7719 -12031 7798 -10655
rect 4290 -12165 7798 -12031
rect 4290 -13541 4369 -12165
rect 4403 -12977 6027 -12165
rect 6061 -12977 7685 -12165
rect 4403 -13467 5413 -12977
rect 6710 -13467 7685 -12977
rect 4403 -13541 6027 -13467
rect 6061 -13541 7685 -13467
rect 7719 -13541 7798 -12165
rect 4290 -13675 7798 -13541
rect 4290 -15051 4369 -13675
rect 4403 -15051 6027 -13675
rect 6061 -15051 7685 -13675
rect 7719 -15051 7798 -13675
rect 4290 -15185 7798 -15051
rect 4290 -16561 4369 -15185
rect 4403 -16561 6027 -15185
rect 6061 -16561 7685 -15185
rect 7719 -16561 7798 -15185
rect 4290 -16695 7798 -16561
rect 4290 -18071 4369 -16695
rect 4403 -18071 6027 -16695
rect 6061 -18071 7685 -16695
rect 7719 -18071 7798 -16695
rect 4290 -18205 7798 -18071
rect 4290 -19581 4369 -18205
rect 4403 -19581 6027 -18205
rect 6061 -19581 7685 -18205
rect 7719 -19581 7798 -18205
rect 4290 -19715 7798 -19581
rect 4290 -21091 4369 -19715
rect 4403 -21091 6027 -19715
rect 6061 -21091 7685 -19715
rect 7719 -21091 7798 -19715
rect 4290 -21225 7798 -21091
rect 4290 -22601 4369 -21225
rect 4403 -22601 6027 -21225
rect 6061 -22601 7685 -21225
rect 7719 -22601 7798 -21225
rect 4290 -22735 7798 -22601
rect 4290 -24111 4369 -22735
rect 4403 -24111 6027 -22735
rect 6061 -24111 7685 -22735
rect 7719 -24111 7798 -22735
rect 4290 -24245 7798 -24111
rect 4290 -25621 4369 -24245
rect 4403 -25621 6027 -24245
rect 6061 -25621 7685 -24245
rect 7719 -25621 7798 -24245
rect 4290 -25771 7798 -25621
rect 4216 -25814 4246 -25771
rect 7834 -25808 7872 -7519
rect 17834 -7518 21491 -7510
rect 12789 -7563 14478 -7554
rect 9858 -7594 10405 -7568
rect 9858 -7628 10176 -7594
rect 10210 -7628 10405 -7594
rect 9858 -7689 10405 -7628
rect 9858 -7850 9897 -7689
rect 9960 -7690 10286 -7689
rect 9960 -7849 10023 -7690
rect 10103 -7849 10174 -7690
rect 10254 -7848 10286 -7690
rect 10366 -7848 10405 -7689
rect 10254 -7849 10405 -7848
rect 9960 -7850 10405 -7849
rect 9858 -7922 10405 -7850
rect 9858 -7956 10176 -7922
rect 10210 -7956 10405 -7922
rect 9858 -7982 10405 -7956
rect 12788 -7595 14478 -7563
rect 12788 -7629 13064 -7595
rect 13098 -7629 13322 -7595
rect 13356 -7629 13580 -7595
rect 13614 -7629 13838 -7595
rect 13872 -7629 14096 -7595
rect 14130 -7629 14478 -7595
rect 12788 -7656 14478 -7629
rect 12788 -7882 12896 -7656
rect 14455 -7882 14478 -7656
rect 12788 -7884 14341 -7882
rect 14454 -7884 14478 -7882
rect 12788 -7923 14478 -7884
rect 12788 -7957 13064 -7923
rect 13098 -7957 13322 -7923
rect 13356 -7957 13580 -7923
rect 13614 -7957 13838 -7923
rect 13872 -7957 14096 -7923
rect 14130 -7957 14478 -7923
rect 12788 -7992 14478 -7957
rect 12789 -7995 14478 -7992
rect 10071 -8567 10197 -8559
rect 10071 -8628 10093 -8567
rect 10173 -8628 10197 -8567
rect 8984 -8654 9262 -8635
rect 8984 -8967 9002 -8654
rect 9241 -8967 9262 -8654
rect 10071 -8788 10197 -8628
rect 10071 -8849 10094 -8788
rect 10174 -8849 10197 -8788
rect 10071 -8942 10197 -8849
rect 8984 -8986 9262 -8967
rect 10070 -9321 10197 -8942
rect 12747 -8571 12873 -8558
rect 12747 -8654 12767 -8571
rect 12865 -8654 12873 -8571
rect 12747 -8766 12873 -8654
rect 12747 -8849 12767 -8766
rect 12865 -8849 12873 -8766
rect 12747 -8953 12873 -8849
rect 15403 -8571 15529 -8559
rect 15403 -8654 15419 -8571
rect 15517 -8654 15529 -8571
rect 15403 -8766 15529 -8654
rect 15403 -8849 15419 -8766
rect 15517 -8849 15529 -8766
rect 15403 -8942 15529 -8849
rect 12747 -9318 12872 -8953
rect 7986 -9349 8378 -9343
rect 10070 -9349 10198 -9321
rect 7986 -9485 10198 -9349
rect 12743 -9366 12872 -9318
rect 12743 -9445 12755 -9366
rect 12850 -9445 12872 -9366
rect 12743 -9462 12872 -9445
rect 7986 -10613 8378 -9485
rect 7986 -10831 8042 -10613
rect 8288 -10831 8378 -10613
rect 7986 -10849 8378 -10831
rect 8857 -9525 9017 -9524
rect 10070 -9525 10196 -9485
rect 11307 -9525 11467 -9524
rect 8857 -9564 11467 -9525
rect 8857 -9598 9242 -9564
rect 9276 -9598 9500 -9564
rect 9534 -9598 9758 -9564
rect 9792 -9598 10016 -9564
rect 10050 -9598 10274 -9564
rect 10308 -9598 10532 -9564
rect 10566 -9598 10790 -9564
rect 10824 -9598 11048 -9564
rect 11082 -9598 11467 -9564
rect 8857 -9624 11467 -9598
rect 8857 -9853 9017 -9624
rect 11307 -9853 11467 -9624
rect 8857 -9874 11467 -9853
rect 8857 -9908 9242 -9874
rect 9276 -9908 9500 -9874
rect 9534 -9908 9758 -9874
rect 9792 -9908 10016 -9874
rect 10050 -9908 10274 -9874
rect 10308 -9908 10532 -9874
rect 10566 -9908 10790 -9874
rect 10824 -9908 11048 -9874
rect 11082 -9908 11467 -9874
rect 8857 -9982 11467 -9908
rect 8857 -10016 9242 -9982
rect 9276 -10016 9500 -9982
rect 9534 -10016 9758 -9982
rect 9792 -10016 10016 -9982
rect 10050 -10016 10274 -9982
rect 10308 -10016 10532 -9982
rect 10566 -10016 10790 -9982
rect 10824 -10016 11048 -9982
rect 11082 -10016 11467 -9982
rect 8857 -10044 11467 -10016
rect 8857 -10263 9017 -10044
rect 11307 -10263 11467 -10044
rect 8857 -10292 11467 -10263
rect 8857 -10326 9242 -10292
rect 9276 -10326 9500 -10292
rect 9534 -10326 9758 -10292
rect 9792 -10326 10016 -10292
rect 10050 -10326 10274 -10292
rect 10308 -10326 10532 -10292
rect 10566 -10326 10790 -10292
rect 10824 -10326 11048 -10292
rect 11082 -10326 11467 -10292
rect 8857 -10400 11467 -10326
rect 8857 -10434 9242 -10400
rect 9276 -10434 9500 -10400
rect 9534 -10434 9758 -10400
rect 9792 -10434 10016 -10400
rect 10050 -10434 10274 -10400
rect 10308 -10434 10532 -10400
rect 10566 -10434 10790 -10400
rect 10824 -10434 11048 -10400
rect 11082 -10434 11467 -10400
rect 8857 -10454 11467 -10434
rect 8857 -10693 9017 -10454
rect 11307 -10693 11467 -10454
rect 8857 -10710 11467 -10693
rect 8857 -10744 9242 -10710
rect 9276 -10744 9500 -10710
rect 9534 -10744 9758 -10710
rect 9792 -10744 10016 -10710
rect 10050 -10744 10274 -10710
rect 10308 -10744 10532 -10710
rect 10566 -10744 10790 -10710
rect 10824 -10744 11048 -10710
rect 11082 -10744 11467 -10710
rect 8857 -10818 11467 -10744
rect 8857 -10852 9242 -10818
rect 9276 -10852 9500 -10818
rect 9534 -10852 9758 -10818
rect 9792 -10852 10016 -10818
rect 10050 -10852 10274 -10818
rect 10308 -10852 10532 -10818
rect 10566 -10852 10790 -10818
rect 10824 -10852 11048 -10818
rect 11082 -10852 11467 -10818
rect 8857 -10884 11467 -10852
rect 8857 -11103 9017 -10884
rect 11307 -11103 11467 -10884
rect 8857 -11128 11467 -11103
rect 8857 -11162 9242 -11128
rect 9276 -11162 9500 -11128
rect 9534 -11162 9758 -11128
rect 9792 -11162 10016 -11128
rect 10050 -11162 10274 -11128
rect 10308 -11162 10532 -11128
rect 10566 -11162 10790 -11128
rect 10824 -11162 11048 -11128
rect 11082 -11162 11467 -11128
rect 8857 -11236 11467 -11162
rect 8857 -11270 9242 -11236
rect 9276 -11270 9500 -11236
rect 9534 -11270 9758 -11236
rect 9792 -11270 10016 -11236
rect 10050 -11270 10274 -11236
rect 10308 -11270 10532 -11236
rect 10566 -11270 10790 -11236
rect 10824 -11270 11048 -11236
rect 11082 -11270 11467 -11236
rect 8857 -11294 11467 -11270
rect 8857 -11523 9017 -11294
rect 11307 -11523 11467 -11294
rect 8857 -11546 11467 -11523
rect 8857 -11580 9242 -11546
rect 9276 -11580 9500 -11546
rect 9534 -11580 9758 -11546
rect 9792 -11580 10016 -11546
rect 10050 -11580 10274 -11546
rect 10308 -11580 10532 -11546
rect 10566 -11580 10790 -11546
rect 10824 -11580 11048 -11546
rect 11082 -11580 11467 -11546
rect 8857 -11654 11467 -11580
rect 8857 -11688 9242 -11654
rect 9276 -11688 9500 -11654
rect 9534 -11688 9758 -11654
rect 9792 -11688 10016 -11654
rect 10050 -11688 10274 -11654
rect 10308 -11688 10532 -11654
rect 10566 -11688 10790 -11654
rect 10824 -11688 11048 -11654
rect 11082 -11688 11467 -11654
rect 8857 -11714 11467 -11688
rect 8857 -11933 9017 -11714
rect 11307 -11933 11467 -11714
rect 8857 -11964 11467 -11933
rect 8857 -11998 9242 -11964
rect 9276 -11998 9500 -11964
rect 9534 -11998 9758 -11964
rect 9792 -11998 10016 -11964
rect 10050 -11998 10274 -11964
rect 10308 -11998 10532 -11964
rect 10566 -11998 10790 -11964
rect 10824 -11998 11048 -11964
rect 11082 -11998 11467 -11964
rect 8857 -12072 11467 -11998
rect 8857 -12106 9242 -12072
rect 9276 -12106 9500 -12072
rect 9534 -12106 9758 -12072
rect 9792 -12106 10016 -12072
rect 10050 -12106 10274 -12072
rect 10308 -12106 10532 -12072
rect 10566 -12106 10790 -12072
rect 10824 -12106 11048 -12072
rect 11082 -12106 11467 -12072
rect 8857 -12124 11467 -12106
rect 8857 -12354 9017 -12124
rect 11307 -12354 11467 -12124
rect 8857 -12382 11467 -12354
rect 8857 -12416 9242 -12382
rect 9276 -12416 9500 -12382
rect 9534 -12416 9758 -12382
rect 9792 -12416 10016 -12382
rect 10050 -12416 10274 -12382
rect 10308 -12416 10532 -12382
rect 10566 -12416 10790 -12382
rect 10824 -12416 11048 -12382
rect 11082 -12416 11467 -12382
rect 8857 -12484 11467 -12416
rect 11527 -9525 11687 -9524
rect 12746 -9525 12872 -9462
rect 15402 -9355 15529 -8942
rect 16398 -8669 16699 -8645
rect 16398 -8990 16433 -8669
rect 16655 -8990 16699 -8669
rect 16398 -9016 16699 -8990
rect 16644 -9253 17522 -9209
rect 15402 -9366 15542 -9355
rect 15402 -9445 15428 -9366
rect 15523 -9445 15542 -9366
rect 15402 -9462 15542 -9445
rect 16644 -9431 16664 -9253
rect 16832 -9429 17324 -9253
rect 17486 -9429 17522 -9253
rect 16832 -9431 17522 -9429
rect 14190 -9524 14350 -9523
rect 15402 -9524 15528 -9462
rect 16644 -9463 17522 -9431
rect 16640 -9524 16800 -9523
rect 13977 -9525 14137 -9524
rect 11527 -9564 14137 -9525
rect 11527 -9598 11912 -9564
rect 11946 -9598 12170 -9564
rect 12204 -9598 12428 -9564
rect 12462 -9598 12686 -9564
rect 12720 -9598 12944 -9564
rect 12978 -9598 13202 -9564
rect 13236 -9598 13460 -9564
rect 13494 -9598 13718 -9564
rect 13752 -9598 14137 -9564
rect 11527 -9624 14137 -9598
rect 11527 -9853 11687 -9624
rect 13977 -9853 14137 -9624
rect 11527 -9874 14137 -9853
rect 11527 -9908 11912 -9874
rect 11946 -9908 12170 -9874
rect 12204 -9908 12428 -9874
rect 12462 -9908 12686 -9874
rect 12720 -9908 12944 -9874
rect 12978 -9908 13202 -9874
rect 13236 -9908 13460 -9874
rect 13494 -9908 13718 -9874
rect 13752 -9908 14137 -9874
rect 11527 -9982 14137 -9908
rect 11527 -10016 11912 -9982
rect 11946 -10016 12170 -9982
rect 12204 -10016 12428 -9982
rect 12462 -10016 12686 -9982
rect 12720 -10016 12944 -9982
rect 12978 -10016 13202 -9982
rect 13236 -10016 13460 -9982
rect 13494 -10016 13718 -9982
rect 13752 -10016 14137 -9982
rect 11527 -10044 14137 -10016
rect 11527 -10263 11687 -10044
rect 13977 -10263 14137 -10044
rect 11527 -10292 14137 -10263
rect 11527 -10326 11912 -10292
rect 11946 -10326 12170 -10292
rect 12204 -10326 12428 -10292
rect 12462 -10326 12686 -10292
rect 12720 -10326 12944 -10292
rect 12978 -10326 13202 -10292
rect 13236 -10326 13460 -10292
rect 13494 -10326 13718 -10292
rect 13752 -10326 14137 -10292
rect 11527 -10400 14137 -10326
rect 11527 -10434 11912 -10400
rect 11946 -10434 12170 -10400
rect 12204 -10434 12428 -10400
rect 12462 -10434 12686 -10400
rect 12720 -10434 12944 -10400
rect 12978 -10434 13202 -10400
rect 13236 -10434 13460 -10400
rect 13494 -10434 13718 -10400
rect 13752 -10434 14137 -10400
rect 11527 -10454 14137 -10434
rect 11527 -10693 11687 -10454
rect 13977 -10693 14137 -10454
rect 11527 -10710 14137 -10693
rect 11527 -10744 11912 -10710
rect 11946 -10744 12170 -10710
rect 12204 -10744 12428 -10710
rect 12462 -10744 12686 -10710
rect 12720 -10744 12944 -10710
rect 12978 -10744 13202 -10710
rect 13236 -10744 13460 -10710
rect 13494 -10744 13718 -10710
rect 13752 -10744 14137 -10710
rect 11527 -10818 14137 -10744
rect 11527 -10852 11912 -10818
rect 11946 -10852 12170 -10818
rect 12204 -10852 12428 -10818
rect 12462 -10852 12686 -10818
rect 12720 -10852 12944 -10818
rect 12978 -10852 13202 -10818
rect 13236 -10852 13460 -10818
rect 13494 -10852 13718 -10818
rect 13752 -10852 14137 -10818
rect 11527 -10884 14137 -10852
rect 11527 -11103 11687 -10884
rect 13977 -11103 14137 -10884
rect 11527 -11128 14137 -11103
rect 11527 -11162 11912 -11128
rect 11946 -11162 12170 -11128
rect 12204 -11162 12428 -11128
rect 12462 -11162 12686 -11128
rect 12720 -11162 12944 -11128
rect 12978 -11162 13202 -11128
rect 13236 -11162 13460 -11128
rect 13494 -11162 13718 -11128
rect 13752 -11162 14137 -11128
rect 11527 -11236 14137 -11162
rect 11527 -11270 11912 -11236
rect 11946 -11270 12170 -11236
rect 12204 -11270 12428 -11236
rect 12462 -11270 12686 -11236
rect 12720 -11270 12944 -11236
rect 12978 -11270 13202 -11236
rect 13236 -11270 13460 -11236
rect 13494 -11270 13718 -11236
rect 13752 -11270 14137 -11236
rect 11527 -11294 14137 -11270
rect 11527 -11523 11687 -11294
rect 13977 -11523 14137 -11294
rect 11527 -11546 14137 -11523
rect 11527 -11580 11912 -11546
rect 11946 -11580 12170 -11546
rect 12204 -11580 12428 -11546
rect 12462 -11580 12686 -11546
rect 12720 -11580 12944 -11546
rect 12978 -11580 13202 -11546
rect 13236 -11580 13460 -11546
rect 13494 -11580 13718 -11546
rect 13752 -11580 14137 -11546
rect 11527 -11654 14137 -11580
rect 11527 -11688 11912 -11654
rect 11946 -11688 12170 -11654
rect 12204 -11688 12428 -11654
rect 12462 -11688 12686 -11654
rect 12720 -11688 12944 -11654
rect 12978 -11688 13202 -11654
rect 13236 -11688 13460 -11654
rect 13494 -11688 13718 -11654
rect 13752 -11688 14137 -11654
rect 11527 -11714 14137 -11688
rect 11527 -11933 11687 -11714
rect 13977 -11933 14137 -11714
rect 11527 -11964 14137 -11933
rect 11527 -11998 11912 -11964
rect 11946 -11998 12170 -11964
rect 12204 -11998 12428 -11964
rect 12462 -11998 12686 -11964
rect 12720 -11998 12944 -11964
rect 12978 -11998 13202 -11964
rect 13236 -11998 13460 -11964
rect 13494 -11998 13718 -11964
rect 13752 -11998 14137 -11964
rect 11527 -12072 14137 -11998
rect 11527 -12106 11912 -12072
rect 11946 -12106 12170 -12072
rect 12204 -12106 12428 -12072
rect 12462 -12106 12686 -12072
rect 12720 -12106 12944 -12072
rect 12978 -12106 13202 -12072
rect 13236 -12106 13460 -12072
rect 13494 -12106 13718 -12072
rect 13752 -12106 14137 -12072
rect 11527 -12124 14137 -12106
rect 11527 -12354 11687 -12124
rect 13977 -12354 14137 -12124
rect 11527 -12382 14137 -12354
rect 11527 -12416 11912 -12382
rect 11946 -12416 12170 -12382
rect 12204 -12416 12428 -12382
rect 12462 -12416 12686 -12382
rect 12720 -12416 12944 -12382
rect 12978 -12416 13202 -12382
rect 13236 -12416 13460 -12382
rect 13494 -12416 13718 -12382
rect 13752 -12416 14137 -12382
rect 11527 -12484 14137 -12416
rect 14190 -9563 16800 -9524
rect 14190 -9597 14575 -9563
rect 14609 -9597 14833 -9563
rect 14867 -9597 15091 -9563
rect 15125 -9597 15349 -9563
rect 15383 -9597 15607 -9563
rect 15641 -9597 15865 -9563
rect 15899 -9597 16123 -9563
rect 16157 -9597 16381 -9563
rect 16415 -9597 16800 -9563
rect 14190 -9623 16800 -9597
rect 14190 -9852 14350 -9623
rect 16640 -9852 16800 -9623
rect 14190 -9873 16800 -9852
rect 14190 -9907 14575 -9873
rect 14609 -9907 14833 -9873
rect 14867 -9907 15091 -9873
rect 15125 -9907 15349 -9873
rect 15383 -9907 15607 -9873
rect 15641 -9907 15865 -9873
rect 15899 -9907 16123 -9873
rect 16157 -9907 16381 -9873
rect 16415 -9907 16800 -9873
rect 14190 -9981 16800 -9907
rect 14190 -10015 14575 -9981
rect 14609 -10015 14833 -9981
rect 14867 -10015 15091 -9981
rect 15125 -10015 15349 -9981
rect 15383 -10015 15607 -9981
rect 15641 -10015 15865 -9981
rect 15899 -10015 16123 -9981
rect 16157 -10015 16381 -9981
rect 16415 -10015 16800 -9981
rect 14190 -10043 16800 -10015
rect 14190 -10262 14350 -10043
rect 16640 -10262 16800 -10043
rect 14190 -10291 16800 -10262
rect 14190 -10325 14575 -10291
rect 14609 -10325 14833 -10291
rect 14867 -10325 15091 -10291
rect 15125 -10325 15349 -10291
rect 15383 -10325 15607 -10291
rect 15641 -10325 15865 -10291
rect 15899 -10325 16123 -10291
rect 16157 -10325 16381 -10291
rect 16415 -10325 16800 -10291
rect 14190 -10399 16800 -10325
rect 14190 -10433 14575 -10399
rect 14609 -10433 14833 -10399
rect 14867 -10433 15091 -10399
rect 15125 -10433 15349 -10399
rect 15383 -10433 15607 -10399
rect 15641 -10433 15865 -10399
rect 15899 -10433 16123 -10399
rect 16157 -10433 16381 -10399
rect 16415 -10433 16800 -10399
rect 14190 -10453 16800 -10433
rect 14190 -10692 14350 -10453
rect 16640 -10692 16800 -10453
rect 14190 -10709 16800 -10692
rect 14190 -10743 14575 -10709
rect 14609 -10743 14833 -10709
rect 14867 -10743 15091 -10709
rect 15125 -10743 15349 -10709
rect 15383 -10743 15607 -10709
rect 15641 -10743 15865 -10709
rect 15899 -10743 16123 -10709
rect 16157 -10743 16381 -10709
rect 16415 -10743 16800 -10709
rect 14190 -10817 16800 -10743
rect 14190 -10851 14575 -10817
rect 14609 -10851 14833 -10817
rect 14867 -10851 15091 -10817
rect 15125 -10851 15349 -10817
rect 15383 -10851 15607 -10817
rect 15641 -10851 15865 -10817
rect 15899 -10851 16123 -10817
rect 16157 -10851 16381 -10817
rect 16415 -10851 16800 -10817
rect 14190 -10883 16800 -10851
rect 14190 -11102 14350 -10883
rect 16640 -11102 16800 -10883
rect 14190 -11127 16800 -11102
rect 14190 -11161 14575 -11127
rect 14609 -11161 14833 -11127
rect 14867 -11161 15091 -11127
rect 15125 -11161 15349 -11127
rect 15383 -11161 15607 -11127
rect 15641 -11161 15865 -11127
rect 15899 -11161 16123 -11127
rect 16157 -11161 16381 -11127
rect 16415 -11161 16800 -11127
rect 14190 -11235 16800 -11161
rect 14190 -11269 14575 -11235
rect 14609 -11269 14833 -11235
rect 14867 -11269 15091 -11235
rect 15125 -11269 15349 -11235
rect 15383 -11269 15607 -11235
rect 15641 -11269 15865 -11235
rect 15899 -11269 16123 -11235
rect 16157 -11269 16381 -11235
rect 16415 -11269 16800 -11235
rect 14190 -11293 16800 -11269
rect 14190 -11522 14350 -11293
rect 16640 -11522 16800 -11293
rect 14190 -11545 16800 -11522
rect 14190 -11579 14575 -11545
rect 14609 -11579 14833 -11545
rect 14867 -11579 15091 -11545
rect 15125 -11579 15349 -11545
rect 15383 -11579 15607 -11545
rect 15641 -11579 15865 -11545
rect 15899 -11579 16123 -11545
rect 16157 -11579 16381 -11545
rect 16415 -11579 16800 -11545
rect 14190 -11653 16800 -11579
rect 14190 -11687 14575 -11653
rect 14609 -11687 14833 -11653
rect 14867 -11687 15091 -11653
rect 15125 -11687 15349 -11653
rect 15383 -11687 15607 -11653
rect 15641 -11687 15865 -11653
rect 15899 -11687 16123 -11653
rect 16157 -11687 16381 -11653
rect 16415 -11687 16800 -11653
rect 14190 -11713 16800 -11687
rect 14190 -11932 14350 -11713
rect 16640 -11932 16800 -11713
rect 14190 -11963 16800 -11932
rect 14190 -11997 14575 -11963
rect 14609 -11997 14833 -11963
rect 14867 -11997 15091 -11963
rect 15125 -11997 15349 -11963
rect 15383 -11997 15607 -11963
rect 15641 -11997 15865 -11963
rect 15899 -11997 16123 -11963
rect 16157 -11997 16381 -11963
rect 16415 -11997 16800 -11963
rect 14190 -12071 16800 -11997
rect 14190 -12105 14575 -12071
rect 14609 -12105 14833 -12071
rect 14867 -12105 15091 -12071
rect 15125 -12105 15349 -12071
rect 15383 -12105 15607 -12071
rect 15641 -12105 15865 -12071
rect 15899 -12105 16123 -12071
rect 16157 -12105 16381 -12071
rect 16415 -12105 16800 -12071
rect 14190 -12123 16800 -12105
rect 14190 -12353 14350 -12123
rect 16640 -12353 16800 -12123
rect 14190 -12381 16800 -12353
rect 14190 -12415 14575 -12381
rect 14609 -12415 14833 -12381
rect 14867 -12415 15091 -12381
rect 15125 -12415 15349 -12381
rect 15383 -12415 15607 -12381
rect 15641 -12415 15865 -12381
rect 15899 -12415 16123 -12381
rect 16157 -12415 16381 -12381
rect 16415 -12415 16800 -12381
rect 14190 -12483 16800 -12415
rect 17294 -10179 17522 -10163
rect 17294 -10355 17324 -10179
rect 17486 -10355 17522 -10179
rect 10107 -12724 10217 -12484
rect 10107 -12764 10137 -12724
rect 10187 -12764 10217 -12724
rect 10107 -13031 10217 -12764
rect 10107 -13071 10140 -13031
rect 10178 -13071 10217 -13031
rect 10107 -13092 10217 -13071
rect 12777 -12724 12887 -12484
rect 12777 -12764 12807 -12724
rect 12857 -12764 12887 -12724
rect 12777 -13031 12887 -12764
rect 12777 -13071 12810 -13031
rect 12848 -13071 12887 -13031
rect 12777 -13095 12887 -13071
rect 15440 -12723 15550 -12483
rect 15440 -12763 15470 -12723
rect 15520 -12763 15550 -12723
rect 15440 -13031 15550 -12763
rect 15440 -13071 15472 -13031
rect 15510 -13071 15550 -13031
rect 15440 -13086 15550 -13071
rect 9950 -13161 10094 -13153
rect 9950 -13267 9970 -13161
rect 10076 -13267 10094 -13161
rect 9950 -13277 10094 -13267
rect 12616 -13161 12760 -13153
rect 12616 -13267 12634 -13161
rect 12740 -13267 12760 -13161
rect 12616 -13277 12760 -13267
rect 15277 -13161 15423 -13153
rect 15277 -13267 15296 -13161
rect 15402 -13267 15423 -13161
rect 15277 -13278 15423 -13267
rect 17294 -14017 17522 -10355
rect 17290 -14061 17522 -14017
rect 8951 -14220 9229 -14206
rect 8951 -14525 8991 -14220
rect 9174 -14525 9229 -14220
rect 17290 -14237 17324 -14061
rect 17486 -14237 17522 -14061
rect 8951 -14557 9229 -14525
rect 10069 -14249 10195 -14241
rect 10069 -14310 10093 -14249
rect 10173 -14310 10195 -14249
rect 10069 -14470 10195 -14310
rect 10069 -14531 10092 -14470
rect 10172 -14531 10195 -14470
rect 10069 -14538 10195 -14531
rect 12740 -14253 12866 -14240
rect 12740 -14336 12748 -14253
rect 12846 -14336 12866 -14253
rect 12740 -14448 12866 -14336
rect 12740 -14531 12748 -14448
rect 12846 -14531 12866 -14448
rect 12740 -14538 12866 -14531
rect 15411 -14253 15537 -14241
rect 15411 -14336 15423 -14253
rect 15521 -14336 15537 -14253
rect 17290 -14271 17522 -14237
rect 15411 -14448 15537 -14336
rect 15411 -14531 15423 -14448
rect 15521 -14531 15537 -14448
rect 15411 -14538 15537 -14531
rect 8032 -15007 9056 -14973
rect 8032 -15059 8856 -15007
rect 8032 -15235 8070 -15059
rect 8232 -15171 8856 -15059
rect 9014 -15171 9056 -15007
rect 8232 -15193 9056 -15171
rect 10070 -15029 10196 -14538
rect 12746 -15029 12872 -14538
rect 10070 -15057 11718 -15029
rect 10070 -15191 11562 -15057
rect 11680 -15191 11718 -15057
rect 12746 -15067 14302 -15029
rect 12746 -15072 14168 -15067
rect 12743 -15179 14168 -15072
rect 8232 -15235 8268 -15193
rect 8032 -15269 8268 -15235
rect 10070 -15201 11718 -15191
rect 12746 -15191 14168 -15179
rect 14280 -15191 14302 -15067
rect 8857 -15242 9017 -15241
rect 10070 -15242 10196 -15201
rect 12746 -15205 14302 -15191
rect 15402 -15039 15528 -14538
rect 17294 -14987 17522 -14971
rect 17294 -15039 17324 -14987
rect 15402 -15163 17324 -15039
rect 17486 -15163 17522 -14987
rect 15402 -15179 17522 -15163
rect 15402 -15181 17292 -15179
rect 11307 -15242 11467 -15241
rect 8857 -15281 11467 -15242
rect 8857 -15315 9242 -15281
rect 9276 -15315 9500 -15281
rect 9534 -15315 9758 -15281
rect 9792 -15315 10016 -15281
rect 10050 -15315 10274 -15281
rect 10308 -15315 10532 -15281
rect 10566 -15315 10790 -15281
rect 10824 -15315 11048 -15281
rect 11082 -15315 11467 -15281
rect 8857 -15341 11467 -15315
rect 8857 -15570 9017 -15341
rect 11307 -15570 11467 -15341
rect 8857 -15591 11467 -15570
rect 8857 -15625 9242 -15591
rect 9276 -15625 9500 -15591
rect 9534 -15625 9758 -15591
rect 9792 -15625 10016 -15591
rect 10050 -15625 10274 -15591
rect 10308 -15625 10532 -15591
rect 10566 -15625 10790 -15591
rect 10824 -15625 11048 -15591
rect 11082 -15625 11467 -15591
rect 8857 -15699 11467 -15625
rect 8857 -15733 9242 -15699
rect 9276 -15733 9500 -15699
rect 9534 -15733 9758 -15699
rect 9792 -15733 10016 -15699
rect 10050 -15733 10274 -15699
rect 10308 -15733 10532 -15699
rect 10566 -15733 10790 -15699
rect 10824 -15733 11048 -15699
rect 11082 -15733 11467 -15699
rect 8857 -15761 11467 -15733
rect 8040 -15985 8268 -15969
rect 8040 -16161 8070 -15985
rect 8232 -16161 8268 -15985
rect 8040 -20041 8268 -16161
rect 8857 -15980 9017 -15761
rect 11307 -15980 11467 -15761
rect 8857 -16009 11467 -15980
rect 8857 -16043 9242 -16009
rect 9276 -16043 9500 -16009
rect 9534 -16043 9758 -16009
rect 9792 -16043 10016 -16009
rect 10050 -16043 10274 -16009
rect 10308 -16043 10532 -16009
rect 10566 -16043 10790 -16009
rect 10824 -16043 11048 -16009
rect 11082 -16043 11467 -16009
rect 8857 -16117 11467 -16043
rect 8857 -16151 9242 -16117
rect 9276 -16151 9500 -16117
rect 9534 -16151 9758 -16117
rect 9792 -16151 10016 -16117
rect 10050 -16151 10274 -16117
rect 10308 -16151 10532 -16117
rect 10566 -16151 10790 -16117
rect 10824 -16151 11048 -16117
rect 11082 -16151 11467 -16117
rect 8857 -16171 11467 -16151
rect 8857 -16410 9017 -16171
rect 11307 -16410 11467 -16171
rect 8857 -16427 11467 -16410
rect 8857 -16461 9242 -16427
rect 9276 -16461 9500 -16427
rect 9534 -16461 9758 -16427
rect 9792 -16461 10016 -16427
rect 10050 -16461 10274 -16427
rect 10308 -16461 10532 -16427
rect 10566 -16461 10790 -16427
rect 10824 -16461 11048 -16427
rect 11082 -16461 11467 -16427
rect 8857 -16535 11467 -16461
rect 8857 -16569 9242 -16535
rect 9276 -16569 9500 -16535
rect 9534 -16569 9758 -16535
rect 9792 -16569 10016 -16535
rect 10050 -16569 10274 -16535
rect 10308 -16569 10532 -16535
rect 10566 -16569 10790 -16535
rect 10824 -16569 11048 -16535
rect 11082 -16569 11467 -16535
rect 8857 -16601 11467 -16569
rect 8857 -16820 9017 -16601
rect 11307 -16820 11467 -16601
rect 8857 -16845 11467 -16820
rect 8857 -16879 9242 -16845
rect 9276 -16879 9500 -16845
rect 9534 -16879 9758 -16845
rect 9792 -16879 10016 -16845
rect 10050 -16879 10274 -16845
rect 10308 -16879 10532 -16845
rect 10566 -16879 10790 -16845
rect 10824 -16879 11048 -16845
rect 11082 -16879 11467 -16845
rect 8857 -16953 11467 -16879
rect 8857 -16987 9242 -16953
rect 9276 -16987 9500 -16953
rect 9534 -16987 9758 -16953
rect 9792 -16987 10016 -16953
rect 10050 -16987 10274 -16953
rect 10308 -16987 10532 -16953
rect 10566 -16987 10790 -16953
rect 10824 -16987 11048 -16953
rect 11082 -16987 11467 -16953
rect 8857 -17011 11467 -16987
rect 8857 -17240 9017 -17011
rect 11307 -17240 11467 -17011
rect 8857 -17263 11467 -17240
rect 8857 -17297 9242 -17263
rect 9276 -17297 9500 -17263
rect 9534 -17297 9758 -17263
rect 9792 -17297 10016 -17263
rect 10050 -17297 10274 -17263
rect 10308 -17297 10532 -17263
rect 10566 -17297 10790 -17263
rect 10824 -17297 11048 -17263
rect 11082 -17297 11467 -17263
rect 8857 -17371 11467 -17297
rect 8857 -17405 9242 -17371
rect 9276 -17405 9500 -17371
rect 9534 -17405 9758 -17371
rect 9792 -17405 10016 -17371
rect 10050 -17405 10274 -17371
rect 10308 -17405 10532 -17371
rect 10566 -17405 10790 -17371
rect 10824 -17405 11048 -17371
rect 11082 -17405 11467 -17371
rect 8857 -17431 11467 -17405
rect 8857 -17650 9017 -17431
rect 11307 -17650 11467 -17431
rect 8857 -17681 11467 -17650
rect 8857 -17715 9242 -17681
rect 9276 -17715 9500 -17681
rect 9534 -17715 9758 -17681
rect 9792 -17715 10016 -17681
rect 10050 -17715 10274 -17681
rect 10308 -17715 10532 -17681
rect 10566 -17715 10790 -17681
rect 10824 -17715 11048 -17681
rect 11082 -17715 11467 -17681
rect 8857 -17789 11467 -17715
rect 8857 -17823 9242 -17789
rect 9276 -17823 9500 -17789
rect 9534 -17823 9758 -17789
rect 9792 -17823 10016 -17789
rect 10050 -17823 10274 -17789
rect 10308 -17823 10532 -17789
rect 10566 -17823 10790 -17789
rect 10824 -17823 11048 -17789
rect 11082 -17823 11467 -17789
rect 8857 -17841 11467 -17823
rect 8857 -18071 9017 -17841
rect 11307 -18071 11467 -17841
rect 8857 -18099 11467 -18071
rect 8857 -18133 9242 -18099
rect 9276 -18133 9500 -18099
rect 9534 -18133 9758 -18099
rect 9792 -18133 10016 -18099
rect 10050 -18133 10274 -18099
rect 10308 -18133 10532 -18099
rect 10566 -18133 10790 -18099
rect 10824 -18133 11048 -18099
rect 11082 -18133 11467 -18099
rect 8857 -18201 11467 -18133
rect 11527 -15242 11687 -15241
rect 12746 -15242 12872 -15205
rect 14190 -15241 14350 -15240
rect 15402 -15241 15528 -15181
rect 16640 -15241 16800 -15240
rect 13977 -15242 14137 -15241
rect 11527 -15281 14137 -15242
rect 11527 -15315 11912 -15281
rect 11946 -15315 12170 -15281
rect 12204 -15315 12428 -15281
rect 12462 -15315 12686 -15281
rect 12720 -15315 12944 -15281
rect 12978 -15315 13202 -15281
rect 13236 -15315 13460 -15281
rect 13494 -15315 13718 -15281
rect 13752 -15315 14137 -15281
rect 11527 -15341 14137 -15315
rect 11527 -15570 11687 -15341
rect 13977 -15570 14137 -15341
rect 11527 -15591 14137 -15570
rect 11527 -15625 11912 -15591
rect 11946 -15625 12170 -15591
rect 12204 -15625 12428 -15591
rect 12462 -15625 12686 -15591
rect 12720 -15625 12944 -15591
rect 12978 -15625 13202 -15591
rect 13236 -15625 13460 -15591
rect 13494 -15625 13718 -15591
rect 13752 -15625 14137 -15591
rect 11527 -15699 14137 -15625
rect 11527 -15733 11912 -15699
rect 11946 -15733 12170 -15699
rect 12204 -15733 12428 -15699
rect 12462 -15733 12686 -15699
rect 12720 -15733 12944 -15699
rect 12978 -15733 13202 -15699
rect 13236 -15733 13460 -15699
rect 13494 -15733 13718 -15699
rect 13752 -15733 14137 -15699
rect 11527 -15761 14137 -15733
rect 11527 -15980 11687 -15761
rect 13977 -15980 14137 -15761
rect 11527 -16009 14137 -15980
rect 11527 -16043 11912 -16009
rect 11946 -16043 12170 -16009
rect 12204 -16043 12428 -16009
rect 12462 -16043 12686 -16009
rect 12720 -16043 12944 -16009
rect 12978 -16043 13202 -16009
rect 13236 -16043 13460 -16009
rect 13494 -16043 13718 -16009
rect 13752 -16043 14137 -16009
rect 11527 -16117 14137 -16043
rect 11527 -16151 11912 -16117
rect 11946 -16151 12170 -16117
rect 12204 -16151 12428 -16117
rect 12462 -16151 12686 -16117
rect 12720 -16151 12944 -16117
rect 12978 -16151 13202 -16117
rect 13236 -16151 13460 -16117
rect 13494 -16151 13718 -16117
rect 13752 -16151 14137 -16117
rect 11527 -16171 14137 -16151
rect 11527 -16410 11687 -16171
rect 13977 -16410 14137 -16171
rect 11527 -16427 14137 -16410
rect 11527 -16461 11912 -16427
rect 11946 -16461 12170 -16427
rect 12204 -16461 12428 -16427
rect 12462 -16461 12686 -16427
rect 12720 -16461 12944 -16427
rect 12978 -16461 13202 -16427
rect 13236 -16461 13460 -16427
rect 13494 -16461 13718 -16427
rect 13752 -16461 14137 -16427
rect 11527 -16535 14137 -16461
rect 11527 -16569 11912 -16535
rect 11946 -16569 12170 -16535
rect 12204 -16569 12428 -16535
rect 12462 -16569 12686 -16535
rect 12720 -16569 12944 -16535
rect 12978 -16569 13202 -16535
rect 13236 -16569 13460 -16535
rect 13494 -16569 13718 -16535
rect 13752 -16569 14137 -16535
rect 11527 -16601 14137 -16569
rect 11527 -16820 11687 -16601
rect 13977 -16820 14137 -16601
rect 11527 -16845 14137 -16820
rect 11527 -16879 11912 -16845
rect 11946 -16879 12170 -16845
rect 12204 -16879 12428 -16845
rect 12462 -16879 12686 -16845
rect 12720 -16879 12944 -16845
rect 12978 -16879 13202 -16845
rect 13236 -16879 13460 -16845
rect 13494 -16879 13718 -16845
rect 13752 -16879 14137 -16845
rect 11527 -16953 14137 -16879
rect 11527 -16987 11912 -16953
rect 11946 -16987 12170 -16953
rect 12204 -16987 12428 -16953
rect 12462 -16987 12686 -16953
rect 12720 -16987 12944 -16953
rect 12978 -16987 13202 -16953
rect 13236 -16987 13460 -16953
rect 13494 -16987 13718 -16953
rect 13752 -16987 14137 -16953
rect 11527 -17011 14137 -16987
rect 11527 -17240 11687 -17011
rect 13977 -17240 14137 -17011
rect 11527 -17263 14137 -17240
rect 11527 -17297 11912 -17263
rect 11946 -17297 12170 -17263
rect 12204 -17297 12428 -17263
rect 12462 -17297 12686 -17263
rect 12720 -17297 12944 -17263
rect 12978 -17297 13202 -17263
rect 13236 -17297 13460 -17263
rect 13494 -17297 13718 -17263
rect 13752 -17297 14137 -17263
rect 11527 -17371 14137 -17297
rect 11527 -17405 11912 -17371
rect 11946 -17405 12170 -17371
rect 12204 -17405 12428 -17371
rect 12462 -17405 12686 -17371
rect 12720 -17405 12944 -17371
rect 12978 -17405 13202 -17371
rect 13236 -17405 13460 -17371
rect 13494 -17405 13718 -17371
rect 13752 -17405 14137 -17371
rect 11527 -17431 14137 -17405
rect 11527 -17650 11687 -17431
rect 13977 -17650 14137 -17431
rect 11527 -17681 14137 -17650
rect 11527 -17715 11912 -17681
rect 11946 -17715 12170 -17681
rect 12204 -17715 12428 -17681
rect 12462 -17715 12686 -17681
rect 12720 -17715 12944 -17681
rect 12978 -17715 13202 -17681
rect 13236 -17715 13460 -17681
rect 13494 -17715 13718 -17681
rect 13752 -17715 14137 -17681
rect 11527 -17789 14137 -17715
rect 11527 -17823 11912 -17789
rect 11946 -17823 12170 -17789
rect 12204 -17823 12428 -17789
rect 12462 -17823 12686 -17789
rect 12720 -17823 12944 -17789
rect 12978 -17823 13202 -17789
rect 13236 -17823 13460 -17789
rect 13494 -17823 13718 -17789
rect 13752 -17823 14137 -17789
rect 11527 -17841 14137 -17823
rect 11527 -18071 11687 -17841
rect 13977 -18071 14137 -17841
rect 11527 -18099 14137 -18071
rect 11527 -18133 11912 -18099
rect 11946 -18133 12170 -18099
rect 12204 -18133 12428 -18099
rect 12462 -18133 12686 -18099
rect 12720 -18133 12944 -18099
rect 12978 -18133 13202 -18099
rect 13236 -18133 13460 -18099
rect 13494 -18133 13718 -18099
rect 13752 -18133 14137 -18099
rect 11527 -18201 14137 -18133
rect 14190 -15280 16800 -15241
rect 14190 -15314 14575 -15280
rect 14609 -15314 14833 -15280
rect 14867 -15314 15091 -15280
rect 15125 -15314 15349 -15280
rect 15383 -15314 15607 -15280
rect 15641 -15314 15865 -15280
rect 15899 -15314 16123 -15280
rect 16157 -15314 16381 -15280
rect 16415 -15314 16800 -15280
rect 14190 -15340 16800 -15314
rect 14190 -15569 14350 -15340
rect 16640 -15569 16800 -15340
rect 14190 -15590 16800 -15569
rect 14190 -15624 14575 -15590
rect 14609 -15624 14833 -15590
rect 14867 -15624 15091 -15590
rect 15125 -15624 15349 -15590
rect 15383 -15624 15607 -15590
rect 15641 -15624 15865 -15590
rect 15899 -15624 16123 -15590
rect 16157 -15624 16381 -15590
rect 16415 -15624 16800 -15590
rect 14190 -15698 16800 -15624
rect 14190 -15732 14575 -15698
rect 14609 -15732 14833 -15698
rect 14867 -15732 15091 -15698
rect 15125 -15732 15349 -15698
rect 15383 -15732 15607 -15698
rect 15641 -15732 15865 -15698
rect 15899 -15732 16123 -15698
rect 16157 -15732 16381 -15698
rect 16415 -15732 16800 -15698
rect 14190 -15760 16800 -15732
rect 14190 -15979 14350 -15760
rect 16640 -15979 16800 -15760
rect 14190 -16008 16800 -15979
rect 14190 -16042 14575 -16008
rect 14609 -16042 14833 -16008
rect 14867 -16042 15091 -16008
rect 15125 -16042 15349 -16008
rect 15383 -16042 15607 -16008
rect 15641 -16042 15865 -16008
rect 15899 -16042 16123 -16008
rect 16157 -16042 16381 -16008
rect 16415 -16042 16800 -16008
rect 14190 -16116 16800 -16042
rect 14190 -16150 14575 -16116
rect 14609 -16150 14833 -16116
rect 14867 -16150 15091 -16116
rect 15125 -16150 15349 -16116
rect 15383 -16150 15607 -16116
rect 15641 -16150 15865 -16116
rect 15899 -16150 16123 -16116
rect 16157 -16150 16381 -16116
rect 16415 -16150 16800 -16116
rect 14190 -16170 16800 -16150
rect 14190 -16409 14350 -16170
rect 16640 -16409 16800 -16170
rect 14190 -16426 16800 -16409
rect 14190 -16460 14575 -16426
rect 14609 -16460 14833 -16426
rect 14867 -16460 15091 -16426
rect 15125 -16460 15349 -16426
rect 15383 -16460 15607 -16426
rect 15641 -16460 15865 -16426
rect 15899 -16460 16123 -16426
rect 16157 -16460 16381 -16426
rect 16415 -16460 16800 -16426
rect 14190 -16534 16800 -16460
rect 14190 -16568 14575 -16534
rect 14609 -16568 14833 -16534
rect 14867 -16568 15091 -16534
rect 15125 -16568 15349 -16534
rect 15383 -16568 15607 -16534
rect 15641 -16568 15865 -16534
rect 15899 -16568 16123 -16534
rect 16157 -16568 16381 -16534
rect 16415 -16568 16800 -16534
rect 14190 -16600 16800 -16568
rect 14190 -16819 14350 -16600
rect 16640 -16819 16800 -16600
rect 14190 -16844 16800 -16819
rect 14190 -16878 14575 -16844
rect 14609 -16878 14833 -16844
rect 14867 -16878 15091 -16844
rect 15125 -16878 15349 -16844
rect 15383 -16878 15607 -16844
rect 15641 -16878 15865 -16844
rect 15899 -16878 16123 -16844
rect 16157 -16878 16381 -16844
rect 16415 -16878 16800 -16844
rect 14190 -16952 16800 -16878
rect 14190 -16986 14575 -16952
rect 14609 -16986 14833 -16952
rect 14867 -16986 15091 -16952
rect 15125 -16986 15349 -16952
rect 15383 -16986 15607 -16952
rect 15641 -16986 15865 -16952
rect 15899 -16986 16123 -16952
rect 16157 -16986 16381 -16952
rect 16415 -16986 16800 -16952
rect 14190 -17010 16800 -16986
rect 14190 -17239 14350 -17010
rect 16640 -17239 16800 -17010
rect 14190 -17262 16800 -17239
rect 14190 -17296 14575 -17262
rect 14609 -17296 14833 -17262
rect 14867 -17296 15091 -17262
rect 15125 -17296 15349 -17262
rect 15383 -17296 15607 -17262
rect 15641 -17296 15865 -17262
rect 15899 -17296 16123 -17262
rect 16157 -17296 16381 -17262
rect 16415 -17296 16800 -17262
rect 14190 -17370 16800 -17296
rect 14190 -17404 14575 -17370
rect 14609 -17404 14833 -17370
rect 14867 -17404 15091 -17370
rect 15125 -17404 15349 -17370
rect 15383 -17404 15607 -17370
rect 15641 -17404 15865 -17370
rect 15899 -17404 16123 -17370
rect 16157 -17404 16381 -17370
rect 16415 -17404 16800 -17370
rect 14190 -17430 16800 -17404
rect 14190 -17649 14350 -17430
rect 16640 -17649 16800 -17430
rect 14190 -17680 16800 -17649
rect 14190 -17714 14575 -17680
rect 14609 -17714 14833 -17680
rect 14867 -17714 15091 -17680
rect 15125 -17714 15349 -17680
rect 15383 -17714 15607 -17680
rect 15641 -17714 15865 -17680
rect 15899 -17714 16123 -17680
rect 16157 -17714 16381 -17680
rect 16415 -17714 16800 -17680
rect 14190 -17788 16800 -17714
rect 14190 -17822 14575 -17788
rect 14609 -17822 14833 -17788
rect 14867 -17822 15091 -17788
rect 15125 -17822 15349 -17788
rect 15383 -17822 15607 -17788
rect 15641 -17822 15865 -17788
rect 15899 -17822 16123 -17788
rect 16157 -17822 16381 -17788
rect 16415 -17822 16800 -17788
rect 14190 -17840 16800 -17822
rect 14190 -18070 14350 -17840
rect 16640 -18070 16800 -17840
rect 14190 -18098 16800 -18070
rect 14190 -18132 14575 -18098
rect 14609 -18132 14833 -18098
rect 14867 -18132 15091 -18098
rect 15125 -18132 15349 -18098
rect 15383 -18132 15607 -18098
rect 15641 -18132 15865 -18098
rect 15899 -18132 16123 -18098
rect 16157 -18132 16381 -18098
rect 16415 -18132 16800 -18098
rect 14190 -18200 16800 -18132
rect 10107 -18441 10217 -18201
rect 10107 -18465 10137 -18441
rect 10106 -18481 10137 -18465
rect 10187 -18465 10217 -18441
rect 12777 -18441 12887 -18201
rect 12777 -18447 12807 -18441
rect 10187 -18481 10218 -18465
rect 10106 -18749 10218 -18481
rect 10106 -18787 10140 -18749
rect 10180 -18787 10218 -18749
rect 10106 -18821 10218 -18787
rect 12776 -18481 12807 -18447
rect 12857 -18447 12887 -18441
rect 15440 -18440 15550 -18200
rect 12857 -18481 12888 -18447
rect 12776 -18749 12888 -18481
rect 12776 -18787 12810 -18749
rect 12850 -18787 12888 -18749
rect 12776 -18809 12888 -18787
rect 15440 -18480 15470 -18440
rect 15520 -18480 15550 -18440
rect 15440 -18747 15550 -18480
rect 15440 -18789 15470 -18747
rect 15512 -18789 15550 -18747
rect 15440 -18803 15550 -18789
rect 9942 -18880 10096 -18870
rect 9942 -18986 9964 -18880
rect 10070 -18986 10096 -18880
rect 9942 -18997 10096 -18986
rect 12626 -18885 12751 -18869
rect 12626 -18979 12640 -18885
rect 12732 -18979 12751 -18885
rect 12626 -18991 12751 -18979
rect 15290 -18885 15415 -18865
rect 15290 -18979 15306 -18885
rect 15398 -18979 15415 -18885
rect 15290 -18991 15415 -18979
rect 16650 -19541 16772 -19513
rect 16206 -19577 16490 -19549
rect 16206 -19578 16247 -19577
rect 16449 -19578 16490 -19577
rect 16206 -19895 16242 -19578
rect 16458 -19895 16490 -19578
rect 16206 -19911 16490 -19895
rect 16650 -19575 16698 -19541
rect 16732 -19575 16772 -19541
rect 8040 -20217 8070 -20041
rect 8232 -20217 8268 -20041
rect 16650 -20005 16772 -19575
rect 17040 -19543 17184 -19515
rect 17040 -19577 17088 -19543
rect 17122 -19577 17184 -19543
rect 16870 -19747 16974 -19728
rect 16870 -19819 16887 -19747
rect 16958 -19819 16974 -19747
rect 16870 -19839 16974 -19819
rect 16650 -20039 16698 -20005
rect 16732 -20039 16772 -20005
rect 8040 -20251 8268 -20217
rect 8950 -20119 9137 -20102
rect 8950 -20391 8963 -20119
rect 9119 -20391 9137 -20119
rect 8950 -20419 9137 -20391
rect 10071 -20174 10197 -20166
rect 10071 -20235 10093 -20174
rect 10173 -20235 10197 -20174
rect 10071 -20395 10197 -20235
rect 10071 -20456 10094 -20395
rect 10174 -20456 10197 -20395
rect 10071 -20873 10197 -20456
rect 8040 -20889 10197 -20873
rect 8040 -21065 8070 -20889
rect 8232 -20916 10197 -20889
rect 12747 -20178 12873 -20165
rect 12747 -20261 12767 -20178
rect 12865 -20261 12873 -20178
rect 12747 -20373 12873 -20261
rect 12747 -20456 12767 -20373
rect 12865 -20456 12873 -20373
rect 12747 -20914 12873 -20456
rect 15403 -20178 15529 -20166
rect 15403 -20261 15419 -20178
rect 15517 -20261 15529 -20178
rect 15403 -20373 15529 -20261
rect 15403 -20456 15419 -20373
rect 15517 -20456 15529 -20373
rect 16650 -20337 16772 -20039
rect 17040 -20007 17184 -19577
rect 17040 -20041 17088 -20007
rect 17122 -20041 17184 -20007
rect 17040 -20169 17184 -20041
rect 16836 -20181 17184 -20169
rect 17365 -20171 17759 -20170
rect 16836 -20219 16848 -20181
rect 16902 -20219 17184 -20181
rect 16836 -20229 17184 -20219
rect 16836 -20231 16922 -20229
rect 16650 -20371 16702 -20337
rect 16736 -20371 16772 -20337
rect 15403 -20537 15529 -20456
rect 16500 -20415 16603 -20389
rect 16500 -20488 16523 -20415
rect 16579 -20488 16603 -20415
rect 16500 -20515 16603 -20488
rect 8232 -21065 10196 -20916
rect 12746 -20934 12873 -20914
rect 12746 -20976 12872 -20934
rect 8040 -21083 10196 -21065
rect 12743 -20987 12872 -20976
rect 12743 -21066 12755 -20987
rect 12850 -21066 12872 -20987
rect 12743 -21083 12872 -21066
rect 8856 -21146 9022 -21143
rect 10070 -21146 10196 -21083
rect 11307 -21146 11467 -21145
rect 8856 -21185 11467 -21146
rect 8856 -21219 9242 -21185
rect 9276 -21219 9500 -21185
rect 9534 -21219 9758 -21185
rect 9792 -21219 10016 -21185
rect 10050 -21219 10274 -21185
rect 10308 -21219 10532 -21185
rect 10566 -21219 10790 -21185
rect 10824 -21219 11048 -21185
rect 11082 -21219 11467 -21185
rect 8856 -21244 11467 -21219
rect 8857 -21245 11467 -21244
rect 8857 -21474 9017 -21245
rect 11307 -21474 11467 -21245
rect 8857 -21495 11467 -21474
rect 8857 -21529 9242 -21495
rect 9276 -21529 9500 -21495
rect 9534 -21529 9758 -21495
rect 9792 -21529 10016 -21495
rect 10050 -21529 10274 -21495
rect 10308 -21529 10532 -21495
rect 10566 -21529 10790 -21495
rect 10824 -21529 11048 -21495
rect 11082 -21529 11467 -21495
rect 8857 -21603 11467 -21529
rect 8857 -21637 9242 -21603
rect 9276 -21637 9500 -21603
rect 9534 -21637 9758 -21603
rect 9792 -21637 10016 -21603
rect 10050 -21637 10274 -21603
rect 10308 -21637 10532 -21603
rect 10566 -21637 10790 -21603
rect 10824 -21637 11048 -21603
rect 11082 -21637 11467 -21603
rect 8857 -21665 11467 -21637
rect 8857 -21884 9017 -21665
rect 11307 -21884 11467 -21665
rect 8857 -21913 11467 -21884
rect 8857 -21947 9242 -21913
rect 9276 -21947 9500 -21913
rect 9534 -21947 9758 -21913
rect 9792 -21947 10016 -21913
rect 10050 -21947 10274 -21913
rect 10308 -21947 10532 -21913
rect 10566 -21947 10790 -21913
rect 10824 -21947 11048 -21913
rect 11082 -21947 11467 -21913
rect 8857 -22021 11467 -21947
rect 8857 -22055 9242 -22021
rect 9276 -22055 9500 -22021
rect 9534 -22055 9758 -22021
rect 9792 -22055 10016 -22021
rect 10050 -22055 10274 -22021
rect 10308 -22055 10532 -22021
rect 10566 -22055 10790 -22021
rect 10824 -22055 11048 -22021
rect 11082 -22055 11467 -22021
rect 8857 -22075 11467 -22055
rect 8857 -22314 9017 -22075
rect 11307 -22314 11467 -22075
rect 8857 -22331 11467 -22314
rect 8857 -22365 9242 -22331
rect 9276 -22365 9500 -22331
rect 9534 -22365 9758 -22331
rect 9792 -22365 10016 -22331
rect 10050 -22365 10274 -22331
rect 10308 -22365 10532 -22331
rect 10566 -22365 10790 -22331
rect 10824 -22365 11048 -22331
rect 11082 -22365 11467 -22331
rect 8857 -22439 11467 -22365
rect 8857 -22473 9242 -22439
rect 9276 -22473 9500 -22439
rect 9534 -22473 9758 -22439
rect 9792 -22473 10016 -22439
rect 10050 -22473 10274 -22439
rect 10308 -22473 10532 -22439
rect 10566 -22473 10790 -22439
rect 10824 -22473 11048 -22439
rect 11082 -22473 11467 -22439
rect 8857 -22505 11467 -22473
rect 8857 -22724 9017 -22505
rect 11307 -22724 11467 -22505
rect 8857 -22749 11467 -22724
rect 8857 -22783 9242 -22749
rect 9276 -22783 9500 -22749
rect 9534 -22783 9758 -22749
rect 9792 -22783 10016 -22749
rect 10050 -22783 10274 -22749
rect 10308 -22783 10532 -22749
rect 10566 -22783 10790 -22749
rect 10824 -22783 11048 -22749
rect 11082 -22783 11467 -22749
rect 8857 -22857 11467 -22783
rect 8857 -22891 9242 -22857
rect 9276 -22891 9500 -22857
rect 9534 -22891 9758 -22857
rect 9792 -22891 10016 -22857
rect 10050 -22891 10274 -22857
rect 10308 -22891 10532 -22857
rect 10566 -22891 10790 -22857
rect 10824 -22891 11048 -22857
rect 11082 -22891 11467 -22857
rect 8857 -22915 11467 -22891
rect 8857 -23144 9017 -22915
rect 11307 -23144 11467 -22915
rect 8857 -23167 11467 -23144
rect 8857 -23201 9242 -23167
rect 9276 -23201 9500 -23167
rect 9534 -23201 9758 -23167
rect 9792 -23201 10016 -23167
rect 10050 -23201 10274 -23167
rect 10308 -23201 10532 -23167
rect 10566 -23201 10790 -23167
rect 10824 -23201 11048 -23167
rect 11082 -23201 11467 -23167
rect 8857 -23275 11467 -23201
rect 8857 -23309 9242 -23275
rect 9276 -23309 9500 -23275
rect 9534 -23309 9758 -23275
rect 9792 -23309 10016 -23275
rect 10050 -23309 10274 -23275
rect 10308 -23309 10532 -23275
rect 10566 -23309 10790 -23275
rect 10824 -23309 11048 -23275
rect 11082 -23309 11467 -23275
rect 8857 -23335 11467 -23309
rect 8857 -23554 9017 -23335
rect 11307 -23554 11467 -23335
rect 8857 -23585 11467 -23554
rect 8857 -23619 9242 -23585
rect 9276 -23619 9500 -23585
rect 9534 -23619 9758 -23585
rect 9792 -23619 10016 -23585
rect 10050 -23619 10274 -23585
rect 10308 -23619 10532 -23585
rect 10566 -23619 10790 -23585
rect 10824 -23619 11048 -23585
rect 11082 -23619 11467 -23585
rect 8857 -23693 11467 -23619
rect 8857 -23727 9242 -23693
rect 9276 -23727 9500 -23693
rect 9534 -23727 9758 -23693
rect 9792 -23727 10016 -23693
rect 10050 -23727 10274 -23693
rect 10308 -23727 10532 -23693
rect 10566 -23727 10790 -23693
rect 10824 -23727 11048 -23693
rect 11082 -23727 11467 -23693
rect 8857 -23745 11467 -23727
rect 8857 -23975 9017 -23745
rect 11307 -23975 11467 -23745
rect 8857 -24003 11467 -23975
rect 8857 -24037 9242 -24003
rect 9276 -24037 9500 -24003
rect 9534 -24037 9758 -24003
rect 9792 -24037 10016 -24003
rect 10050 -24037 10274 -24003
rect 10308 -24037 10532 -24003
rect 10566 -24037 10790 -24003
rect 10824 -24037 11048 -24003
rect 11082 -24037 11467 -24003
rect 8857 -24105 11467 -24037
rect 11527 -21146 11687 -21145
rect 12746 -21146 12872 -21083
rect 15402 -20940 15529 -20537
rect 16650 -20531 16772 -20371
rect 17040 -20337 17184 -20229
rect 17222 -20183 17759 -20171
rect 17222 -20227 17236 -20183
rect 17284 -20227 17759 -20183
rect 17222 -20235 17759 -20227
rect 17040 -20371 17092 -20337
rect 17126 -20371 17184 -20337
rect 16887 -20415 16990 -20387
rect 16887 -20488 16912 -20415
rect 16968 -20488 16990 -20415
rect 16887 -20513 16990 -20488
rect 16650 -20565 16702 -20531
rect 16736 -20565 16772 -20531
rect 16650 -20693 16772 -20565
rect 17040 -20531 17184 -20371
rect 17040 -20565 17092 -20531
rect 17126 -20565 17184 -20531
rect 17040 -20593 17184 -20565
rect 16498 -20741 17498 -20693
rect 15402 -20976 15528 -20940
rect 15402 -20987 15542 -20976
rect 15402 -21066 15428 -20987
rect 15523 -21066 15542 -20987
rect 15402 -21083 15542 -21066
rect 16498 -21031 16542 -20741
rect 16792 -20743 17498 -20741
rect 16792 -21031 17164 -20743
rect 16498 -21039 17164 -21031
rect 17416 -21039 17498 -20743
rect 14190 -21145 14350 -21144
rect 15402 -21145 15528 -21083
rect 16498 -21085 17498 -21039
rect 16640 -21145 16800 -21144
rect 13977 -21146 14137 -21145
rect 11527 -21185 14137 -21146
rect 11527 -21219 11912 -21185
rect 11946 -21219 12170 -21185
rect 12204 -21219 12428 -21185
rect 12462 -21219 12686 -21185
rect 12720 -21219 12944 -21185
rect 12978 -21219 13202 -21185
rect 13236 -21219 13460 -21185
rect 13494 -21219 13718 -21185
rect 13752 -21219 14137 -21185
rect 11527 -21245 14137 -21219
rect 11527 -21474 11687 -21245
rect 13977 -21474 14137 -21245
rect 11527 -21495 14137 -21474
rect 11527 -21529 11912 -21495
rect 11946 -21529 12170 -21495
rect 12204 -21529 12428 -21495
rect 12462 -21529 12686 -21495
rect 12720 -21529 12944 -21495
rect 12978 -21529 13202 -21495
rect 13236 -21529 13460 -21495
rect 13494 -21529 13718 -21495
rect 13752 -21529 14137 -21495
rect 11527 -21603 14137 -21529
rect 11527 -21637 11912 -21603
rect 11946 -21637 12170 -21603
rect 12204 -21637 12428 -21603
rect 12462 -21637 12686 -21603
rect 12720 -21637 12944 -21603
rect 12978 -21637 13202 -21603
rect 13236 -21637 13460 -21603
rect 13494 -21637 13718 -21603
rect 13752 -21637 14137 -21603
rect 11527 -21665 14137 -21637
rect 11527 -21884 11687 -21665
rect 13977 -21884 14137 -21665
rect 11527 -21913 14137 -21884
rect 11527 -21947 11912 -21913
rect 11946 -21947 12170 -21913
rect 12204 -21947 12428 -21913
rect 12462 -21947 12686 -21913
rect 12720 -21947 12944 -21913
rect 12978 -21947 13202 -21913
rect 13236 -21947 13460 -21913
rect 13494 -21947 13718 -21913
rect 13752 -21947 14137 -21913
rect 11527 -22021 14137 -21947
rect 11527 -22055 11912 -22021
rect 11946 -22055 12170 -22021
rect 12204 -22055 12428 -22021
rect 12462 -22055 12686 -22021
rect 12720 -22055 12944 -22021
rect 12978 -22055 13202 -22021
rect 13236 -22055 13460 -22021
rect 13494 -22055 13718 -22021
rect 13752 -22055 14137 -22021
rect 11527 -22075 14137 -22055
rect 11527 -22314 11687 -22075
rect 13977 -22314 14137 -22075
rect 11527 -22331 14137 -22314
rect 11527 -22365 11912 -22331
rect 11946 -22365 12170 -22331
rect 12204 -22365 12428 -22331
rect 12462 -22365 12686 -22331
rect 12720 -22365 12944 -22331
rect 12978 -22365 13202 -22331
rect 13236 -22365 13460 -22331
rect 13494 -22365 13718 -22331
rect 13752 -22365 14137 -22331
rect 11527 -22439 14137 -22365
rect 11527 -22473 11912 -22439
rect 11946 -22473 12170 -22439
rect 12204 -22473 12428 -22439
rect 12462 -22473 12686 -22439
rect 12720 -22473 12944 -22439
rect 12978 -22473 13202 -22439
rect 13236 -22473 13460 -22439
rect 13494 -22473 13718 -22439
rect 13752 -22473 14137 -22439
rect 11527 -22505 14137 -22473
rect 11527 -22724 11687 -22505
rect 13977 -22724 14137 -22505
rect 11527 -22749 14137 -22724
rect 11527 -22783 11912 -22749
rect 11946 -22783 12170 -22749
rect 12204 -22783 12428 -22749
rect 12462 -22783 12686 -22749
rect 12720 -22783 12944 -22749
rect 12978 -22783 13202 -22749
rect 13236 -22783 13460 -22749
rect 13494 -22783 13718 -22749
rect 13752 -22783 14137 -22749
rect 11527 -22857 14137 -22783
rect 11527 -22891 11912 -22857
rect 11946 -22891 12170 -22857
rect 12204 -22891 12428 -22857
rect 12462 -22891 12686 -22857
rect 12720 -22891 12944 -22857
rect 12978 -22891 13202 -22857
rect 13236 -22891 13460 -22857
rect 13494 -22891 13718 -22857
rect 13752 -22891 14137 -22857
rect 11527 -22915 14137 -22891
rect 11527 -23144 11687 -22915
rect 13977 -23144 14137 -22915
rect 11527 -23167 14137 -23144
rect 11527 -23201 11912 -23167
rect 11946 -23201 12170 -23167
rect 12204 -23201 12428 -23167
rect 12462 -23201 12686 -23167
rect 12720 -23201 12944 -23167
rect 12978 -23201 13202 -23167
rect 13236 -23201 13460 -23167
rect 13494 -23201 13718 -23167
rect 13752 -23201 14137 -23167
rect 11527 -23275 14137 -23201
rect 11527 -23309 11912 -23275
rect 11946 -23309 12170 -23275
rect 12204 -23309 12428 -23275
rect 12462 -23309 12686 -23275
rect 12720 -23309 12944 -23275
rect 12978 -23309 13202 -23275
rect 13236 -23309 13460 -23275
rect 13494 -23309 13718 -23275
rect 13752 -23309 14137 -23275
rect 11527 -23335 14137 -23309
rect 11527 -23554 11687 -23335
rect 13977 -23554 14137 -23335
rect 11527 -23585 14137 -23554
rect 11527 -23619 11912 -23585
rect 11946 -23619 12170 -23585
rect 12204 -23619 12428 -23585
rect 12462 -23619 12686 -23585
rect 12720 -23619 12944 -23585
rect 12978 -23619 13202 -23585
rect 13236 -23619 13460 -23585
rect 13494 -23619 13718 -23585
rect 13752 -23619 14137 -23585
rect 11527 -23693 14137 -23619
rect 11527 -23727 11912 -23693
rect 11946 -23727 12170 -23693
rect 12204 -23727 12428 -23693
rect 12462 -23727 12686 -23693
rect 12720 -23727 12944 -23693
rect 12978 -23727 13202 -23693
rect 13236 -23727 13460 -23693
rect 13494 -23727 13718 -23693
rect 13752 -23727 14137 -23693
rect 11527 -23745 14137 -23727
rect 11527 -23975 11687 -23745
rect 13977 -23975 14137 -23745
rect 11527 -24003 14137 -23975
rect 11527 -24037 11912 -24003
rect 11946 -24037 12170 -24003
rect 12204 -24037 12428 -24003
rect 12462 -24037 12686 -24003
rect 12720 -24037 12944 -24003
rect 12978 -24037 13202 -24003
rect 13236 -24037 13460 -24003
rect 13494 -24037 13718 -24003
rect 13752 -24037 14137 -24003
rect 11527 -24105 14137 -24037
rect 14190 -21184 16800 -21145
rect 14190 -21218 14575 -21184
rect 14609 -21218 14833 -21184
rect 14867 -21218 15091 -21184
rect 15125 -21218 15349 -21184
rect 15383 -21218 15607 -21184
rect 15641 -21218 15865 -21184
rect 15899 -21218 16123 -21184
rect 16157 -21218 16381 -21184
rect 16415 -21218 16800 -21184
rect 14190 -21244 16800 -21218
rect 14190 -21473 14350 -21244
rect 16640 -21473 16800 -21244
rect 14190 -21494 16800 -21473
rect 14190 -21528 14575 -21494
rect 14609 -21528 14833 -21494
rect 14867 -21528 15091 -21494
rect 15125 -21528 15349 -21494
rect 15383 -21528 15607 -21494
rect 15641 -21528 15865 -21494
rect 15899 -21528 16123 -21494
rect 16157 -21528 16381 -21494
rect 16415 -21528 16800 -21494
rect 14190 -21602 16800 -21528
rect 14190 -21636 14575 -21602
rect 14609 -21636 14833 -21602
rect 14867 -21636 15091 -21602
rect 15125 -21636 15349 -21602
rect 15383 -21636 15607 -21602
rect 15641 -21636 15865 -21602
rect 15899 -21636 16123 -21602
rect 16157 -21636 16381 -21602
rect 16415 -21636 16800 -21602
rect 14190 -21664 16800 -21636
rect 14190 -21883 14350 -21664
rect 16640 -21883 16800 -21664
rect 14190 -21912 16800 -21883
rect 14190 -21946 14575 -21912
rect 14609 -21946 14833 -21912
rect 14867 -21946 15091 -21912
rect 15125 -21946 15349 -21912
rect 15383 -21946 15607 -21912
rect 15641 -21946 15865 -21912
rect 15899 -21946 16123 -21912
rect 16157 -21946 16381 -21912
rect 16415 -21946 16800 -21912
rect 14190 -22020 16800 -21946
rect 14190 -22054 14575 -22020
rect 14609 -22054 14833 -22020
rect 14867 -22054 15091 -22020
rect 15125 -22054 15349 -22020
rect 15383 -22054 15607 -22020
rect 15641 -22054 15865 -22020
rect 15899 -22054 16123 -22020
rect 16157 -22054 16381 -22020
rect 16415 -22054 16800 -22020
rect 14190 -22074 16800 -22054
rect 14190 -22313 14350 -22074
rect 16640 -22313 16800 -22074
rect 14190 -22330 16800 -22313
rect 14190 -22364 14575 -22330
rect 14609 -22364 14833 -22330
rect 14867 -22364 15091 -22330
rect 15125 -22364 15349 -22330
rect 15383 -22364 15607 -22330
rect 15641 -22364 15865 -22330
rect 15899 -22364 16123 -22330
rect 16157 -22364 16381 -22330
rect 16415 -22364 16800 -22330
rect 14190 -22438 16800 -22364
rect 14190 -22472 14575 -22438
rect 14609 -22472 14833 -22438
rect 14867 -22472 15091 -22438
rect 15125 -22472 15349 -22438
rect 15383 -22472 15607 -22438
rect 15641 -22472 15865 -22438
rect 15899 -22472 16123 -22438
rect 16157 -22472 16381 -22438
rect 16415 -22472 16800 -22438
rect 14190 -22504 16800 -22472
rect 14190 -22723 14350 -22504
rect 16640 -22723 16800 -22504
rect 14190 -22748 16800 -22723
rect 14190 -22782 14575 -22748
rect 14609 -22782 14833 -22748
rect 14867 -22782 15091 -22748
rect 15125 -22782 15349 -22748
rect 15383 -22782 15607 -22748
rect 15641 -22782 15865 -22748
rect 15899 -22782 16123 -22748
rect 16157 -22782 16381 -22748
rect 16415 -22782 16800 -22748
rect 14190 -22856 16800 -22782
rect 14190 -22890 14575 -22856
rect 14609 -22890 14833 -22856
rect 14867 -22890 15091 -22856
rect 15125 -22890 15349 -22856
rect 15383 -22890 15607 -22856
rect 15641 -22890 15865 -22856
rect 15899 -22890 16123 -22856
rect 16157 -22890 16381 -22856
rect 16415 -22890 16800 -22856
rect 14190 -22914 16800 -22890
rect 14190 -23143 14350 -22914
rect 16640 -23143 16800 -22914
rect 14190 -23166 16800 -23143
rect 14190 -23200 14575 -23166
rect 14609 -23200 14833 -23166
rect 14867 -23200 15091 -23166
rect 15125 -23200 15349 -23166
rect 15383 -23200 15607 -23166
rect 15641 -23200 15865 -23166
rect 15899 -23200 16123 -23166
rect 16157 -23200 16381 -23166
rect 16415 -23200 16800 -23166
rect 14190 -23274 16800 -23200
rect 14190 -23308 14575 -23274
rect 14609 -23308 14833 -23274
rect 14867 -23308 15091 -23274
rect 15125 -23308 15349 -23274
rect 15383 -23308 15607 -23274
rect 15641 -23308 15865 -23274
rect 15899 -23308 16123 -23274
rect 16157 -23308 16381 -23274
rect 16415 -23308 16800 -23274
rect 14190 -23334 16800 -23308
rect 14190 -23553 14350 -23334
rect 16640 -23553 16800 -23334
rect 14190 -23584 16800 -23553
rect 14190 -23618 14575 -23584
rect 14609 -23618 14833 -23584
rect 14867 -23618 15091 -23584
rect 15125 -23618 15349 -23584
rect 15383 -23618 15607 -23584
rect 15641 -23618 15865 -23584
rect 15899 -23618 16123 -23584
rect 16157 -23618 16381 -23584
rect 16415 -23618 16800 -23584
rect 14190 -23692 16800 -23618
rect 14190 -23726 14575 -23692
rect 14609 -23726 14833 -23692
rect 14867 -23726 15091 -23692
rect 15125 -23726 15349 -23692
rect 15383 -23726 15607 -23692
rect 15641 -23726 15865 -23692
rect 15899 -23726 16123 -23692
rect 16157 -23726 16381 -23692
rect 16415 -23726 16800 -23692
rect 14190 -23744 16800 -23726
rect 14190 -23974 14350 -23744
rect 16640 -23974 16800 -23744
rect 14190 -24002 16800 -23974
rect 14190 -24036 14575 -24002
rect 14609 -24036 14833 -24002
rect 14867 -24036 15091 -24002
rect 15125 -24036 15349 -24002
rect 15383 -24036 15607 -24002
rect 15641 -24036 15865 -24002
rect 15899 -24036 16123 -24002
rect 16157 -24036 16381 -24002
rect 16415 -24036 16800 -24002
rect 14190 -24104 16800 -24036
rect 17122 -23033 17498 -23021
rect 17122 -23267 17202 -23033
rect 17426 -23267 17498 -23033
rect 10107 -24345 10217 -24105
rect 10107 -24371 10137 -24345
rect 10106 -24385 10137 -24371
rect 10187 -24385 10217 -24345
rect 10106 -24654 10217 -24385
rect 10106 -24690 10138 -24654
rect 10178 -24690 10217 -24654
rect 10106 -24709 10217 -24690
rect 12777 -24345 12887 -24105
rect 12777 -24385 12807 -24345
rect 12857 -24385 12887 -24345
rect 12777 -24651 12887 -24385
rect 12777 -24694 12808 -24651
rect 12852 -24694 12887 -24651
rect 12777 -24709 12887 -24694
rect 15440 -24344 15550 -24104
rect 15440 -24384 15470 -24344
rect 15520 -24384 15550 -24344
rect 15440 -24650 15550 -24384
rect 15440 -24692 15470 -24650
rect 15514 -24692 15550 -24650
rect 15440 -24716 15550 -24692
rect 9942 -24781 10096 -24760
rect 9942 -24875 9972 -24781
rect 10064 -24875 10096 -24781
rect 9942 -24887 10096 -24875
rect 12616 -24781 12763 -24765
rect 12616 -24875 12642 -24781
rect 12734 -24875 12763 -24781
rect 12616 -24888 12763 -24875
rect 15284 -24781 15431 -24767
rect 15284 -24875 15308 -24781
rect 15400 -24875 15431 -24781
rect 15284 -24890 15431 -24875
rect 7986 -25151 8490 -25029
rect 17122 -25151 17498 -23267
rect 7986 -25413 8086 -25151
rect 8380 -25253 17498 -25151
rect 8380 -25413 17496 -25253
rect 7986 -25457 17496 -25413
rect 7986 -25563 8490 -25457
rect 7833 -25814 7872 -25808
rect 4216 -25848 7872 -25814
rect 17834 -25764 17875 -7518
rect 17910 -7634 21419 -7518
rect 17910 -9010 17990 -7634
rect 18024 -9010 19648 -7634
rect 19682 -9010 21306 -7634
rect 21340 -9010 21419 -7634
rect 17910 -9144 21419 -9010
rect 17910 -10520 17990 -9144
rect 18024 -10520 19648 -9144
rect 19682 -10520 21306 -9144
rect 21340 -10520 21419 -9144
rect 17910 -10654 21419 -10520
rect 17910 -12030 17990 -10654
rect 18024 -12030 19648 -10654
rect 19682 -12030 21306 -10654
rect 21340 -12030 21419 -10654
rect 17910 -12164 21419 -12030
rect 17910 -13540 17990 -12164
rect 18024 -13391 19648 -12164
rect 19682 -13391 21306 -12164
rect 18024 -13540 19172 -13391
rect 20172 -13540 21306 -13391
rect 21340 -13540 21419 -12164
rect 17910 -13674 19172 -13540
rect 20172 -13674 21419 -13540
rect 17910 -15050 17990 -13674
rect 18024 -13987 19172 -13674
rect 20172 -13987 21306 -13674
rect 18024 -15050 19648 -13987
rect 19682 -15050 21306 -13987
rect 21340 -15050 21419 -13674
rect 17910 -15184 21419 -15050
rect 17910 -16560 17990 -15184
rect 18024 -16560 19648 -15184
rect 19682 -16560 21306 -15184
rect 21340 -16560 21419 -15184
rect 17910 -16694 21419 -16560
rect 17910 -18070 17990 -16694
rect 18024 -18070 19648 -16694
rect 19682 -18070 21306 -16694
rect 21340 -18070 21419 -16694
rect 17910 -18204 21419 -18070
rect 17910 -19580 17990 -18204
rect 18024 -19580 19648 -18204
rect 19682 -19580 21306 -18204
rect 21340 -19580 21419 -18204
rect 17910 -19714 21419 -19580
rect 17910 -21090 17990 -19714
rect 18024 -21090 19648 -19714
rect 19682 -21090 21306 -19714
rect 21340 -21090 21419 -19714
rect 17910 -21224 21419 -21090
rect 17910 -22600 17990 -21224
rect 18024 -22600 19648 -21224
rect 19682 -22600 21306 -21224
rect 21340 -22600 21419 -21224
rect 17910 -22734 21419 -22600
rect 17910 -24110 17990 -22734
rect 18024 -24110 19648 -22734
rect 19682 -24110 21306 -22734
rect 21340 -24110 21419 -22734
rect 17910 -24244 21419 -24110
rect 17910 -25620 17990 -24244
rect 18024 -25620 19648 -24244
rect 19682 -25620 21306 -24244
rect 21340 -25620 21419 -24244
rect 17910 -25764 21419 -25620
rect 21454 -25764 21491 -7518
rect 17834 -25809 17874 -25764
rect 21459 -25809 21491 -25764
rect 17834 -25844 21491 -25809
<< via1 >>
rect -18978 55462 -17592 56190
rect -14978 55462 -13592 56190
rect -10978 55462 -9592 56190
rect -6978 55462 -5592 56190
rect -2978 55462 -1592 56190
rect 1022 55462 2408 56190
rect 5022 55462 6408 56190
rect 9022 55462 10408 56190
rect 13022 55462 14408 56190
rect 17022 55462 18408 56190
rect 21022 55462 22408 56190
rect 25022 55462 26408 56190
rect 29022 55462 30408 56190
rect 33022 55462 34408 56190
rect 37022 55462 38408 56190
rect -20714 53298 -19328 54026
rect 37064 52260 38450 52988
rect -20714 49298 -19328 50026
rect -16260 49662 -16184 49684
rect -16260 49265 -16240 49662
rect -16240 49265 -16202 49662
rect -16202 49265 -16184 49662
rect -16260 49248 -16184 49265
rect -15940 49662 -15864 49684
rect -15940 49265 -15922 49662
rect -15922 49265 -15884 49662
rect -15884 49265 -15864 49662
rect -15940 49248 -15864 49265
rect -15624 49662 -15548 49684
rect -15624 49265 -15604 49662
rect -15604 49265 -15566 49662
rect -15566 49265 -15548 49662
rect -15624 49248 -15548 49265
rect -15304 49662 -15228 49684
rect -15304 49265 -15286 49662
rect -15286 49265 -15248 49662
rect -15248 49265 -15228 49662
rect -15304 49248 -15228 49265
rect 37064 48260 38450 48988
rect -20714 45298 -19328 46026
rect -16256 44505 -16184 44522
rect -16256 44108 -16240 44505
rect -16240 44108 -16202 44505
rect -16202 44108 -16184 44505
rect -16256 44090 -16184 44108
rect -15940 44505 -15868 44522
rect -15940 44108 -15922 44505
rect -15922 44108 -15884 44505
rect -15884 44108 -15868 44505
rect -15940 44090 -15868 44108
rect -15620 44505 -15548 44522
rect -15620 44108 -15604 44505
rect -15604 44108 -15566 44505
rect -15566 44108 -15548 44505
rect -15620 44090 -15548 44108
rect -15304 44505 -15232 44522
rect -15304 44108 -15286 44505
rect -15286 44108 -15248 44505
rect -15248 44108 -15232 44505
rect -15304 44090 -15232 44108
rect 37064 44260 38450 44988
rect -20714 41298 -19328 42026
rect -16204 42384 -16132 42400
rect -16204 41987 -16188 42384
rect -16188 41987 -16150 42384
rect -16150 41987 -16132 42384
rect -16204 41968 -16132 41987
rect -15134 42348 -15062 42372
rect -15134 41951 -15116 42348
rect -15116 41951 -15078 42348
rect -15078 41951 -15062 42348
rect -15134 41940 -15062 41951
rect 37064 40260 38450 40988
rect -20714 37298 -19328 38026
rect -16206 37227 -16132 37244
rect -16206 36830 -16188 37227
rect -16188 36830 -16150 37227
rect -16150 36830 -16132 37227
rect -16206 36812 -16132 36830
rect -15134 37191 -15060 37204
rect -15134 36794 -15116 37191
rect -15116 36794 -15078 37191
rect -15078 36794 -15060 37191
rect -15134 36772 -15060 36794
rect -20714 33298 -19328 34026
rect -20714 29298 -19328 30026
rect -20714 25298 -19328 26026
rect -16214 35884 -16140 35908
rect -16214 35487 -16196 35884
rect -16196 35487 -16158 35884
rect -16158 35487 -16140 35884
rect -16214 35476 -16140 35487
rect -13876 36162 -13688 36338
rect -11578 36390 -11378 36624
rect 37064 36260 38450 36988
rect -15190 35902 -15116 35918
rect -15190 35505 -15170 35902
rect -15170 35505 -15132 35902
rect -15132 35505 -15116 35902
rect -15190 35486 -15116 35505
rect 11372 34134 11636 34230
rect -16212 30727 -16142 30744
rect -16212 30330 -16196 30727
rect -16196 30330 -16158 30727
rect -16158 30330 -16142 30727
rect -16212 30310 -16142 30330
rect -15186 30745 -15116 30764
rect -15186 30348 -15170 30745
rect -15170 30348 -15132 30745
rect -15132 30348 -15116 30745
rect -15186 30330 -15116 30348
rect -16192 29132 -16120 29156
rect -16192 28735 -16174 29132
rect -16174 28735 -16136 29132
rect -16136 28735 -16120 29132
rect -16192 28718 -16120 28735
rect -15866 29132 -15794 29156
rect -15866 28735 -15856 29132
rect -15856 28735 -15818 29132
rect -15818 28735 -15794 29132
rect -15866 28718 -15794 28735
rect -15554 29132 -15482 29160
rect -15554 28735 -15538 29132
rect -15538 28735 -15500 29132
rect -15500 28735 -15482 29132
rect -15554 28722 -15482 28735
rect -15236 29132 -15164 29152
rect -15236 28735 -15220 29132
rect -15220 28735 -15182 29132
rect -15182 28735 -15164 29132
rect -15236 28714 -15164 28735
rect 9172 28064 9526 28258
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -96044 17274 -95512 17740
rect -96044 15274 -95512 15740
rect -96044 13274 -95512 13740
rect -96044 11274 -95512 11740
rect -96044 9274 -95512 9740
rect -96044 7274 -95512 7740
rect -96044 5274 -95512 5740
rect -20714 21298 -19328 22026
rect -27644 19274 -27112 19740
rect -16192 23975 -16120 23992
rect -16192 23578 -16174 23975
rect -16174 23578 -16136 23975
rect -16136 23578 -16120 23975
rect -16192 23554 -16120 23578
rect -15876 23975 -15804 23992
rect -15876 23578 -15856 23975
rect -15856 23578 -15818 23975
rect -15818 23578 -15804 23975
rect -15876 23554 -15804 23578
rect -15552 23975 -15480 23992
rect -15552 23578 -15538 23975
rect -15538 23578 -15500 23975
rect -15500 23578 -15480 23975
rect -15236 23975 -15164 23998
rect -15236 23590 -15220 23975
rect -15220 23590 -15182 23975
rect -15182 23590 -15164 23975
rect -15552 23554 -15480 23578
rect 37064 32260 38450 32988
rect 37064 28260 38450 28988
rect 37064 24260 38450 24988
rect 9218 20792 9482 21060
rect -27644 17274 -27112 17740
rect -20714 17298 -19328 18026
rect 16524 20618 16754 20860
rect 37064 20260 38450 20988
rect 13138 18134 13424 18404
rect 37064 16260 38450 16988
rect -27644 15274 -27112 15740
rect -18052 14180 -16666 14908
rect -14052 14180 -12666 14908
rect -10052 14180 -8666 14908
rect -6052 14180 -4666 14908
rect -2052 14180 -666 14908
rect 1948 14180 3334 14908
rect 5948 14180 7334 14908
rect 9948 14180 11334 14908
rect 13948 14180 15334 14908
rect 17948 14180 19334 14908
rect 21948 14180 23334 14908
rect 25948 14180 27334 14908
rect 29948 14180 31334 14908
rect 33948 14180 35334 14908
rect -27644 13274 -27112 13740
rect -27644 11274 -27112 11740
rect 18000 11574 18960 12068
rect -27644 9274 -27112 9740
rect -27644 7274 -27112 7740
rect 5368 10124 5800 10140
rect 5368 10086 5386 10124
rect 5386 10086 5783 10124
rect 5783 10086 5800 10124
rect 5368 10070 5800 10086
rect 9650 10124 10082 10140
rect 9650 10086 9667 10124
rect 9667 10086 10064 10124
rect 10064 10086 10082 10124
rect 9650 10070 10082 10086
rect 10564 10126 10998 10144
rect 10564 10088 10582 10126
rect 10582 10088 10979 10126
rect 10979 10088 10998 10126
rect 10564 10070 10998 10088
rect 5368 9806 5800 9822
rect 5368 9768 5386 9806
rect 5386 9768 5783 9806
rect 5783 9768 5800 9806
rect 5368 9752 5800 9768
rect 9650 9806 10082 9822
rect 9650 9768 9667 9806
rect 9667 9768 10064 9806
rect 10064 9768 10082 9806
rect 9650 9752 10082 9768
rect 5368 9488 5800 9504
rect 5368 9450 5386 9488
rect 5386 9450 5783 9488
rect 5783 9450 5800 9488
rect 5368 9434 5800 9450
rect 10564 9808 10998 9824
rect 10564 9770 10582 9808
rect 10582 9770 10979 9808
rect 10979 9770 10998 9808
rect 10564 9750 10998 9770
rect 14846 10126 15274 10142
rect 14846 10088 14863 10126
rect 14863 10088 15260 10126
rect 15260 10088 15274 10126
rect 14846 10072 15274 10088
rect 14848 9808 15276 9822
rect 14848 9770 14863 9808
rect 14863 9770 15260 9808
rect 15260 9770 15276 9808
rect 14848 9752 15276 9770
rect 9650 9488 10082 9504
rect 9650 9450 9667 9488
rect 9667 9450 10064 9488
rect 10064 9450 10082 9488
rect 9650 9434 10082 9450
rect 10562 9490 10996 9510
rect 10562 9452 10582 9490
rect 10582 9452 10979 9490
rect 10979 9452 10996 9490
rect 10562 9436 10996 9452
rect 14848 9490 15276 9506
rect 14848 9452 14863 9490
rect 14863 9452 15260 9490
rect 15260 9452 15276 9490
rect 14848 9436 15276 9452
rect 5368 9170 5802 9186
rect 5368 9132 5386 9170
rect 5386 9132 5783 9170
rect 5783 9132 5802 9170
rect 5368 9112 5802 9132
rect 5366 8852 5800 8870
rect 5366 8814 5386 8852
rect 5386 8814 5783 8852
rect 5783 8814 5800 8852
rect 5366 8796 5800 8814
rect 9650 9170 10082 9188
rect 9650 9132 9667 9170
rect 9667 9132 10064 9170
rect 10064 9132 10082 9170
rect 9650 9116 10082 9132
rect 9650 8852 10082 8870
rect 9650 8814 9667 8852
rect 9667 8814 10064 8852
rect 10064 8814 10082 8852
rect 9650 8798 10082 8814
rect 5368 8534 5800 8550
rect 5368 8496 5386 8534
rect 5386 8496 5783 8534
rect 5783 8496 5800 8534
rect 5368 8480 5800 8496
rect 10564 9172 10996 9188
rect 10564 9134 10582 9172
rect 10582 9134 10979 9172
rect 10979 9134 10996 9172
rect 10564 9118 10996 9134
rect 14846 9172 15278 9188
rect 14846 9134 14863 9172
rect 14863 9134 15260 9172
rect 15260 9134 15278 9172
rect 14846 9118 15278 9134
rect 10564 8854 10996 8870
rect 10564 8816 10582 8854
rect 10582 8816 10979 8854
rect 10979 8816 10996 8854
rect 10564 8800 10996 8816
rect 14846 8854 15278 8870
rect 14846 8816 14863 8854
rect 14863 8816 15260 8854
rect 15260 8816 15278 8854
rect 14846 8800 15278 8816
rect 9650 8534 10082 8552
rect 9650 8496 9667 8534
rect 9667 8496 10064 8534
rect 10064 8496 10082 8534
rect 9650 8478 10082 8496
rect 10564 8536 10996 8552
rect 10564 8498 10582 8536
rect 10582 8498 10979 8536
rect 10979 8498 10996 8536
rect 10564 8482 10996 8498
rect 14846 8536 15278 8552
rect 14846 8498 14863 8536
rect 14863 8498 15260 8536
rect 15260 8498 15278 8536
rect 14846 8482 15278 8498
rect 5368 8216 5794 8234
rect 5368 8178 5386 8216
rect 5386 8178 5783 8216
rect 5783 8178 5794 8216
rect 5368 8162 5794 8178
rect 5368 7898 5794 7916
rect 5368 7860 5386 7898
rect 5386 7860 5783 7898
rect 5783 7860 5794 7898
rect 5368 7844 5794 7860
rect 9650 8216 10082 8232
rect 9650 8178 9667 8216
rect 9667 8178 10064 8216
rect 10064 8178 10082 8216
rect 9650 8160 10082 8178
rect 10562 8218 11000 8236
rect 10562 8180 10582 8218
rect 10582 8180 10979 8218
rect 10979 8180 11000 8218
rect 10562 8162 11000 8180
rect 14846 8218 15278 8234
rect 14846 8180 14863 8218
rect 14863 8180 15260 8218
rect 15260 8180 15278 8218
rect 14846 8164 15278 8180
rect 9650 7898 10082 7916
rect 9650 7860 9667 7898
rect 9667 7860 10064 7898
rect 10064 7860 10082 7898
rect 9650 7844 10082 7860
rect 10562 7900 10998 7918
rect 10562 7862 10582 7900
rect 10582 7862 10979 7900
rect 10979 7862 10998 7900
rect 10562 7848 10998 7862
rect 5368 7580 5800 7598
rect 5368 7542 5386 7580
rect 5386 7542 5783 7580
rect 5783 7542 5800 7580
rect 5368 7526 5800 7542
rect 9652 7580 10080 7598
rect 9652 7542 9667 7580
rect 9667 7542 10064 7580
rect 10064 7542 10080 7580
rect 9652 7526 10080 7542
rect 10562 7582 10998 7598
rect 10562 7544 10582 7582
rect 10582 7544 10979 7582
rect 10979 7544 10998 7582
rect 10562 7528 10998 7544
rect 14846 7900 15282 7916
rect 14846 7862 14863 7900
rect 14863 7862 15260 7900
rect 15260 7862 15282 7900
rect 14846 7846 15282 7862
rect 14846 7582 15282 7598
rect 14846 7544 14863 7582
rect 14863 7544 15260 7582
rect 15260 7544 15282 7582
rect 14846 7528 15282 7544
rect 3932 6526 4052 6604
rect -27644 5274 -27112 5740
rect 1374 5776 1700 6016
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect -61788 3670 -61770 3722
rect -61770 3670 -61736 3722
rect -61370 3666 -61352 3718
rect -61352 3666 -61318 3718
rect -61844 3088 -61818 3184
rect -61818 3088 -61788 3184
rect -61426 3098 -61400 3184
rect -61400 3098 -61374 3184
rect 988 4816 1048 4880
rect 1386 4798 1394 4862
rect 1394 4798 1428 4862
rect 1428 4798 1450 4862
rect 1492 4904 1534 4974
rect 1534 4904 1568 4974
rect 1568 4904 1570 4974
rect 1616 4698 1622 4764
rect 1622 4698 1656 4764
rect 1656 4698 1688 4764
rect 1836 4912 1840 4978
rect 1840 4912 1874 4978
rect 1874 4912 1908 4978
rect 1068 4266 1098 4324
rect 1098 4266 1126 4324
rect 1844 4264 1876 4322
rect 1876 4264 1902 4322
rect 6262 5854 6588 6094
rect 6174 4834 6234 4898
rect 6572 4816 6580 4880
rect 6580 4816 6614 4880
rect 6614 4816 6636 4880
rect 6678 4922 6720 4992
rect 6720 4922 6754 4992
rect 6754 4922 6756 4992
rect 6802 4716 6808 4782
rect 6808 4716 6842 4782
rect 6842 4716 6874 4782
rect 7022 4930 7026 4996
rect 7026 4930 7060 4996
rect 7060 4930 7094 4996
rect 7630 6306 7682 6406
rect 7810 6318 7862 6402
rect 8534 6326 8612 6424
rect 10312 6320 10400 6452
rect 7918 6066 8094 6118
rect 7456 5936 7564 6022
rect 12778 6106 12860 6192
rect 14218 6120 14278 6174
rect 14794 6176 14856 6236
rect 11574 5642 11900 5882
rect 11350 4846 11410 4910
rect 6254 4284 6284 4342
rect 6284 4284 6312 4342
rect 7030 4282 7062 4340
rect 7062 4282 7088 4340
rect 7950 4408 8056 4462
rect 11748 4828 11756 4892
rect 11756 4828 11790 4892
rect 11790 4828 11812 4892
rect 11854 4934 11896 5004
rect 11896 4934 11930 5004
rect 11930 4934 11932 5004
rect 11978 4728 11984 4794
rect 11984 4728 12018 4794
rect 12018 4728 12050 4794
rect 12198 4942 12202 5008
rect 12202 4942 12236 5008
rect 12236 4942 12270 5008
rect 11430 4296 11460 4354
rect 11460 4296 11488 4354
rect 2210 3812 2286 3880
rect 12206 4294 12238 4352
rect 12238 4294 12264 4352
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect 10738 3716 10862 3768
rect -61864 2826 -61806 2878
rect -61464 2826 -61406 2878
rect 10728 2536 10846 2598
rect 17010 5584 17336 5824
rect 16664 5008 16746 5108
rect 17006 4638 17066 4702
rect 17404 4620 17412 4684
rect 17412 4620 17446 4684
rect 17446 4620 17468 4684
rect 17510 4726 17552 4796
rect 17552 4726 17586 4796
rect 17586 4726 17588 4796
rect 17634 4520 17640 4586
rect 17640 4520 17674 4586
rect 17674 4520 17706 4586
rect 17854 4734 17858 4800
rect 17858 4734 17892 4800
rect 17892 4734 17926 4800
rect 17086 4088 17116 4146
rect 17116 4088 17144 4146
rect 17862 4086 17894 4144
rect 17894 4086 17920 4144
rect 12876 3414 13064 3506
rect 12308 2096 12452 2228
rect 3524 1204 4484 1698
rect 10946 1020 11906 1514
rect 26138 3246 26538 3638
rect 26876 2794 26928 2796
rect 26876 2482 26886 2794
rect 26886 2482 26920 2794
rect 26920 2482 26928 2794
rect 26876 2478 26928 2482
rect 27082 2520 27090 2832
rect 27090 2520 27124 2832
rect 27124 2520 27134 2832
rect 26690 2190 26780 2264
rect 26874 2196 26936 2202
rect 26874 2072 26886 2196
rect 26886 2072 26920 2196
rect 26920 2072 26936 2196
rect 26874 2068 26936 2072
rect 27488 2802 27540 2804
rect 27488 2490 27498 2802
rect 27498 2490 27532 2802
rect 27532 2490 27540 2802
rect 27488 2486 27540 2490
rect 27694 2528 27702 2840
rect 27702 2528 27736 2840
rect 27736 2528 27746 2840
rect 27486 2204 27548 2210
rect 27486 2080 27498 2204
rect 27498 2080 27532 2204
rect 27532 2080 27548 2204
rect 27486 2076 27548 2080
rect 28066 2798 28118 2800
rect 28066 2486 28076 2798
rect 28076 2486 28110 2798
rect 28110 2486 28118 2798
rect 28066 2482 28118 2486
rect 28272 2524 28280 2836
rect 28280 2524 28314 2836
rect 28314 2524 28324 2836
rect 28064 2200 28126 2206
rect 28064 2076 28076 2200
rect 28076 2076 28110 2200
rect 28110 2076 28126 2200
rect 28064 2072 28126 2076
rect 28640 2806 28692 2808
rect 28640 2494 28650 2806
rect 28650 2494 28684 2806
rect 28684 2494 28692 2806
rect 28640 2490 28692 2494
rect 28846 2532 28854 2844
rect 28854 2532 28888 2844
rect 28888 2532 28898 2844
rect 28638 2208 28700 2214
rect 28638 2084 28650 2208
rect 28650 2084 28684 2208
rect 28684 2084 28700 2208
rect 28638 2080 28700 2084
rect 29218 2806 29270 2808
rect 29218 2494 29228 2806
rect 29228 2494 29262 2806
rect 29262 2494 29270 2806
rect 29218 2490 29270 2494
rect 29424 2532 29432 2844
rect 29432 2532 29466 2844
rect 29466 2532 29476 2844
rect 29216 2208 29278 2214
rect 29216 2084 29228 2208
rect 29228 2084 29262 2208
rect 29262 2084 29278 2208
rect 29216 2080 29278 2084
rect 29796 2806 29848 2808
rect 29796 2494 29806 2806
rect 29806 2494 29840 2806
rect 29840 2494 29848 2806
rect 29796 2490 29848 2494
rect 30002 2532 30010 2844
rect 30010 2532 30044 2844
rect 30044 2532 30054 2844
rect 29794 2208 29856 2214
rect 29794 2084 29806 2208
rect 29806 2084 29840 2208
rect 29840 2084 29856 2208
rect 29794 2080 29856 2084
rect 30378 2810 30430 2812
rect 30378 2498 30388 2810
rect 30388 2498 30422 2810
rect 30422 2498 30430 2810
rect 30378 2494 30430 2498
rect 30584 2536 30592 2848
rect 30592 2536 30626 2848
rect 30626 2536 30636 2848
rect 30376 2212 30438 2218
rect 30376 2088 30388 2212
rect 30388 2088 30422 2212
rect 30422 2088 30438 2212
rect 30376 2084 30438 2088
rect 30954 2806 31006 2808
rect 30954 2494 30964 2806
rect 30964 2494 30998 2806
rect 30998 2494 31006 2806
rect 30954 2490 31006 2494
rect 31160 2532 31168 2844
rect 31168 2532 31202 2844
rect 31202 2532 31212 2844
rect 30952 2208 31014 2214
rect 30952 2084 30964 2208
rect 30964 2084 30998 2208
rect 30998 2084 31014 2208
rect 30952 2080 31014 2084
rect 31524 2802 31576 2804
rect 31524 2490 31534 2802
rect 31534 2490 31568 2802
rect 31568 2490 31576 2802
rect 31524 2486 31576 2490
rect 31730 2528 31738 2840
rect 31738 2528 31772 2840
rect 31772 2528 31782 2840
rect 31522 2204 31584 2210
rect 31320 2012 31382 2074
rect 31522 2080 31534 2204
rect 31534 2080 31568 2204
rect 31568 2080 31584 2204
rect 31522 2076 31584 2080
rect 17578 1338 18538 1832
rect 32424 1746 32904 2206
rect 28270 428 28280 740
rect 28280 428 28314 740
rect 28314 428 28324 740
rect 28470 466 28480 778
rect 28480 466 28514 778
rect 28514 466 28524 778
rect 28270 -78 28280 234
rect 28280 -78 28314 234
rect 28314 -78 28324 234
rect 28470 -40 28480 272
rect 28480 -40 28514 272
rect 28514 -40 28524 272
rect 28672 426 28682 738
rect 28682 426 28716 738
rect 28716 426 28726 738
rect 28270 -586 28280 -274
rect 28280 -586 28314 -274
rect 28314 -586 28324 -274
rect 28470 -548 28480 -236
rect 28480 -548 28514 -236
rect 28514 -548 28524 -236
rect 28670 -78 28680 234
rect 28680 -78 28714 234
rect 28714 -78 28724 234
rect 28670 -586 28680 -274
rect 28680 -586 28714 -274
rect 28714 -586 28724 -274
rect 9031 -1196 9083 -1184
rect 9031 -1230 9039 -1196
rect 9039 -1230 9073 -1196
rect 9073 -1230 9083 -1196
rect 9031 -1236 9083 -1230
rect 11497 -1196 11549 -1183
rect 11497 -1230 11505 -1196
rect 11505 -1230 11539 -1196
rect 11539 -1230 11549 -1196
rect 11497 -1235 11549 -1230
rect 10478 -1266 10530 -1256
rect 10478 -1301 10488 -1266
rect 10488 -1301 10522 -1266
rect 10522 -1301 10530 -1266
rect 10478 -1308 10530 -1301
rect 10205 -1332 10257 -1325
rect 10205 -1366 10215 -1332
rect 10215 -1366 10249 -1332
rect 10249 -1366 10257 -1332
rect 10205 -1377 10257 -1366
rect 10775 -1265 10827 -1257
rect 10775 -1299 10783 -1265
rect 10783 -1299 10817 -1265
rect 10817 -1299 10827 -1265
rect 10775 -1309 10827 -1299
rect 11220 -1264 11272 -1254
rect 11220 -1298 11230 -1264
rect 11230 -1298 11264 -1264
rect 11264 -1298 11272 -1264
rect 11220 -1306 11272 -1298
rect 13244 -1264 13296 -1254
rect 13244 -1298 13251 -1264
rect 13251 -1298 13285 -1264
rect 13285 -1298 13296 -1264
rect 13244 -1306 13296 -1298
rect 12674 -1332 12726 -1327
rect 12674 -1366 12681 -1332
rect 12681 -1366 12715 -1332
rect 12715 -1366 12726 -1332
rect 12674 -1379 12726 -1366
rect 11221 -2032 11273 -2025
rect 11221 -2066 11230 -2032
rect 11230 -2066 11265 -2032
rect 11265 -2066 11273 -2032
rect 11221 -2077 11273 -2066
rect 10166 -2100 10181 -2086
rect 10181 -2100 10215 -2086
rect 10215 -2100 10218 -2086
rect 10166 -2138 10218 -2100
rect 10264 -2096 10316 -2088
rect 10264 -2130 10273 -2096
rect 10273 -2130 10307 -2096
rect 10307 -2130 10316 -2096
rect 10264 -2140 10316 -2130
rect 11500 -2028 11552 -2016
rect 11500 -2062 11505 -2028
rect 11505 -2062 11539 -2028
rect 11539 -2062 11552 -2028
rect 11500 -2068 11552 -2062
rect 12674 -2134 12726 -2128
rect 12674 -2168 12681 -2134
rect 12681 -2168 12715 -2134
rect 12715 -2168 12726 -2134
rect 12674 -2180 12726 -2168
rect 13242 -2097 13294 -2090
rect 13242 -2131 13249 -2097
rect 13249 -2131 13283 -2097
rect 13283 -2131 13294 -2097
rect 13242 -2142 13294 -2131
rect -7725 -4539 -7673 -4495
rect -7725 -4547 -7703 -4539
rect -7703 -4547 -7673 -4539
rect -8858 -4614 -8806 -4606
rect -8858 -4648 -8851 -4614
rect -8851 -4648 -8813 -4614
rect -8813 -4648 -8806 -4614
rect -8858 -4658 -8806 -4648
rect -7089 -4515 -7037 -4507
rect -7089 -4549 -7082 -4515
rect -7082 -4549 -7044 -4515
rect -7044 -4549 -7037 -4515
rect -7089 -4559 -7037 -4549
rect -5609 -4539 -5557 -4495
rect -5609 -4547 -5587 -4539
rect -5587 -4547 -5557 -4539
rect -6742 -4614 -6690 -4606
rect -6742 -4648 -6735 -4614
rect -6735 -4648 -6697 -4614
rect -6697 -4648 -6690 -4614
rect -6742 -4658 -6690 -4648
rect -4973 -4515 -4921 -4507
rect -4973 -4549 -4966 -4515
rect -4966 -4549 -4928 -4515
rect -4928 -4549 -4921 -4515
rect -4973 -4559 -4921 -4549
rect -3493 -4539 -3441 -4495
rect -3493 -4547 -3471 -4539
rect -3471 -4547 -3441 -4539
rect -4626 -4614 -4574 -4606
rect -4626 -4648 -4619 -4614
rect -4619 -4648 -4581 -4614
rect -4581 -4648 -4574 -4614
rect -4626 -4658 -4574 -4648
rect -2857 -4515 -2805 -4507
rect -2857 -4549 -2850 -4515
rect -2850 -4549 -2812 -4515
rect -2812 -4549 -2805 -4515
rect -2857 -4559 -2805 -4549
rect -1377 -4539 -1325 -4495
rect -1377 -4547 -1355 -4539
rect -1355 -4547 -1325 -4539
rect -2510 -4614 -2458 -4606
rect -2510 -4648 -2503 -4614
rect -2503 -4648 -2465 -4614
rect -2465 -4648 -2458 -4614
rect -2510 -4658 -2458 -4648
rect -741 -4515 -689 -4507
rect -741 -4549 -734 -4515
rect -734 -4549 -696 -4515
rect -696 -4549 -689 -4515
rect -741 -4559 -689 -4549
rect 739 -4539 791 -4495
rect 739 -4547 761 -4539
rect 761 -4547 791 -4539
rect -394 -4614 -342 -4606
rect -394 -4648 -387 -4614
rect -387 -4648 -349 -4614
rect -349 -4648 -342 -4614
rect -394 -4658 -342 -4648
rect 1375 -4515 1427 -4507
rect 1375 -4549 1382 -4515
rect 1382 -4549 1420 -4515
rect 1420 -4549 1427 -4515
rect 1375 -4559 1427 -4549
rect 2855 -4539 2907 -4495
rect 2855 -4547 2877 -4539
rect 2877 -4547 2907 -4539
rect 1722 -4614 1774 -4606
rect 1722 -4648 1729 -4614
rect 1729 -4648 1767 -4614
rect 1767 -4648 1774 -4614
rect 1722 -4658 1774 -4648
rect 3491 -4515 3543 -4507
rect 3491 -4549 3498 -4515
rect 3498 -4549 3536 -4515
rect 3536 -4549 3543 -4515
rect 3491 -4559 3543 -4549
rect 4971 -4539 5023 -4495
rect 4971 -4547 4993 -4539
rect 4993 -4547 5023 -4539
rect 3838 -4614 3890 -4606
rect 3838 -4648 3845 -4614
rect 3845 -4648 3883 -4614
rect 3883 -4648 3890 -4614
rect 3838 -4658 3890 -4648
rect 5607 -4515 5659 -4507
rect 5607 -4549 5614 -4515
rect 5614 -4549 5652 -4515
rect 5652 -4549 5659 -4515
rect 5607 -4559 5659 -4549
rect 7087 -4539 7139 -4495
rect 7087 -4547 7109 -4539
rect 7109 -4547 7139 -4539
rect 5954 -4614 6006 -4606
rect 5954 -4648 5961 -4614
rect 5961 -4648 5999 -4614
rect 5999 -4648 6006 -4614
rect 5954 -4658 6006 -4648
rect 7723 -4515 7775 -4507
rect 7723 -4549 7730 -4515
rect 7730 -4549 7768 -4515
rect 7768 -4549 7775 -4515
rect 7723 -4559 7775 -4549
rect 9203 -4539 9255 -4495
rect 9203 -4547 9225 -4539
rect 9225 -4547 9255 -4539
rect 8070 -4614 8122 -4606
rect 8070 -4648 8077 -4614
rect 8077 -4648 8115 -4614
rect 8115 -4648 8122 -4614
rect 8070 -4658 8122 -4648
rect 9839 -4515 9891 -4507
rect 9839 -4549 9846 -4515
rect 9846 -4549 9884 -4515
rect 9884 -4549 9891 -4515
rect 9839 -4559 9891 -4549
rect 11319 -4539 11371 -4495
rect 11319 -4547 11341 -4539
rect 11341 -4547 11371 -4539
rect 10186 -4614 10238 -4606
rect 10186 -4648 10193 -4614
rect 10193 -4648 10231 -4614
rect 10231 -4648 10238 -4614
rect 10186 -4658 10238 -4648
rect 11955 -4515 12007 -4507
rect 11955 -4549 11962 -4515
rect 11962 -4549 12000 -4515
rect 12000 -4549 12007 -4515
rect 11955 -4559 12007 -4549
rect 13435 -4539 13487 -4495
rect 13435 -4547 13457 -4539
rect 13457 -4547 13487 -4539
rect 12302 -4614 12354 -4606
rect 12302 -4648 12309 -4614
rect 12309 -4648 12347 -4614
rect 12347 -4648 12354 -4614
rect 12302 -4658 12354 -4648
rect 14071 -4515 14123 -4507
rect 14071 -4549 14078 -4515
rect 14078 -4549 14116 -4515
rect 14116 -4549 14123 -4515
rect 14071 -4559 14123 -4549
rect 15551 -4539 15603 -4495
rect 15551 -4547 15573 -4539
rect 15573 -4547 15603 -4539
rect 14418 -4614 14470 -4606
rect 14418 -4648 14425 -4614
rect 14425 -4648 14463 -4614
rect 14463 -4648 14470 -4614
rect 14418 -4658 14470 -4648
rect 16187 -4515 16239 -4507
rect 16187 -4549 16194 -4515
rect 16194 -4549 16232 -4515
rect 16232 -4549 16239 -4515
rect 16187 -4559 16239 -4549
rect 17667 -4539 17719 -4495
rect 17667 -4547 17689 -4539
rect 17689 -4547 17719 -4539
rect 16534 -4614 16586 -4606
rect 16534 -4648 16541 -4614
rect 16541 -4648 16579 -4614
rect 16579 -4648 16586 -4614
rect 16534 -4658 16586 -4648
rect 18303 -4515 18355 -4507
rect 18303 -4549 18310 -4515
rect 18310 -4549 18348 -4515
rect 18348 -4549 18355 -4515
rect 18303 -4559 18355 -4549
rect 19783 -4539 19835 -4495
rect 19783 -4547 19805 -4539
rect 19805 -4547 19835 -4539
rect 18650 -4614 18702 -4606
rect 18650 -4648 18657 -4614
rect 18657 -4648 18695 -4614
rect 18695 -4648 18702 -4614
rect 18650 -4658 18702 -4648
rect 20419 -4515 20471 -4507
rect 20419 -4549 20426 -4515
rect 20426 -4549 20464 -4515
rect 20464 -4549 20471 -4515
rect 20419 -4559 20471 -4549
rect 21899 -4539 21951 -4495
rect 21899 -4547 21921 -4539
rect 21921 -4547 21951 -4539
rect 20766 -4614 20818 -4606
rect 20766 -4648 20773 -4614
rect 20773 -4648 20811 -4614
rect 20811 -4648 20818 -4614
rect 20766 -4658 20818 -4648
rect 22535 -4515 22587 -4507
rect 22535 -4549 22542 -4515
rect 22542 -4549 22580 -4515
rect 22580 -4549 22587 -4515
rect 22535 -4559 22587 -4549
rect 24015 -4539 24067 -4495
rect 24015 -4547 24037 -4539
rect 24037 -4547 24067 -4539
rect 22882 -4614 22934 -4606
rect 22882 -4648 22889 -4614
rect 22889 -4648 22927 -4614
rect 22927 -4648 22934 -4614
rect 22882 -4658 22934 -4648
rect 24651 -4515 24703 -4507
rect 24651 -4549 24658 -4515
rect 24658 -4549 24696 -4515
rect 24696 -4549 24703 -4515
rect 24651 -4559 24703 -4549
rect 26131 -4539 26183 -4495
rect 26131 -4547 26153 -4539
rect 26153 -4547 26183 -4539
rect 24998 -4614 25050 -4606
rect 24998 -4648 25005 -4614
rect 25005 -4648 25043 -4614
rect 25043 -4648 25050 -4614
rect 24998 -4658 25050 -4648
rect 26767 -4515 26819 -4507
rect 26767 -4549 26774 -4515
rect 26774 -4549 26812 -4515
rect 26812 -4549 26819 -4515
rect 26767 -4559 26819 -4549
rect 28247 -4539 28299 -4495
rect 28247 -4547 28269 -4539
rect 28269 -4547 28299 -4539
rect 27114 -4614 27166 -4606
rect 27114 -4648 27121 -4614
rect 27121 -4648 27159 -4614
rect 27159 -4648 27166 -4614
rect 27114 -4658 27166 -4648
rect 28883 -4515 28935 -4507
rect 28883 -4549 28890 -4515
rect 28890 -4549 28928 -4515
rect 28928 -4549 28935 -4515
rect 28883 -4559 28935 -4549
rect 30363 -4539 30415 -4495
rect 30363 -4547 30385 -4539
rect 30385 -4547 30415 -4539
rect 29230 -4614 29282 -4606
rect 29230 -4648 29237 -4614
rect 29237 -4648 29275 -4614
rect 29275 -4648 29282 -4614
rect 29230 -4658 29282 -4648
rect 30999 -4515 31051 -4507
rect 30999 -4549 31006 -4515
rect 31006 -4549 31044 -4515
rect 31044 -4549 31051 -4515
rect 30999 -4559 31051 -4549
rect 32479 -4539 32531 -4495
rect 32479 -4547 32501 -4539
rect 32501 -4547 32531 -4539
rect 31346 -4614 31398 -4606
rect 31346 -4648 31353 -4614
rect 31353 -4648 31391 -4614
rect 31391 -4648 31398 -4614
rect 31346 -4658 31398 -4648
rect 33115 -4515 33167 -4507
rect 33115 -4549 33122 -4515
rect 33122 -4549 33160 -4515
rect 33160 -4549 33167 -4515
rect 33115 -4559 33167 -4549
rect 5413 -13467 6027 -12977
rect 6027 -13467 6061 -12977
rect 6061 -13467 6710 -12977
rect 9897 -7850 9960 -7689
rect 10023 -7849 10103 -7690
rect 10174 -7849 10254 -7690
rect 10286 -7848 10366 -7689
rect 12896 -7882 14455 -7656
rect 14341 -7884 14454 -7882
rect 9002 -8657 9241 -8654
rect 9002 -8959 9036 -8657
rect 9036 -8959 9209 -8657
rect 9209 -8959 9241 -8657
rect 9002 -8967 9241 -8959
rect 8042 -10831 8288 -10613
rect 16433 -8670 16655 -8669
rect 16433 -8989 16436 -8670
rect 16436 -8989 16651 -8670
rect 16651 -8989 16655 -8670
rect 16433 -8990 16655 -8989
rect 17324 -9429 17486 -9253
rect 17324 -10355 17486 -10179
rect 9970 -13267 10076 -13161
rect 12634 -13267 12740 -13161
rect 15296 -13267 15402 -13161
rect 8991 -14525 9174 -14220
rect 17324 -14237 17486 -14061
rect 8070 -15235 8232 -15059
rect 17324 -15163 17486 -14987
rect 8070 -16161 8232 -15985
rect 9964 -18986 10070 -18880
rect 12640 -18979 12732 -18885
rect 15306 -18979 15398 -18885
rect 16242 -19892 16247 -19578
rect 16247 -19892 16449 -19578
rect 16449 -19892 16458 -19578
rect 16242 -19895 16458 -19892
rect 8070 -20217 8232 -20041
rect 16887 -19819 16958 -19747
rect 8963 -20123 9119 -20119
rect 8963 -20387 8970 -20123
rect 8970 -20387 9113 -20123
rect 9113 -20387 9119 -20123
rect 8963 -20391 9119 -20387
rect 8070 -21065 8232 -20889
rect 16523 -20488 16579 -20415
rect 16912 -20488 16915 -20415
rect 16915 -20488 16961 -20415
rect 16961 -20488 16968 -20415
rect 17164 -21033 17414 -20743
rect 17414 -21033 17416 -20743
rect 17164 -21039 17416 -21033
rect 17202 -23267 17426 -23033
rect 9972 -24875 10064 -24781
rect 12642 -24875 12734 -24781
rect 15308 -24875 15400 -24781
rect 8086 -25413 8380 -25151
rect 19172 -13540 19648 -13391
rect 19648 -13540 19682 -13391
rect 19682 -13540 20172 -13391
rect 19172 -13674 20172 -13540
rect 19172 -13987 19648 -13674
rect 19648 -13987 19682 -13674
rect 19682 -13987 20172 -13674
<< metal2 >>
rect -19220 56190 -17382 56450
rect -19220 55462 -18978 56190
rect -17592 55462 -17382 56190
rect -19220 55220 -17382 55462
rect -15220 56190 -13382 56450
rect -15220 55462 -14978 56190
rect -13592 55462 -13382 56190
rect -15220 55220 -13382 55462
rect -11220 56190 -9382 56450
rect -11220 55462 -10978 56190
rect -9592 55462 -9382 56190
rect -11220 55220 -9382 55462
rect -7220 56190 -5382 56450
rect -7220 55462 -6978 56190
rect -5592 55462 -5382 56190
rect -7220 55220 -5382 55462
rect -3220 56190 -1382 56450
rect -3220 55462 -2978 56190
rect -1592 55462 -1382 56190
rect -3220 55220 -1382 55462
rect 780 56190 2618 56450
rect 780 55462 1022 56190
rect 2408 55462 2618 56190
rect 780 55220 2618 55462
rect 4780 56190 6618 56450
rect 4780 55462 5022 56190
rect 6408 55462 6618 56190
rect 4780 55220 6618 55462
rect 8780 56190 10618 56450
rect 8780 55462 9022 56190
rect 10408 55462 10618 56190
rect 8780 55220 10618 55462
rect 12780 56190 14618 56450
rect 12780 55462 13022 56190
rect 14408 55462 14618 56190
rect 12780 55220 14618 55462
rect 16780 56190 18618 56450
rect 16780 55462 17022 56190
rect 18408 55462 18618 56190
rect 16780 55220 18618 55462
rect 20780 56190 22618 56450
rect 20780 55462 21022 56190
rect 22408 55462 22618 56190
rect 20780 55220 22618 55462
rect 24780 56190 26618 56450
rect 24780 55462 25022 56190
rect 26408 55462 26618 56190
rect 24780 55220 26618 55462
rect 28780 56190 30618 56450
rect 28780 55462 29022 56190
rect 30408 55462 30618 56190
rect 28780 55220 30618 55462
rect 32780 56190 34618 56450
rect 32780 55462 33022 56190
rect 34408 55462 34618 56190
rect 32780 55220 34618 55462
rect 36780 56190 38618 56450
rect 36780 55462 37022 56190
rect 38408 55462 38618 56190
rect 36780 55220 38618 55462
rect -20956 54026 -19118 54286
rect -20956 53298 -20714 54026
rect -19328 53298 -19118 54026
rect -20956 53056 -19118 53298
rect -312 52964 23168 53816
rect 36822 52988 38660 53256
rect -312 52442 23260 52964
rect -20956 50026 -19118 50286
rect -20956 49298 -20714 50026
rect -19328 49298 -19118 50026
rect -20956 49056 -19118 49298
rect -16462 49684 -14894 49700
rect -16462 49248 -16260 49684
rect -16184 49248 -15940 49684
rect -15864 49248 -15624 49684
rect -15548 49248 -15304 49684
rect -15228 49248 -14894 49684
rect -20956 46026 -19118 46286
rect -20956 45298 -20714 46026
rect -19328 45298 -19118 46026
rect -20956 45056 -19118 45298
rect -16462 44522 -14894 49248
rect -16462 44090 -16256 44522
rect -16184 44090 -15940 44522
rect -15868 44090 -15620 44522
rect -15548 44090 -15304 44522
rect -15232 44090 -14894 44522
rect -16462 42400 -14894 44090
rect -20956 42026 -19118 42286
rect -20956 41298 -20714 42026
rect -19328 41298 -19118 42026
rect -20956 41056 -19118 41298
rect -16462 41968 -16204 42400
rect -16132 42372 -14894 42400
rect -260 44978 1042 52442
rect 21958 52102 23260 52442
rect 5844 51868 18096 52002
rect 5844 51076 16720 51868
rect 17836 51076 18096 51868
rect 5844 50944 18096 51076
rect 21958 51314 22192 52102
rect 23050 51314 23260 52102
rect 36822 52260 37064 52988
rect 38450 52260 38660 52988
rect 36822 52018 38660 52260
rect 5850 44996 7042 50944
rect -260 44958 1044 44978
rect -260 44886 388 44958
rect 550 44886 1044 44958
rect -260 43522 1044 44886
rect 5850 44924 6284 44996
rect 6446 44924 7042 44996
rect 5850 44884 7042 44924
rect 16662 45004 17854 50944
rect 16662 44932 17176 45004
rect 17338 44932 17854 45004
rect -260 42770 -14 43522
rect 668 42770 1044 43522
rect -260 42560 1044 42770
rect 5776 43194 7052 44884
rect 5776 42980 6278 43194
rect 6536 42980 7052 43194
rect -260 42382 1042 42560
rect 5776 42466 7052 42980
rect 16662 44052 17854 44932
rect 16662 42588 16860 44052
rect 17822 42588 17854 44052
rect -16132 41968 -15134 42372
rect -16462 41940 -15134 41968
rect -15062 41940 -14894 42372
rect 5850 42248 7042 42466
rect 16662 42202 17854 42588
rect 21958 44928 23260 51314
rect 36822 48988 38660 49256
rect 36822 48260 37064 48988
rect 38450 48260 38660 48988
rect 36822 48018 38660 48260
rect 21958 44856 22446 44928
rect 22608 44856 23260 44928
rect 21958 44304 23260 44856
rect 21958 42840 22142 44304
rect 23104 42840 23260 44304
rect 36822 44988 38660 45256
rect 36822 44260 37064 44988
rect 38450 44260 38660 44988
rect 36822 44018 38660 44260
rect 21958 42450 23260 42840
rect -20956 38026 -19118 38286
rect -20956 37298 -20714 38026
rect -19328 37298 -19118 38026
rect -20956 37056 -19118 37298
rect -16462 37244 -14894 41940
rect 36822 40988 38660 41256
rect 36822 40260 37064 40988
rect 38450 40260 38660 40988
rect 36822 40018 38660 40260
rect -16462 36812 -16206 37244
rect -16132 37204 -14894 37244
rect -16132 36812 -15134 37204
rect -16462 36772 -15134 36812
rect -15060 36772 -14894 37204
rect -16462 35918 -14894 36772
rect -244 38840 1176 39110
rect -244 37376 -54 38840
rect 908 37376 1176 38840
rect 13756 38836 16472 39012
rect 5476 38474 6124 38698
rect -11614 36624 -11334 36712
rect -13924 36338 -13646 36440
rect -13924 36162 -13876 36338
rect -13688 36162 -13646 36338
rect -11614 36390 -11578 36624
rect -11378 36390 -11334 36624
rect -11614 36314 -11334 36390
rect -13924 36074 -13646 36162
rect -16462 35908 -15190 35918
rect -16462 35476 -16214 35908
rect -16140 35486 -15190 35908
rect -15116 35486 -14894 35918
rect -16140 35476 -14894 35486
rect -20956 34026 -19118 34286
rect -20956 33298 -20714 34026
rect -19328 33298 -19118 34026
rect -20956 33056 -19118 33298
rect -16462 30764 -14894 35476
rect -16462 30744 -15186 30764
rect -16462 30310 -16212 30744
rect -16142 30330 -15186 30744
rect -15116 30330 -14894 30764
rect -16142 30310 -14894 30330
rect -20956 30026 -19118 30286
rect -20956 29298 -20714 30026
rect -19328 29298 -19118 30026
rect -20956 29056 -19118 29298
rect -16462 29160 -14894 30310
rect -16462 29156 -15554 29160
rect -16462 28718 -16192 29156
rect -16120 28718 -15866 29156
rect -15794 28722 -15554 29156
rect -15482 29152 -14894 29160
rect -15482 28722 -15236 29152
rect -15794 28718 -15236 28722
rect -16462 28714 -15236 28718
rect -15164 28714 -14894 29152
rect -20956 26026 -19118 26286
rect -20956 25298 -20714 26026
rect -19328 25298 -19118 26026
rect -20956 25056 -19118 25298
rect -16462 23998 -14894 28714
rect -244 34194 1176 37376
rect 5982 37010 6124 38474
rect 5476 35990 6124 37010
rect 13756 38566 17326 38836
rect 13756 37102 16472 38566
rect 17206 37102 17326 38566
rect 13756 36270 17326 37102
rect -244 34122 508 34194
rect 670 34122 1176 34194
rect -8390 27902 -6772 28176
rect -8390 27104 -8174 27902
rect -6984 27104 -6772 27902
rect -8390 26888 -6772 27104
rect -16462 23992 -15236 23998
rect -16462 23554 -16192 23992
rect -16120 23554 -15876 23992
rect -15804 23554 -15552 23992
rect -15480 23590 -15236 23992
rect -15164 23590 -14894 23998
rect -15480 23554 -14894 23590
rect -16462 22684 -14894 23554
rect -8264 23736 -8188 26888
rect -244 26256 1176 34122
rect 4910 34264 6124 35990
rect 4910 34192 5434 34264
rect 5596 34192 6124 34264
rect 4910 27450 6124 34192
rect 11324 34230 11700 34274
rect 11324 34134 11372 34230
rect 11636 34134 11700 34230
rect 11324 34106 11700 34134
rect 16112 34116 17326 36270
rect 16112 34044 16704 34116
rect 16866 34044 17326 34116
rect 8960 28258 9880 28336
rect 8960 28064 9172 28258
rect 9526 28064 9880 28258
rect 8960 28032 9880 28064
rect 16112 27450 17326 34044
rect 21702 38750 23122 39018
rect 21702 37286 21866 38750
rect 22828 37286 23122 38750
rect 21702 34204 23122 37286
rect 36822 36988 38660 37256
rect 36822 36260 37064 36988
rect 38450 36260 38660 36988
rect 36822 36018 38660 36260
rect 21702 34132 22228 34204
rect 22390 34132 23122 34204
rect -248 26050 1176 26256
rect -248 25118 20 26050
rect 728 25732 1176 26050
rect 4888 27028 17418 27450
rect 4888 25912 15928 27028
rect 17090 25912 17418 27028
rect 728 25118 1154 25732
rect 4888 25664 17418 25912
rect 21702 26142 23122 34132
rect 36822 32988 38660 33256
rect 36822 32260 37064 32988
rect 38450 32260 38660 32988
rect 36822 32018 38660 32260
rect 36822 28988 38660 29256
rect 36822 28260 37064 28988
rect 38450 28260 38660 28988
rect 36822 28018 38660 28260
rect 21702 25640 23154 26142
rect -248 24716 1154 25118
rect 21752 24716 23154 25640
rect 36822 24988 38660 25256
rect -20956 22026 -19118 22286
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -96266 13740 -95320 15274
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -96266 4182 -95320 5274
rect -27834 19740 -26806 21200
rect -20956 21298 -20714 22026
rect -19328 21298 -19118 22026
rect -20956 21056 -19118 21298
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -27834 17740 -26806 19274
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -27834 15740 -26806 17274
rect -20956 18026 -19118 18286
rect -20956 17298 -20714 18026
rect -19328 17298 -19118 18026
rect -20956 17056 -19118 17298
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -27834 13740 -26806 15274
rect -18294 14908 -16456 15184
rect -18294 14180 -18052 14908
rect -16666 14606 -16456 14908
rect -16314 14606 -16142 22684
rect -8264 21828 -8192 23736
rect -454 23404 23316 24716
rect 36822 24260 37064 24988
rect 38450 24260 38660 24988
rect 36822 24018 38660 24260
rect 21752 23336 23154 23404
rect -8264 21762 -8190 21828
rect -8262 20788 -8190 21762
rect 9136 21060 9548 21130
rect 9136 20792 9218 21060
rect 9482 20792 9548 21060
rect 36822 20988 38660 21256
rect -8262 20730 -8188 20788
rect -8260 19778 -8188 20730
rect 9136 20726 9548 20792
rect 16440 20860 16836 20964
rect 16440 20618 16524 20860
rect 16754 20618 16836 20860
rect 16440 20528 16836 20618
rect 36822 20260 37064 20988
rect 38450 20260 38660 20988
rect 36822 20018 38660 20260
rect -8260 19690 -8184 19778
rect -8256 16636 -8184 19690
rect 13066 18404 13490 18476
rect 13066 18134 13138 18404
rect 13424 18134 13490 18404
rect 13066 18052 13490 18134
rect -8258 16580 -8184 16636
rect 36822 16988 38660 17256
rect -8258 15610 -8186 16580
rect 36822 16260 37064 16988
rect 38450 16260 38660 16988
rect 36822 16018 38660 16260
rect -8258 15538 -8182 15610
rect -16666 14536 -16142 14606
rect -16666 14180 -16456 14536
rect -16314 14508 -16142 14536
rect -14294 15084 -14106 15180
rect -13566 15084 -12456 15180
rect -14294 14908 -12456 15084
rect -18294 13938 -16456 14180
rect -14294 14180 -14052 14908
rect -12666 14180 -12456 14908
rect -14294 13938 -12456 14180
rect -10294 14908 -8456 15180
rect -10294 14180 -10052 14908
rect -8666 14582 -8456 14908
rect -8254 14582 -8182 15538
rect -6294 14908 -4456 15180
rect -8666 14524 -8176 14582
rect -8666 14180 -8456 14524
rect -8254 14512 -8182 14524
rect -10294 13938 -8456 14180
rect -6294 14180 -6052 14908
rect -4666 14180 -4456 14908
rect -6294 13938 -4456 14180
rect -2294 14908 -456 15180
rect -2294 14180 -2052 14908
rect -666 14180 -456 14908
rect -2294 13938 -456 14180
rect 1706 14908 3544 15180
rect 1706 14180 1948 14908
rect 3334 14180 3544 14908
rect 1706 13938 3544 14180
rect 5706 14908 7544 15180
rect 5706 14180 5948 14908
rect 7334 14180 7544 14908
rect 5706 13938 7544 14180
rect 9706 14908 11544 15180
rect 9706 14180 9948 14908
rect 11334 14180 11544 14908
rect 9706 13938 11544 14180
rect 13706 14908 15544 15180
rect 13706 14180 13948 14908
rect 15334 14180 15544 14908
rect 13706 13938 15544 14180
rect 17706 14908 19544 15180
rect 17706 14180 17948 14908
rect 19334 14180 19544 14908
rect 17706 13938 19544 14180
rect 21706 14908 23544 15180
rect 21706 14180 21948 14908
rect 23334 14180 23544 14908
rect 21706 13938 23544 14180
rect 25706 14908 27544 15180
rect 25706 14180 25948 14908
rect 27334 14180 27544 14908
rect 25706 13938 27544 14180
rect 29706 14908 31544 15180
rect 29706 14180 29948 14908
rect 31334 14180 31544 14908
rect 29706 13938 31544 14180
rect 33706 14908 35544 15180
rect 33706 14180 33948 14908
rect 35334 14180 35544 14908
rect 33706 13938 35544 14180
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -27834 11740 -26806 13274
rect 17792 12068 19104 12262
rect 9300 11810 9356 11820
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect 9296 11804 14830 11810
rect 17792 11804 18000 12068
rect 9296 11718 18000 11804
rect -27834 9740 -26806 11274
rect 5354 10140 5804 10154
rect 5354 10070 5368 10140
rect 5800 10070 5804 10140
rect 5354 9822 5804 10070
rect 5354 9752 5368 9822
rect 5800 9752 5804 9822
rect 5354 9742 5804 9752
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect 5356 9508 5810 9524
rect 5356 9434 5368 9508
rect 5800 9434 5810 9508
rect 5356 9418 5810 9434
rect -27834 7740 -26806 9274
rect 5356 9188 5816 9202
rect 5356 9112 5368 9188
rect 5800 9186 5816 9188
rect 5802 9112 5816 9186
rect 5356 8870 5816 9112
rect 5356 8796 5366 8870
rect 5356 8794 5368 8796
rect 5802 8794 5816 8870
rect 5356 8782 5816 8794
rect 5360 8556 5808 8560
rect 3940 8550 5808 8556
rect 3940 8480 5368 8550
rect 5800 8480 5808 8550
rect 3940 8468 5808 8480
rect 3940 8466 5546 8468
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -27834 5740 -26806 7274
rect 3966 8288 4022 8466
rect 3966 6634 4018 8288
rect 5354 8236 5804 8244
rect 5354 8234 5806 8236
rect 5354 8162 5368 8234
rect 5794 8162 5806 8234
rect 5354 7998 5806 8162
rect 9300 8062 9356 11718
rect 14486 11686 18000 11718
rect 9862 10222 13710 10260
rect 9862 10158 9912 10222
rect 9644 10140 10098 10158
rect 9644 10070 9650 10140
rect 10082 10070 10098 10140
rect 9644 10052 10098 10070
rect 10552 10144 11002 10154
rect 10552 10070 10564 10144
rect 10998 10070 11002 10144
rect 9642 9822 10098 9836
rect 9642 9752 9650 9822
rect 10082 9752 10098 9822
rect 9642 9504 10098 9752
rect 10552 9824 11002 10070
rect 10552 9750 10564 9824
rect 10998 9750 11002 9824
rect 10552 9738 11002 9750
rect 9642 9434 9650 9504
rect 10082 9434 10098 9504
rect 9642 9420 10098 9434
rect 10552 9510 11006 9520
rect 10552 9436 10562 9510
rect 10996 9436 11006 9510
rect 10552 9426 11006 9436
rect 10738 9332 10784 9426
rect 10738 9294 12820 9332
rect 9636 9188 10092 9206
rect 9636 9116 9650 9188
rect 10082 9116 10092 9188
rect 9636 8870 10092 9116
rect 9636 8798 9650 8870
rect 10082 8798 10092 8870
rect 9636 8552 10092 8798
rect 10554 9188 11000 9200
rect 10554 9118 10564 9188
rect 10996 9118 11000 9188
rect 10554 8870 11000 9118
rect 10554 8800 10564 8870
rect 10996 8800 11000 8870
rect 10554 8788 11000 8800
rect 9636 8478 9650 8552
rect 10082 8478 10092 8552
rect 9636 8466 10092 8478
rect 10554 8552 11002 8562
rect 10554 8482 10564 8552
rect 10996 8482 11002 8552
rect 10554 8472 11002 8482
rect 10770 8412 10836 8472
rect 12128 8412 12200 8418
rect 10770 8350 12200 8412
rect 10770 8348 10836 8350
rect 9646 8232 10092 8250
rect 9646 8160 9650 8232
rect 10082 8160 10092 8232
rect 9646 8062 10092 8160
rect 10556 8236 11010 8246
rect 10556 8162 10562 8236
rect 11000 8162 11010 8236
rect 10556 8152 11010 8162
rect 7640 7998 7676 8004
rect 9300 8002 10092 8062
rect 10818 8074 10856 8152
rect 10818 8026 11706 8074
rect 5354 7956 7676 7998
rect 5354 7916 5806 7956
rect 5354 7844 5368 7916
rect 5794 7844 5806 7916
rect 5354 7842 5806 7844
rect 5354 7832 5804 7842
rect 5360 7600 5808 7610
rect 5118 7598 5808 7600
rect 5118 7544 5368 7598
rect 5118 6654 5166 7544
rect 5360 7526 5368 7544
rect 5800 7526 5808 7598
rect 5360 7516 5808 7526
rect 3910 6604 4078 6634
rect 3910 6526 3932 6604
rect 4052 6526 4078 6604
rect 3910 6492 4078 6526
rect 5112 6188 5172 6654
rect 7640 6426 7676 7956
rect 9646 7916 10092 8002
rect 9646 7844 9650 7916
rect 10082 7844 10092 7916
rect 9646 7832 10092 7844
rect 10552 7918 11006 7934
rect 10552 7848 10562 7918
rect 10998 7848 11006 7918
rect 10552 7734 11006 7848
rect 7806 7682 11006 7734
rect 7806 7680 7982 7682
rect 7806 6426 7870 7680
rect 9646 7598 10094 7608
rect 9646 7526 9652 7598
rect 10080 7526 10094 7598
rect 9646 7514 10094 7526
rect 10552 7598 11006 7682
rect 10552 7528 10562 7598
rect 10998 7528 11006 7598
rect 9794 7480 9850 7514
rect 10552 7508 11006 7528
rect 8530 7444 9850 7480
rect 8530 7440 9834 7444
rect 8530 6444 8586 7440
rect 10298 6452 10416 6478
rect 7618 6406 7694 6426
rect 7618 6306 7630 6406
rect 7682 6306 7694 6406
rect 7618 6286 7694 6306
rect 7794 6402 7880 6426
rect 7794 6318 7810 6402
rect 7862 6318 7880 6402
rect 7794 6294 7880 6318
rect 8522 6424 8622 6444
rect 8522 6326 8534 6424
rect 8612 6326 8622 6424
rect 8522 6294 8622 6326
rect 10298 6320 10312 6452
rect 10400 6438 10416 6452
rect 11640 6438 11706 8026
rect 10400 6378 11706 6438
rect 10400 6372 11702 6378
rect 10400 6320 10416 6372
rect 10298 6300 10416 6320
rect 6168 6188 6682 6190
rect 5112 6154 6682 6188
rect 5114 6150 6682 6154
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 1280 5776 1374 6016
rect 1700 5776 1794 6016
rect 1280 5678 1794 5776
rect 6168 6094 6682 6150
rect 7894 6118 8126 6142
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 7694 6108 7766 6110
rect 7894 6108 7918 6118
rect 7694 6068 7918 6108
rect 7440 6022 7580 6040
rect 7440 5936 7456 6022
rect 7564 5936 7580 6022
rect 7440 5916 7580 5936
rect 6168 5756 6682 5854
rect 7460 5608 7564 5916
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -96396 3740 -62544 3910
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -61816 3722 -61296 3892
rect -27834 3846 -26806 5274
rect 984 5556 7564 5608
rect 984 5040 1058 5556
rect 7694 5410 7766 6068
rect 7894 6066 7918 6068
rect 8094 6066 8126 6118
rect 7894 6046 8126 6066
rect 11480 5882 11994 5978
rect 11480 5642 11574 5882
rect 11900 5766 11994 5882
rect 12128 5766 12200 8350
rect 12778 6204 12820 9294
rect 12764 6192 12872 6204
rect 12764 6106 12778 6192
rect 12860 6106 12872 6192
rect 13670 6166 13710 10222
rect 14486 7740 14546 11686
rect 17792 11574 18000 11686
rect 18960 11574 19104 12068
rect 17792 11354 19104 11574
rect 14834 10142 15292 10154
rect 14834 10072 14846 10142
rect 15274 10072 15292 10142
rect 14834 9822 15292 10072
rect 14834 9752 14848 9822
rect 15276 9752 15292 9822
rect 14834 9652 15292 9752
rect 14834 9600 15294 9652
rect 14834 9506 15292 9600
rect 14834 9436 14848 9506
rect 15276 9436 15292 9506
rect 14834 9416 15292 9436
rect 15416 9200 15494 9202
rect 15144 9198 15494 9200
rect 14842 9188 15494 9198
rect 14842 9118 14846 9188
rect 15278 9118 15494 9188
rect 14842 9108 15494 9118
rect 15144 9104 15494 9108
rect 14842 8870 15288 8882
rect 14842 8800 14846 8870
rect 15278 8800 15288 8870
rect 14842 8552 15288 8800
rect 14842 8482 14846 8552
rect 15278 8482 15288 8552
rect 14842 8470 15288 8482
rect 14836 8234 15290 8246
rect 14836 8164 14846 8234
rect 15278 8164 15290 8234
rect 14836 8152 15290 8164
rect 14838 7916 15294 7930
rect 14838 7846 14846 7916
rect 15282 7846 15294 7916
rect 14838 7740 15294 7846
rect 14486 7662 15294 7740
rect 14838 7598 15294 7662
rect 14838 7528 14846 7598
rect 15282 7528 15294 7598
rect 14838 7512 15294 7528
rect 15416 6280 15494 9104
rect 14776 6236 14874 6254
rect 14196 6174 14294 6180
rect 14196 6166 14218 6174
rect 13670 6120 14218 6166
rect 14278 6120 14294 6174
rect 14776 6176 14794 6236
rect 14856 6214 14874 6236
rect 15414 6214 15496 6280
rect 14856 6192 15496 6214
rect 14856 6186 15494 6192
rect 14856 6176 14874 6186
rect 14776 6158 14874 6176
rect 13670 6118 14294 6120
rect 12764 6088 12872 6106
rect 14196 6104 14294 6118
rect 16916 5824 17430 5920
rect 11900 5690 12202 5766
rect 11900 5642 11994 5690
rect 12128 5684 12200 5690
rect 11480 5544 11994 5642
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect 2064 5354 7766 5410
rect 1192 5040 1246 5042
rect 970 5034 1246 5040
rect 1386 5036 1456 5040
rect 1384 5034 1456 5036
rect 970 4880 1456 5034
rect 1484 4978 1912 5040
rect 2064 4978 2140 5354
rect 7694 5352 7766 5354
rect 16638 5108 16776 5134
rect 11554 5070 11608 5072
rect 11332 5064 11608 5070
rect 11748 5066 11818 5070
rect 11746 5064 11818 5066
rect 6378 5058 6432 5060
rect 1484 4974 1836 4978
rect 1484 4904 1492 4974
rect 1570 4912 1836 4974
rect 1908 4912 2140 4978
rect 1570 4910 2140 4912
rect 1570 4904 1912 4910
rect 2064 4906 2140 4910
rect 6156 5052 6432 5058
rect 6572 5054 6642 5058
rect 6570 5052 6642 5054
rect 1484 4886 1912 4904
rect 1494 4884 1912 4886
rect 6156 4898 6642 5052
rect 6670 4996 7098 5058
rect 6670 4992 7022 4996
rect 6670 4922 6678 4992
rect 6756 4930 7022 4992
rect 7094 4930 7098 4996
rect 6756 4922 7098 4930
rect 6670 4904 7098 4922
rect 6680 4902 7098 4904
rect 11332 4910 11818 5064
rect 11846 5008 12274 5070
rect 11846 5004 12198 5008
rect 11846 4934 11854 5004
rect 11932 4942 12198 5004
rect 12270 4942 12274 5008
rect 16638 5008 16664 5108
rect 16746 5008 16776 5108
rect 16638 4978 16776 5008
rect 11932 4934 12274 4942
rect 11846 4916 12274 4934
rect 11856 4914 12274 4916
rect 11890 4910 12244 4914
rect 6714 4898 7068 4902
rect 1528 4880 1882 4884
rect 970 4816 988 4880
rect 1048 4862 1456 4880
rect 1048 4816 1386 4862
rect 970 4798 1386 4816
rect 1450 4798 1456 4862
rect 970 4640 1456 4798
rect 6156 4834 6174 4898
rect 6234 4880 6642 4898
rect 6234 4834 6572 4880
rect 6156 4816 6572 4834
rect 6636 4816 6642 4880
rect 2014 4774 2068 4780
rect 1606 4764 2068 4774
rect 1606 4698 1616 4764
rect 1688 4698 2068 4764
rect 1606 4688 2068 4698
rect 970 4638 1210 4640
rect 1242 4638 1456 4640
rect 1384 4636 1456 4638
rect 1050 4324 1912 4402
rect 1050 4266 1068 4324
rect 1126 4322 1912 4324
rect 1126 4266 1844 4322
rect 1050 4264 1844 4266
rect 1902 4264 1912 4322
rect 1050 4200 1912 4264
rect 2014 3866 2068 4688
rect 6156 4658 6642 4816
rect 11332 4846 11350 4910
rect 11410 4892 11818 4910
rect 11410 4846 11748 4892
rect 11332 4828 11748 4846
rect 11812 4828 11818 4892
rect 17210 4862 17264 4864
rect 6792 4782 7252 4792
rect 6792 4716 6802 4782
rect 6874 4772 7252 4782
rect 7700 4772 7746 4776
rect 6874 4732 7746 4772
rect 6874 4716 7252 4732
rect 6792 4706 7252 4716
rect 6156 4656 6396 4658
rect 6428 4656 6642 4658
rect 6570 4654 6642 4656
rect 7700 4454 7746 4732
rect 11332 4670 11818 4828
rect 16988 4856 17264 4862
rect 17404 4858 17474 4862
rect 17402 4856 17474 4858
rect 12374 4804 12432 4806
rect 11968 4794 12432 4804
rect 11968 4728 11978 4794
rect 12050 4728 12432 4794
rect 11968 4718 12432 4728
rect 11332 4668 11572 4670
rect 11604 4668 11818 4670
rect 11746 4666 11818 4668
rect 7924 4462 8082 4474
rect 7924 4454 7950 4462
rect 7700 4420 7950 4454
rect 6236 4342 7098 4420
rect 7702 4414 7950 4420
rect 7924 4408 7950 4414
rect 8056 4408 8082 4462
rect 7924 4394 8082 4408
rect 6236 4284 6254 4342
rect 6312 4340 7098 4342
rect 6312 4284 7030 4340
rect 6236 4282 7030 4284
rect 7088 4282 7098 4340
rect 6236 4218 7098 4282
rect 11412 4354 12274 4432
rect 11412 4296 11430 4354
rect 11488 4352 12274 4354
rect 11488 4296 12206 4352
rect 11412 4294 12206 4296
rect 12264 4294 12274 4352
rect 11412 4230 12274 4294
rect 12374 4044 12432 4718
rect 16988 4702 17474 4856
rect 17502 4800 17930 4862
rect 17502 4796 17854 4800
rect 17502 4726 17510 4796
rect 17588 4734 17854 4796
rect 17926 4734 17930 4800
rect 17588 4726 17930 4734
rect 17502 4708 17930 4726
rect 17512 4706 17930 4708
rect 17546 4702 17900 4706
rect 16988 4638 17006 4702
rect 17066 4684 17474 4702
rect 17066 4638 17404 4684
rect 16988 4620 17404 4638
rect 17468 4620 17474 4684
rect 16988 4462 17474 4620
rect 17624 4586 18084 4596
rect 17624 4520 17634 4586
rect 17706 4520 18084 4586
rect 17624 4510 18084 4520
rect 16988 4460 17228 4462
rect 17260 4460 17474 4462
rect 17402 4458 17474 4460
rect 17068 4146 17930 4224
rect 17068 4088 17086 4146
rect 17144 4144 17930 4146
rect 17144 4088 17862 4144
rect 17068 4086 17862 4088
rect 17920 4086 17930 4144
rect 2190 3880 2310 3902
rect 2190 3866 2210 3880
rect -61816 3670 -61788 3722
rect -61736 3718 -61296 3722
rect -61736 3670 -61370 3718
rect -61816 3666 -61370 3670
rect -61318 3666 -61296 3718
rect -61816 3490 -61296 3666
rect -60278 3740 -26756 3846
rect 2014 3824 2210 3866
rect 2016 3816 2210 3824
rect 2190 3812 2210 3816
rect 2286 3812 2310 3880
rect 2190 3786 2310 3812
rect -96396 2966 -62544 3274
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect 10712 3772 10888 3786
rect 10712 3716 10738 3772
rect 10862 3716 10888 3772
rect 10712 3698 10888 3716
rect 12376 3476 12428 4044
rect 17068 4022 17930 4086
rect 16228 3804 16448 3842
rect 16228 3686 16256 3804
rect 16414 3766 16448 3804
rect 18030 3766 18082 4510
rect 16414 3698 18084 3766
rect 16414 3686 16448 3698
rect 16228 3656 16448 3686
rect 26112 3638 26592 3676
rect 12850 3506 13108 3516
rect 12850 3476 12876 3506
rect 12374 3422 12876 3476
rect -61858 3184 -61358 3244
rect -60278 3224 -26756 3274
rect -61858 3088 -61844 3184
rect -61788 3098 -61426 3184
rect -61374 3098 -61358 3184
rect -61788 3088 -61358 3098
rect -61858 3046 -61358 3088
rect -61896 2882 -61292 2894
rect -61896 2826 -61864 2882
rect -61806 2826 -61464 2882
rect -61406 2826 -61292 2882
rect -61896 2812 -61292 2826
rect 10714 2598 10860 2608
rect 10714 2536 10728 2598
rect 10846 2536 10860 2598
rect 10714 2524 10860 2536
rect 12376 2270 12428 3422
rect 12850 3414 12876 3422
rect 13064 3414 13108 3506
rect 12850 3402 13108 3414
rect 26112 3246 26138 3638
rect 26538 3272 26592 3638
rect 26538 3246 26600 3272
rect 26112 3242 26600 3246
rect 26112 3216 26474 3242
rect 26206 3174 26474 3216
rect 26208 3164 26474 3174
rect 26802 3164 31696 3176
rect 26208 3094 31696 3164
rect 26874 2806 26932 3094
rect 27078 2832 27136 2844
rect 26872 2796 26934 2806
rect 26872 2478 26876 2796
rect 26928 2558 26934 2796
rect 27078 2558 27082 2832
rect 26928 2520 27082 2558
rect 27134 2520 27136 2832
rect 26928 2518 27136 2520
rect 26928 2478 26934 2518
rect 27078 2508 27136 2518
rect 27484 2804 27546 3094
rect 26872 2470 26934 2478
rect 27484 2486 27488 2804
rect 27540 2566 27546 2804
rect 27690 2840 27748 2852
rect 27690 2566 27694 2840
rect 27540 2528 27694 2566
rect 27746 2528 27748 2840
rect 28064 2810 28122 3094
rect 28268 2836 28326 2848
rect 27540 2526 27748 2528
rect 27540 2486 27546 2526
rect 27690 2516 27748 2526
rect 28062 2800 28124 2810
rect 27484 2476 27546 2486
rect 28062 2482 28066 2800
rect 28118 2562 28124 2800
rect 28268 2562 28272 2836
rect 28118 2524 28272 2562
rect 28324 2524 28326 2836
rect 28118 2522 28326 2524
rect 28118 2482 28124 2522
rect 28268 2512 28326 2522
rect 28632 2808 28700 3094
rect 28062 2474 28124 2482
rect 28632 2490 28640 2808
rect 28692 2570 28700 2808
rect 28842 2844 28900 2856
rect 28842 2570 28846 2844
rect 28692 2532 28846 2570
rect 28898 2532 28900 2844
rect 28692 2530 28900 2532
rect 28692 2490 28700 2530
rect 28842 2520 28900 2530
rect 29212 2808 29276 3094
rect 28632 2478 28700 2490
rect 29212 2490 29218 2808
rect 29270 2570 29276 2808
rect 29420 2844 29478 2856
rect 29420 2570 29424 2844
rect 29270 2532 29424 2570
rect 29476 2532 29478 2844
rect 29270 2530 29478 2532
rect 29270 2490 29276 2530
rect 29420 2520 29478 2530
rect 29788 2818 29850 3094
rect 29998 2844 30056 2856
rect 29788 2808 29854 2818
rect 29212 2482 29276 2490
rect 29788 2490 29796 2808
rect 29848 2570 29854 2808
rect 29998 2570 30002 2844
rect 29848 2532 30002 2570
rect 30054 2532 30056 2844
rect 29848 2530 30056 2532
rect 29848 2490 29854 2530
rect 29998 2520 30056 2530
rect 30368 2822 30430 3094
rect 30580 2848 30638 2860
rect 30368 2812 30436 2822
rect 29788 2482 29854 2490
rect 30368 2494 30378 2812
rect 30430 2574 30436 2812
rect 30580 2574 30584 2848
rect 30430 2536 30584 2574
rect 30636 2536 30638 2848
rect 30430 2534 30638 2536
rect 30430 2494 30436 2534
rect 30580 2524 30638 2534
rect 30950 2818 31006 3094
rect 31156 2844 31214 2856
rect 30950 2808 31012 2818
rect 30368 2486 30436 2494
rect 30950 2490 30954 2808
rect 31006 2570 31012 2808
rect 31156 2570 31160 2844
rect 31006 2532 31160 2570
rect 31212 2532 31214 2844
rect 31006 2530 31214 2532
rect 31006 2490 31012 2530
rect 31156 2520 31214 2530
rect 31520 2804 31582 3094
rect 29788 2474 29850 2482
rect 30368 2480 30430 2486
rect 30950 2482 31012 2490
rect 31520 2486 31524 2804
rect 31576 2566 31582 2804
rect 31726 2840 31784 2852
rect 31726 2566 31730 2840
rect 31576 2528 31730 2566
rect 31782 2528 31784 2840
rect 31576 2526 31784 2528
rect 31576 2486 31582 2526
rect 31726 2516 31784 2526
rect 30950 2474 31006 2482
rect 31520 2476 31582 2486
rect 26874 2468 26932 2470
rect 12272 2228 12500 2270
rect 12272 2096 12308 2228
rect 12452 2096 12500 2228
rect 26678 2264 26796 2280
rect 26678 2190 26690 2264
rect 26780 2190 26796 2264
rect 30376 2224 30436 2226
rect 29794 2220 29854 2222
rect 26876 2210 26936 2212
rect 26678 2176 26796 2190
rect 26872 2202 26936 2210
rect 12272 2064 12500 2096
rect 26872 2068 26874 2202
rect 3316 1698 4628 1892
rect 17370 1832 18682 2026
rect 26872 1950 26936 2068
rect 27486 2210 27548 2216
rect 28636 2214 28700 2220
rect 27486 2068 27548 2076
rect 28064 2206 28126 2214
rect 27486 1950 27546 2068
rect 28064 2058 28126 2072
rect 28636 2080 28638 2214
rect 28636 2072 28700 2080
rect 29216 2214 29278 2220
rect 28636 2070 28698 2072
rect 28064 1950 28124 2058
rect 28636 1950 28696 2070
rect 29216 2062 29278 2080
rect 29218 1950 29278 2062
rect 29794 2214 29856 2220
rect 29794 2072 29856 2080
rect 30376 2218 30438 2224
rect 30376 2076 30438 2084
rect 30952 2214 31014 2220
rect 31534 2216 31582 2218
rect 31522 2210 31584 2216
rect 29794 1950 29854 2072
rect 30376 1950 30436 2076
rect 30952 2068 31014 2080
rect 30954 1950 31014 2068
rect 31306 2074 31396 2090
rect 31306 2012 31320 2074
rect 31382 2012 31396 2074
rect 31306 1998 31396 2012
rect 31522 2068 31584 2076
rect 32364 2206 32976 2274
rect 26872 1948 31298 1950
rect 31522 1948 31582 2068
rect 32364 2064 32424 2206
rect 31830 1970 32424 2064
rect 31830 1948 31902 1970
rect 26872 1898 31902 1948
rect 31296 1896 31902 1898
rect 31830 1894 31902 1896
rect 3316 1204 3524 1698
rect 4484 1204 4628 1698
rect 3316 984 4628 1204
rect 10738 1514 12050 1708
rect 10738 1020 10946 1514
rect 11906 1020 12050 1514
rect 17370 1338 17578 1832
rect 18538 1338 18682 1832
rect 32364 1746 32424 1970
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 17370 1118 18682 1338
rect 10738 800 12050 1020
rect 28468 778 28528 790
rect 28266 740 28326 754
rect 28266 428 28270 740
rect 28324 708 28326 740
rect 28468 708 28470 778
rect 28324 654 28470 708
rect 28324 428 28326 654
rect 28266 234 28326 428
rect 28266 -78 28270 234
rect 28324 28 28326 234
rect 28468 466 28470 654
rect 28524 708 28528 778
rect 28668 738 28728 750
rect 28668 708 28672 738
rect 28524 654 28672 708
rect 28524 466 28528 654
rect 28468 272 28528 466
rect 28468 28 28470 272
rect 28324 -26 28470 28
rect 28324 -78 28326 -26
rect 28266 -274 28326 -78
rect 28266 -416 28270 -274
rect 28262 -470 28270 -416
rect 28266 -586 28270 -470
rect 28324 -416 28326 -274
rect 28468 -40 28470 -26
rect 28524 28 28528 272
rect 28668 426 28672 654
rect 28726 708 28728 738
rect 28726 654 28730 708
rect 28726 426 28728 654
rect 28668 234 28728 426
rect 28668 28 28670 234
rect 28524 -26 28670 28
rect 28524 -40 28528 -26
rect 28468 -236 28528 -40
rect 28468 -414 28470 -236
rect 28466 -416 28470 -414
rect 28324 -470 28470 -416
rect 28324 -586 28326 -470
rect 28468 -548 28470 -470
rect 28524 -414 28528 -236
rect 28668 -78 28670 -26
rect 28724 -78 28728 234
rect 28668 -274 28728 -78
rect 28668 -414 28670 -274
rect 28524 -468 28670 -414
rect 28524 -548 28528 -468
rect 28468 -560 28528 -548
rect 28266 -602 28326 -586
rect 28668 -586 28670 -468
rect 28724 -586 28728 -274
rect 28668 -600 28728 -586
rect 9025 -847 10957 -804
rect 13408 -805 13447 -804
rect 9025 -859 10890 -847
rect 9025 -1184 9089 -859
rect 9025 -1236 9031 -1184
rect 9083 -1236 9089 -1184
rect 9025 -1239 9089 -1236
rect 10461 -1256 10546 -1234
rect 10919 -1251 10955 -847
rect 11491 -855 13447 -805
rect 11491 -1183 11556 -855
rect 11491 -1235 11497 -1183
rect 11549 -1235 11556 -1183
rect 11491 -1239 11556 -1235
rect 10461 -1308 10478 -1256
rect 10530 -1308 10546 -1256
rect 10197 -1325 10265 -1323
rect 10197 -1336 10205 -1325
rect 9841 -1373 10205 -1336
rect 9841 -2099 9894 -1373
rect 10197 -1377 10205 -1373
rect 10257 -1377 10265 -1325
rect 10197 -1384 10265 -1377
rect 10461 -1377 10546 -1308
rect 10769 -1257 10955 -1251
rect 10769 -1309 10775 -1257
rect 10827 -1309 10955 -1257
rect 10769 -1315 10955 -1309
rect 11061 -1254 11282 -1248
rect 13408 -1249 13447 -855
rect 11061 -1286 11220 -1254
rect 11061 -1377 11091 -1286
rect 11140 -1306 11220 -1286
rect 11272 -1306 11282 -1254
rect 11140 -1314 11282 -1306
rect 13232 -1254 13447 -1249
rect 13232 -1306 13244 -1254
rect 13296 -1306 13447 -1254
rect 13232 -1313 13447 -1306
rect 10461 -1415 11091 -1377
rect 10870 -1419 11091 -1415
rect 12664 -1327 12738 -1323
rect 12664 -1379 12674 -1327
rect 12726 -1379 12738 -1327
rect 10870 -1444 10906 -1419
rect 10878 -1651 10906 -1444
rect 12664 -1432 12738 -1379
rect 12664 -1488 13663 -1432
rect 9842 -2443 9894 -2099
rect 10075 -1680 10906 -1651
rect 10075 -1684 10124 -1680
rect 10456 -1684 10906 -1680
rect 10075 -2050 10103 -1684
rect 11490 -1699 13447 -1670
rect 11490 -2016 11561 -1699
rect 10759 -2019 10907 -2018
rect 10759 -2025 11279 -2019
rect 10075 -2086 10221 -2050
rect 10759 -2077 11221 -2025
rect 11273 -2077 11279 -2025
rect 11490 -2068 11500 -2016
rect 11552 -2068 11561 -2016
rect 11490 -2070 11561 -2068
rect 10759 -2082 11279 -2077
rect 10075 -2138 10166 -2086
rect 10218 -2138 10221 -2086
rect 10075 -2150 10221 -2138
rect 10258 -2083 11279 -2082
rect 10258 -2088 10811 -2083
rect 13402 -2086 13447 -1699
rect 10258 -2140 10264 -2088
rect 10316 -2140 10811 -2088
rect 13236 -2090 13447 -2086
rect 10258 -2146 10811 -2140
rect 12664 -2128 12739 -2123
rect 12664 -2180 12674 -2128
rect 12726 -2180 12739 -2128
rect 13236 -2142 13242 -2090
rect 13294 -2142 13447 -2090
rect 13236 -2146 13447 -2142
rect 13402 -2147 13447 -2146
rect 12664 -2443 12739 -2180
rect 13603 -2443 13663 -1488
rect 9842 -2480 13665 -2443
rect 9842 -2482 12677 -2480
rect 12738 -2481 13665 -2480
rect -7749 -4432 32575 -4363
rect -7749 -4495 -7629 -4432
rect -7749 -4547 -7725 -4495
rect -7673 -4547 -7629 -4495
rect -7749 -4569 -7629 -4547
rect -7113 -4507 -7020 -4464
rect -7113 -4559 -7089 -4507
rect -7037 -4559 -7020 -4507
rect -7113 -4598 -7020 -4559
rect -5633 -4495 -5513 -4432
rect -5633 -4547 -5609 -4495
rect -5557 -4547 -5513 -4495
rect -5633 -4569 -5513 -4547
rect -4997 -4507 -4904 -4464
rect -4997 -4559 -4973 -4507
rect -4921 -4559 -4904 -4507
rect -4997 -4598 -4904 -4559
rect -3517 -4495 -3397 -4432
rect -3517 -4547 -3493 -4495
rect -3441 -4547 -3397 -4495
rect -3517 -4569 -3397 -4547
rect -2881 -4507 -2788 -4464
rect -2881 -4559 -2857 -4507
rect -2805 -4559 -2788 -4507
rect -2881 -4598 -2788 -4559
rect -1401 -4495 -1281 -4432
rect -1401 -4547 -1377 -4495
rect -1325 -4547 -1281 -4495
rect -1401 -4569 -1281 -4547
rect -765 -4507 -672 -4464
rect -765 -4559 -741 -4507
rect -689 -4559 -672 -4507
rect -765 -4598 -672 -4559
rect 715 -4495 835 -4432
rect 715 -4547 739 -4495
rect 791 -4547 835 -4495
rect 715 -4569 835 -4547
rect 1351 -4507 1444 -4464
rect 1351 -4559 1375 -4507
rect 1427 -4559 1444 -4507
rect 1351 -4598 1444 -4559
rect 2831 -4495 2951 -4432
rect 2831 -4547 2855 -4495
rect 2907 -4547 2951 -4495
rect 2831 -4569 2951 -4547
rect 3467 -4507 3560 -4464
rect 3467 -4559 3491 -4507
rect 3543 -4559 3560 -4507
rect 3467 -4598 3560 -4559
rect 4947 -4495 5067 -4432
rect 4947 -4547 4971 -4495
rect 5023 -4547 5067 -4495
rect 4947 -4569 5067 -4547
rect 5583 -4507 5676 -4464
rect 5583 -4559 5607 -4507
rect 5659 -4559 5676 -4507
rect 5583 -4598 5676 -4559
rect 7063 -4495 7183 -4432
rect 7063 -4547 7087 -4495
rect 7139 -4547 7183 -4495
rect 7063 -4569 7183 -4547
rect 7699 -4507 7792 -4464
rect 7699 -4559 7723 -4507
rect 7775 -4559 7792 -4507
rect 7699 -4598 7792 -4559
rect 9179 -4495 9299 -4432
rect 9179 -4547 9203 -4495
rect 9255 -4547 9299 -4495
rect 9179 -4569 9299 -4547
rect 9815 -4507 9908 -4464
rect 9815 -4559 9839 -4507
rect 9891 -4559 9908 -4507
rect 9815 -4598 9908 -4559
rect 11295 -4495 11415 -4432
rect 11295 -4547 11319 -4495
rect 11371 -4547 11415 -4495
rect 11295 -4569 11415 -4547
rect 11931 -4507 12024 -4464
rect 11931 -4559 11955 -4507
rect 12007 -4559 12024 -4507
rect 11931 -4598 12024 -4559
rect 13411 -4495 13531 -4432
rect 13411 -4547 13435 -4495
rect 13487 -4547 13531 -4495
rect 13411 -4569 13531 -4547
rect 14047 -4507 14140 -4464
rect 14047 -4559 14071 -4507
rect 14123 -4559 14140 -4507
rect 14047 -4598 14140 -4559
rect 15527 -4495 15647 -4432
rect 15527 -4547 15551 -4495
rect 15603 -4547 15647 -4495
rect 15527 -4569 15647 -4547
rect 16163 -4507 16256 -4464
rect 16163 -4559 16187 -4507
rect 16239 -4559 16256 -4507
rect 16163 -4598 16256 -4559
rect 17643 -4495 17763 -4432
rect 17643 -4547 17667 -4495
rect 17719 -4547 17763 -4495
rect 17643 -4569 17763 -4547
rect 18279 -4507 18372 -4464
rect 18279 -4559 18303 -4507
rect 18355 -4559 18372 -4507
rect 18279 -4598 18372 -4559
rect 19759 -4495 19879 -4432
rect 19759 -4547 19783 -4495
rect 19835 -4547 19879 -4495
rect 19759 -4569 19879 -4547
rect 20395 -4507 20488 -4464
rect 20395 -4559 20419 -4507
rect 20471 -4559 20488 -4507
rect 20395 -4598 20488 -4559
rect 21875 -4495 21995 -4432
rect 21875 -4547 21899 -4495
rect 21951 -4547 21995 -4495
rect 21875 -4569 21995 -4547
rect 22511 -4507 22604 -4464
rect 22511 -4559 22535 -4507
rect 22587 -4559 22604 -4507
rect 22511 -4598 22604 -4559
rect 23991 -4495 24111 -4432
rect 23991 -4547 24015 -4495
rect 24067 -4547 24111 -4495
rect 23991 -4569 24111 -4547
rect 24627 -4507 24720 -4464
rect 24627 -4559 24651 -4507
rect 24703 -4559 24720 -4507
rect 24627 -4598 24720 -4559
rect 26107 -4495 26227 -4432
rect 26107 -4547 26131 -4495
rect 26183 -4547 26227 -4495
rect 26107 -4569 26227 -4547
rect 26743 -4507 26836 -4464
rect 26743 -4559 26767 -4507
rect 26819 -4559 26836 -4507
rect 26743 -4598 26836 -4559
rect 28223 -4495 28343 -4432
rect 28223 -4547 28247 -4495
rect 28299 -4547 28343 -4495
rect 28223 -4569 28343 -4547
rect 28859 -4507 28952 -4464
rect 28859 -4559 28883 -4507
rect 28935 -4559 28952 -4507
rect 28859 -4598 28952 -4559
rect 30339 -4495 30459 -4432
rect 30339 -4547 30363 -4495
rect 30415 -4547 30459 -4495
rect 30339 -4569 30459 -4547
rect 30975 -4507 31068 -4464
rect 30975 -4559 30999 -4507
rect 31051 -4559 31068 -4507
rect 30975 -4598 31068 -4559
rect 32455 -4495 32575 -4432
rect 32455 -4547 32479 -4495
rect 32531 -4547 32575 -4495
rect 32455 -4569 32575 -4547
rect 33091 -4507 33184 -4464
rect 33091 -4559 33115 -4507
rect 33167 -4559 33184 -4507
rect 33091 -4598 33184 -4559
rect -8909 -4606 -7020 -4598
rect -8909 -4658 -8858 -4606
rect -8806 -4658 -7020 -4606
rect -8909 -4667 -7020 -4658
rect -6793 -4606 -4904 -4598
rect -6793 -4658 -6742 -4606
rect -6690 -4658 -4904 -4606
rect -6793 -4667 -4904 -4658
rect -4677 -4606 -2788 -4598
rect -4677 -4658 -4626 -4606
rect -4574 -4658 -2788 -4606
rect -4677 -4667 -2788 -4658
rect -2561 -4606 -672 -4598
rect -2561 -4658 -2510 -4606
rect -2458 -4658 -672 -4606
rect -2561 -4667 -672 -4658
rect -445 -4606 1444 -4598
rect -445 -4658 -394 -4606
rect -342 -4658 1444 -4606
rect -445 -4667 1444 -4658
rect 1671 -4606 3560 -4598
rect 1671 -4658 1722 -4606
rect 1774 -4658 3560 -4606
rect 1671 -4667 3560 -4658
rect 3787 -4606 5676 -4598
rect 3787 -4658 3838 -4606
rect 3890 -4658 5676 -4606
rect 3787 -4667 5676 -4658
rect 5903 -4606 7792 -4598
rect 5903 -4658 5954 -4606
rect 6006 -4658 7792 -4606
rect 5903 -4667 7792 -4658
rect 8019 -4606 9908 -4598
rect 8019 -4658 8070 -4606
rect 8122 -4658 9908 -4606
rect 8019 -4667 9908 -4658
rect 10135 -4606 12024 -4598
rect 10135 -4658 10186 -4606
rect 10238 -4658 12024 -4606
rect 10135 -4667 12024 -4658
rect 12251 -4606 14140 -4598
rect 12251 -4658 12302 -4606
rect 12354 -4658 14140 -4606
rect 12251 -4667 14140 -4658
rect 14367 -4606 16256 -4598
rect 14367 -4658 14418 -4606
rect 14470 -4658 16256 -4606
rect 14367 -4667 16256 -4658
rect 16483 -4606 18372 -4598
rect 16483 -4658 16534 -4606
rect 16586 -4658 18372 -4606
rect 16483 -4667 18372 -4658
rect 18599 -4606 20488 -4598
rect 18599 -4658 18650 -4606
rect 18702 -4658 20488 -4606
rect 18599 -4667 20488 -4658
rect 20715 -4606 22604 -4598
rect 20715 -4658 20766 -4606
rect 20818 -4658 22604 -4606
rect 20715 -4667 22604 -4658
rect 22831 -4606 24720 -4598
rect 22831 -4658 22882 -4606
rect 22934 -4658 24720 -4606
rect 22831 -4667 24720 -4658
rect 24947 -4606 26836 -4598
rect 24947 -4658 24998 -4606
rect 25050 -4658 26836 -4606
rect 24947 -4667 26836 -4658
rect 27063 -4606 28952 -4598
rect 27063 -4658 27114 -4606
rect 27166 -4658 28952 -4606
rect 27063 -4667 28952 -4658
rect 29179 -4606 31068 -4598
rect 29179 -4658 29230 -4606
rect 29282 -4658 31068 -4606
rect 29179 -4667 31068 -4658
rect 31295 -4606 33184 -4598
rect 31295 -4658 31346 -4606
rect 31398 -4658 33184 -4606
rect 31295 -4667 33184 -4658
rect 12828 -7629 14422 -7627
rect 12828 -7656 17524 -7629
rect 8082 -7689 10389 -7662
rect 8082 -7850 9897 -7689
rect 9960 -7690 10286 -7689
rect 9960 -7849 10023 -7690
rect 10103 -7849 10174 -7690
rect 10254 -7848 10286 -7690
rect 10366 -7848 10389 -7689
rect 10254 -7849 10389 -7848
rect 9960 -7850 10389 -7849
rect 8082 -7887 10389 -7850
rect 12828 -7882 12896 -7656
rect 14455 -7882 17524 -7656
rect 12828 -7884 14341 -7882
rect 14454 -7884 17524 -7882
rect 12828 -7906 17524 -7884
rect 12828 -7907 14422 -7906
rect 8984 -8654 9262 -8635
rect 8984 -8967 9002 -8654
rect 9241 -8967 9262 -8654
rect 8984 -8986 9262 -8967
rect 16398 -8656 16699 -8645
rect 16398 -9006 16412 -8656
rect 16685 -9006 16699 -8656
rect 16398 -9016 16699 -9006
rect 17292 -9253 17522 -9211
rect 17292 -9429 17324 -9253
rect 17486 -9429 17522 -9253
rect 17292 -10179 17522 -9429
rect 17292 -10355 17324 -10179
rect 17486 -10355 17522 -10179
rect 17292 -10371 17522 -10355
rect 7986 -10613 8378 -10557
rect 7986 -10831 8042 -10613
rect 8288 -10831 8378 -10613
rect 7986 -11325 8378 -10831
rect 7986 -11549 8076 -11325
rect 8324 -11549 8378 -11325
rect 7986 -11587 8378 -11549
rect 5190 -12920 7102 -12739
rect 5190 -13561 5392 -12920
rect 6904 -13561 7102 -12920
rect 9950 -13161 10094 -13153
rect 9950 -13267 9970 -13161
rect 10076 -13267 10094 -13161
rect 9950 -13277 10094 -13267
rect 12616 -13161 12760 -13153
rect 12616 -13267 12634 -13161
rect 12740 -13267 12760 -13161
rect 12616 -13277 12760 -13267
rect 15277 -13161 15423 -13153
rect 15277 -13267 15296 -13161
rect 15402 -13267 15423 -13161
rect 15277 -13278 15423 -13267
rect 5190 -13772 7102 -13561
rect 18860 -13362 20667 -13165
rect 17292 -14061 17522 -14019
rect 8951 -14220 9229 -14206
rect 8951 -14525 8991 -14220
rect 9174 -14525 9229 -14220
rect 8951 -14557 9229 -14525
rect 17292 -14237 17324 -14061
rect 17486 -14237 17522 -14061
rect 17292 -14987 17522 -14237
rect 18860 -14064 19119 -13362
rect 20321 -14064 20667 -13362
rect 18860 -14314 20667 -14064
rect 8038 -15059 8268 -15017
rect 8038 -15235 8070 -15059
rect 8232 -15235 8268 -15059
rect 17292 -15163 17324 -14987
rect 17486 -15163 17522 -14987
rect 17292 -15179 17522 -15163
rect 8038 -15985 8268 -15235
rect 8038 -16161 8070 -15985
rect 8232 -16161 8268 -15985
rect 8038 -16177 8268 -16161
rect 9942 -18880 10096 -18870
rect 9942 -18986 9964 -18880
rect 10070 -18986 10096 -18880
rect 9942 -18997 10096 -18986
rect 12626 -18885 12751 -18869
rect 12626 -18979 12640 -18885
rect 12732 -18979 12751 -18885
rect 12626 -18991 12751 -18979
rect 15290 -18885 15415 -18865
rect 15290 -18979 15306 -18885
rect 15398 -18979 15415 -18885
rect 15290 -18991 15415 -18979
rect 16195 -19562 16511 -19542
rect 16195 -19911 16230 -19562
rect 16476 -19911 16511 -19562
rect 16851 -19728 16995 -19714
rect 16851 -19839 16870 -19728
rect 16974 -19839 16995 -19728
rect 16851 -19853 16995 -19839
rect 16195 -19922 16511 -19911
rect 8040 -20041 8268 -19999
rect 8040 -20217 8070 -20041
rect 8232 -20217 8268 -20041
rect 8040 -20889 8268 -20217
rect 8932 -20119 9165 -20099
rect 8932 -20129 8963 -20119
rect 9119 -20129 9165 -20119
rect 8932 -20385 8952 -20129
rect 9133 -20385 9165 -20129
rect 8932 -20391 8963 -20385
rect 9119 -20391 9165 -20385
rect 8932 -20424 9165 -20391
rect 16500 -20399 16603 -20389
rect 16500 -20503 16510 -20399
rect 16589 -20503 16603 -20399
rect 16500 -20515 16603 -20503
rect 16887 -20400 16990 -20387
rect 16887 -20503 16900 -20400
rect 16974 -20503 16990 -20400
rect 16887 -20513 16990 -20503
rect 8040 -21065 8070 -20889
rect 8232 -21065 8268 -20889
rect 8040 -21081 8268 -21065
rect 17122 -20743 17498 -20693
rect 17122 -21039 17164 -20743
rect 17416 -21039 17498 -20743
rect 17122 -23033 17498 -21039
rect 17122 -23267 17202 -23033
rect 17426 -23267 17498 -23033
rect 17122 -23299 17498 -23267
rect 9942 -24781 10096 -24760
rect 9942 -24875 9972 -24781
rect 10064 -24875 10096 -24781
rect 9942 -24887 10096 -24875
rect 12616 -24781 12763 -24765
rect 12616 -24875 12642 -24781
rect 12734 -24875 12763 -24781
rect 12616 -24888 12763 -24875
rect 15284 -24781 15431 -24767
rect 15284 -24875 15308 -24781
rect 15400 -24875 15431 -24781
rect 15284 -24890 15431 -24875
rect 7986 -25151 8498 -25033
rect 7986 -25413 8086 -25151
rect 8380 -25413 8498 -25151
rect 7986 -25573 8498 -25413
<< via2 >>
rect -18978 55462 -17592 56190
rect -14978 55462 -13592 56190
rect -10978 55462 -9592 56190
rect -6978 55462 -5592 56190
rect -2978 55462 -1592 56190
rect 1022 55462 2408 56190
rect 5022 55462 6408 56190
rect 9022 55462 10408 56190
rect 13022 55462 14408 56190
rect 17022 55462 18408 56190
rect 21022 55462 22408 56190
rect 25022 55462 26408 56190
rect 29022 55462 30408 56190
rect 33022 55462 34408 56190
rect 37022 55462 38408 56190
rect -20714 53298 -19328 54026
rect -20714 49298 -19328 50026
rect -20714 45298 -19328 46026
rect -20714 41298 -19328 42026
rect 16720 51076 17836 51868
rect 22192 51314 23050 52102
rect 37064 52260 38450 52988
rect 388 44886 550 44958
rect 6284 44924 6446 44996
rect 17176 44932 17338 45004
rect 37064 48260 38450 48988
rect 22446 44856 22608 44928
rect 37064 44260 38450 44988
rect -20714 37298 -19328 38026
rect 37064 40260 38450 40988
rect -13876 36162 -13688 36338
rect -11578 36390 -11378 36624
rect -20714 33298 -19328 34026
rect -20714 29298 -19328 30026
rect -20714 25298 -19328 26026
rect 508 34122 670 34194
rect -8174 27104 -6984 27902
rect 5434 34192 5596 34264
rect 11372 34134 11636 34230
rect 16704 34044 16866 34116
rect 9172 28064 9526 28258
rect 37064 36260 38450 36988
rect 22228 34132 22390 34204
rect 20 25118 728 26050
rect 15928 25912 17090 27028
rect 37064 32260 38450 32988
rect 37064 28260 38450 28988
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -96044 17274 -95512 17740
rect -96044 15274 -95512 15740
rect -96044 13274 -95512 13740
rect -96044 11274 -95512 11740
rect -96044 9274 -95512 9740
rect -96044 7274 -95512 7740
rect -96044 5274 -95512 5740
rect -20714 21298 -19328 22026
rect -27644 19274 -27112 19740
rect -27644 17274 -27112 17740
rect -20714 17298 -19328 18026
rect -27644 15274 -27112 15740
rect -18052 14180 -16666 14908
rect 37064 24260 38450 24988
rect 9218 20792 9482 21060
rect 16524 20618 16754 20860
rect 37064 20260 38450 20988
rect 13138 18134 13424 18404
rect 37064 16260 38450 16988
rect -14052 14180 -12666 14908
rect -10052 14180 -8666 14908
rect -6052 14180 -4666 14908
rect -2052 14180 -666 14908
rect 1948 14180 3334 14908
rect 5948 14180 7334 14908
rect 9948 14180 11334 14908
rect 13948 14180 15334 14908
rect 17948 14180 19334 14908
rect 21948 14180 23334 14908
rect 25948 14180 27334 14908
rect 29948 14180 31334 14908
rect 33948 14180 35334 14908
rect -27644 13274 -27112 13740
rect -27644 11274 -27112 11740
rect -27644 9274 -27112 9740
rect 5368 9504 5800 9508
rect 5368 9434 5800 9504
rect 5368 9186 5800 9188
rect 5368 9114 5800 9186
rect 5368 8796 5800 8870
rect 5800 8796 5802 8870
rect 5368 8794 5802 8796
rect -27644 7274 -27112 7740
rect 10564 10072 10996 10144
rect 10564 9752 10996 9824
rect -27644 5274 -27112 5740
rect 1374 5776 1700 6016
rect 6262 5854 6588 6094
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect 11574 5642 11900 5882
rect 18000 11574 18960 12068
rect 14846 8164 15278 8234
rect 17010 5584 17336 5824
rect 16664 5008 16746 5108
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect 10738 3768 10862 3772
rect 10738 3716 10862 3768
rect 16256 3686 16414 3804
rect -61864 2878 -61806 2882
rect -61864 2826 -61806 2878
rect -61464 2878 -61406 2882
rect -61464 2826 -61406 2878
rect 10728 2536 10846 2598
rect 26138 3246 26538 3638
rect 26690 2190 26780 2264
rect 31320 2012 31382 2074
rect 3524 1204 4484 1698
rect 10946 1020 11906 1514
rect 17578 1338 18538 1832
rect 32424 1746 32904 2206
rect 9002 -8967 9241 -8654
rect 16412 -8669 16685 -8656
rect 16412 -8990 16433 -8669
rect 16433 -8990 16655 -8669
rect 16655 -8990 16685 -8669
rect 16412 -9006 16685 -8990
rect 8076 -11549 8324 -11325
rect 5392 -12977 6904 -12920
rect 5392 -13467 5413 -12977
rect 5413 -13467 6710 -12977
rect 6710 -13467 6904 -12977
rect 5392 -13561 6904 -13467
rect 9970 -13267 10076 -13161
rect 12634 -13267 12740 -13161
rect 15296 -13267 15402 -13161
rect 8991 -14525 9174 -14220
rect 19119 -13391 20321 -13362
rect 19119 -13987 19172 -13391
rect 19172 -13987 20172 -13391
rect 20172 -13987 20321 -13391
rect 19119 -14064 20321 -13987
rect 9964 -18986 10070 -18880
rect 12640 -18979 12732 -18885
rect 15306 -18979 15398 -18885
rect 16230 -19578 16476 -19562
rect 16230 -19895 16242 -19578
rect 16242 -19895 16458 -19578
rect 16458 -19895 16476 -19578
rect 16230 -19911 16476 -19895
rect 16870 -19747 16974 -19728
rect 16870 -19819 16887 -19747
rect 16887 -19819 16958 -19747
rect 16958 -19819 16974 -19747
rect 16870 -19839 16974 -19819
rect 8952 -20385 8963 -20129
rect 8963 -20385 9119 -20129
rect 9119 -20385 9133 -20129
rect 16510 -20415 16589 -20399
rect 16510 -20488 16523 -20415
rect 16523 -20488 16579 -20415
rect 16579 -20488 16589 -20415
rect 16510 -20503 16589 -20488
rect 16900 -20415 16974 -20400
rect 16900 -20488 16912 -20415
rect 16912 -20488 16968 -20415
rect 16968 -20488 16974 -20415
rect 16900 -20503 16974 -20488
rect 9972 -24875 10064 -24781
rect 12642 -24875 12734 -24781
rect 15308 -24875 15400 -24781
rect 8086 -25413 8380 -25151
<< metal3 >>
rect -19220 56190 -17382 56450
rect -19220 55462 -18978 56190
rect -17592 55462 -17382 56190
rect -19220 55220 -17382 55462
rect -15220 56190 -13382 56450
rect -15220 55462 -14978 56190
rect -13592 55462 -13382 56190
rect -15220 55220 -13382 55462
rect -11220 56190 -9382 56450
rect -11220 55462 -10978 56190
rect -9592 55462 -9382 56190
rect -11220 55220 -9382 55462
rect -7220 56190 -5382 56450
rect -7220 55462 -6978 56190
rect -5592 55462 -5382 56190
rect -7220 55220 -5382 55462
rect -3220 56190 -1382 56450
rect -3220 55462 -2978 56190
rect -1592 55462 -1382 56190
rect -3220 55220 -1382 55462
rect 780 56190 2618 56450
rect 780 55462 1022 56190
rect 2408 55462 2618 56190
rect 780 55220 2618 55462
rect 4780 56190 6618 56450
rect 4780 55462 5022 56190
rect 6408 55462 6618 56190
rect 4780 55220 6618 55462
rect 8780 56190 10618 56450
rect 8780 55462 9022 56190
rect 10408 55462 10618 56190
rect 8780 55220 10618 55462
rect 12780 56190 14618 56450
rect 12780 55462 13022 56190
rect 14408 55462 14618 56190
rect 12780 55220 14618 55462
rect 16780 56190 18618 56450
rect 16780 55462 17022 56190
rect 18408 55462 18618 56190
rect 16780 55220 18618 55462
rect 20780 56190 22618 56450
rect 20780 55462 21022 56190
rect 22408 55462 22618 56190
rect 20780 55220 22618 55462
rect 24780 56190 26618 56450
rect 24780 55462 25022 56190
rect 26408 55462 26618 56190
rect 24780 55220 26618 55462
rect 28780 56190 30618 56450
rect 28780 55462 29022 56190
rect 30408 55462 30618 56190
rect 28780 55220 30618 55462
rect 32780 56190 34618 56450
rect 32780 55462 33022 56190
rect 34408 55462 34618 56190
rect 32780 55220 34618 55462
rect 36780 56190 38618 56450
rect 36780 55462 37022 56190
rect 38408 55462 38618 56190
rect 36780 55220 38618 55462
rect -20956 54026 -19118 54286
rect -20956 53298 -20714 54026
rect -19328 53298 -19118 54026
rect -20956 53056 -19118 53298
rect 36822 52988 38660 53256
rect 22030 52238 32260 52264
rect 36822 52260 37064 52988
rect 38450 52260 38660 52988
rect 22030 52102 32348 52238
rect -14642 51868 18546 52000
rect -14642 51076 16720 51868
rect 17836 51076 18546 51868
rect 22030 51314 22192 52102
rect 23050 51314 32348 52102
rect 36822 52018 38660 52260
rect 22030 51220 32348 51314
rect -14642 50738 18546 51076
rect -20956 50026 -19118 50286
rect -20956 49298 -20714 50026
rect -19328 49298 -19118 50026
rect -20956 49056 -19118 49298
rect -20956 46026 -19118 46286
rect -20956 45298 -20714 46026
rect -19328 45298 -19118 46026
rect -20956 45056 -19118 45298
rect -20956 42026 -19118 42286
rect -20956 41298 -20714 42026
rect -19328 41298 -19118 42026
rect -20956 41056 -19118 41298
rect -20956 38026 -19118 38286
rect -20956 37298 -20714 38026
rect -19328 37298 -19118 38026
rect -20956 37056 -19118 37298
rect -14362 36338 -13054 50738
rect -8835 45298 29386 50416
rect -8835 45296 16552 45298
rect -8835 45266 5958 45296
rect -8835 45144 40 45266
rect 930 45144 5958 45266
rect 6860 45144 16552 45296
rect 18186 45246 29386 45298
rect 18186 45144 22154 45246
rect 23066 45144 29386 45246
rect -14362 36162 -13876 36338
rect -13688 36162 -13054 36338
rect -11614 36624 -11334 36712
rect -11614 36390 -11578 36624
rect -11378 36390 -11334 36624
rect -11614 36314 -11334 36390
rect -20956 34026 -19118 34286
rect -20956 33298 -20714 34026
rect -19328 33298 -19118 34026
rect -20956 33056 -19118 33298
rect -20956 30026 -19118 30286
rect -20956 29298 -20714 30026
rect -19328 29298 -19118 30026
rect -20956 29056 -19118 29298
rect -20956 26026 -19118 26286
rect -20956 25298 -20714 26026
rect -19328 25298 -19118 26026
rect -20956 25056 -19118 25298
rect -14362 22596 -13054 36162
rect -8802 33710 -3695 45144
rect 6260 44996 6478 45026
rect 364 44958 582 44988
rect 6260 44968 6284 44996
rect 364 44930 388 44958
rect 362 44886 388 44930
rect 550 44886 582 44958
rect 362 44828 582 44886
rect 6258 44924 6284 44968
rect 6446 44924 6478 44996
rect 17152 45004 17370 45034
rect 17152 44976 17176 45004
rect 6258 44828 6478 44924
rect 17150 44932 17176 44976
rect 17338 44932 17370 45004
rect 17150 44868 17370 44932
rect 22422 44928 22640 44958
rect 22422 44900 22446 44928
rect -3298 44690 1748 44828
rect -3298 39814 1752 44690
rect 2226 44674 7272 44828
rect 2226 41396 7286 44674
rect -3298 39710 1748 39814
rect 2226 39710 7272 41396
rect 7731 39710 12777 44828
rect 13215 39750 18261 44868
rect 22420 44856 22446 44900
rect 22608 44856 22640 44928
rect 22420 44828 22640 44856
rect 24147 44828 29254 45144
rect 18740 39710 23786 44828
rect 24147 39710 29286 44828
rect 7772 39292 12746 39710
rect 2208 39239 7194 39252
rect -3196 34194 1790 39192
rect 2208 34264 7278 39239
rect 2208 34226 5434 34264
rect -3196 34166 508 34194
rect 482 34122 508 34166
rect 670 34166 1790 34194
rect 5408 34192 5434 34226
rect 5596 34226 7278 34264
rect 7772 34266 12759 39292
rect 7772 34238 12746 34266
rect 13275 34247 18261 39352
rect 24147 39272 29254 39710
rect 13275 34246 18142 34247
rect 5596 34192 5628 34226
rect 6939 34224 7278 34226
rect 11040 34230 12086 34238
rect 670 34122 702 34166
rect 482 34046 702 34122
rect 5408 34116 5628 34192
rect 11040 34134 11372 34230
rect 11636 34134 12086 34230
rect 11040 34082 12086 34134
rect 16672 34116 16930 34246
rect 18740 34204 23786 39272
rect 18740 34166 22228 34204
rect 16672 34070 16704 34116
rect 16678 34044 16704 34070
rect 16866 34070 16930 34116
rect 22202 34132 22228 34166
rect 22390 34166 23786 34204
rect 24147 34166 29286 39272
rect 22390 34132 22422 34166
rect 16866 34044 16898 34070
rect 22202 34056 22422 34132
rect 16678 33968 16898 34044
rect -3298 33710 1748 33728
rect 2226 33710 7272 33728
rect 7731 33710 12777 33728
rect 13215 33710 16372 33768
rect -8901 33678 16372 33710
rect 17296 33710 18261 33768
rect 24147 33728 29254 34166
rect 18740 33710 23786 33728
rect 24147 33710 29286 33728
rect 17296 33678 29286 33710
rect -8901 28616 29286 33678
rect -8901 28471 29254 28616
rect -8402 27902 -6746 28471
rect 8960 28258 9880 28336
rect 8960 28064 9172 28258
rect 9526 28064 9880 28258
rect 8960 28032 9880 28064
rect -8402 27104 -8174 27902
rect -6984 27104 -6746 27902
rect 15928 27260 17416 27400
rect -8402 26890 -6746 27104
rect 15604 27028 17416 27260
rect -8390 26888 -6772 26890
rect -240 26050 1286 26608
rect -240 25118 20 26050
rect 728 25118 1286 26050
rect 15604 25912 15928 27028
rect 17090 25912 17416 27028
rect 15604 25342 17416 25912
rect -240 22596 1286 25118
rect 15622 22624 17148 25342
rect 30162 24238 32348 51220
rect 36822 48988 38660 49256
rect 36822 48260 37064 48988
rect 38450 48260 38660 48988
rect 36822 48018 38660 48260
rect 36822 44988 38660 45256
rect 36822 44260 37064 44988
rect 38450 44260 38660 44988
rect 36822 44018 38660 44260
rect 36822 40988 38660 41256
rect 36822 40260 37064 40988
rect 38450 40260 38660 40988
rect 36822 40018 38660 40260
rect 36822 36988 38660 37256
rect 36822 36260 37064 36988
rect 38450 36260 38660 36988
rect 36822 36018 38660 36260
rect 36822 32988 38660 33256
rect 36822 32260 37064 32988
rect 38450 32260 38660 32988
rect 36822 32018 38660 32260
rect 36822 28988 38660 29256
rect 36822 28260 37064 28988
rect 38450 28260 38660 28988
rect 36822 28018 38660 28260
rect 36822 24988 38660 25256
rect 36822 24260 37064 24988
rect 38450 24260 38660 24988
rect 9478 22596 11254 22624
rect -20956 22026 -19118 22286
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -96266 13740 -95320 15274
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -96266 4182 -95320 5274
rect -27834 19740 -26806 21200
rect -20956 21298 -20714 22026
rect -19328 21298 -19118 22026
rect -14362 21616 11254 22596
rect -20956 21056 -19118 21298
rect -14268 21060 11254 21616
rect -14268 20792 9218 21060
rect 9482 20820 11254 21060
rect 15604 21818 17416 22624
rect 30022 21818 32394 24238
rect 36822 24018 38660 24260
rect 15604 20860 32394 21818
rect 9482 20792 11206 20820
rect -14268 20260 11206 20792
rect 15604 20618 16524 20860
rect 16754 20618 32394 20860
rect 15604 19958 32394 20618
rect 36822 20988 38660 21256
rect 36822 20260 37064 20988
rect 38450 20260 38660 20988
rect 36822 20018 38660 20260
rect 30022 19912 32394 19958
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -27834 17740 -26806 19274
rect 13066 18404 13490 18476
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -27834 15740 -26806 17274
rect -20956 18026 -19118 18286
rect 13066 18134 13138 18404
rect 13424 18134 13490 18404
rect 13066 18052 13490 18134
rect -20956 17298 -20714 18026
rect -19328 17298 -19118 18026
rect -20956 17056 -19118 17298
rect 36822 16988 38660 17256
rect 36822 16260 37064 16988
rect 38450 16260 38660 16988
rect 36822 16018 38660 16260
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -27834 13740 -26806 15274
rect -18294 14908 -16456 15184
rect -18294 14180 -18052 14908
rect -16666 14180 -16456 14908
rect -18294 13938 -16456 14180
rect -14294 15084 -14106 15180
rect -13566 15084 -12456 15180
rect -14294 14908 -12456 15084
rect -14294 14180 -14052 14908
rect -12666 14180 -12456 14908
rect -14294 13938 -12456 14180
rect -10294 14908 -8456 15180
rect -10294 14180 -10052 14908
rect -8666 14180 -8456 14908
rect -10294 13938 -8456 14180
rect -6294 14908 -4456 15180
rect -6294 14180 -6052 14908
rect -4666 14180 -4456 14908
rect -6294 13938 -4456 14180
rect -2294 14908 -456 15180
rect -2294 14180 -2052 14908
rect -666 14180 -456 14908
rect -2294 13938 -456 14180
rect 1706 14908 3544 15180
rect 1706 14180 1948 14908
rect 3334 14180 3544 14908
rect 1706 13938 3544 14180
rect 5706 14908 7544 15180
rect 5706 14180 5948 14908
rect 7334 14180 7544 14908
rect 5706 13938 7544 14180
rect 9706 14908 11544 15180
rect 9706 14180 9948 14908
rect 11334 14180 11544 14908
rect 9706 13938 11544 14180
rect 13706 14908 15544 15180
rect 13706 14180 13948 14908
rect 15334 14180 15544 14908
rect 13706 13938 15544 14180
rect 17706 14908 19544 15180
rect 17706 14180 17948 14908
rect 19334 14180 19544 14908
rect 17706 13938 19544 14180
rect 21706 14908 23544 15180
rect 21706 14180 21948 14908
rect 23334 14180 23544 14908
rect 21706 13938 23544 14180
rect 25706 14908 27544 15180
rect 25706 14180 25948 14908
rect 27334 14180 27544 14908
rect 25706 13938 27544 14180
rect 29706 14908 31544 15180
rect 29706 14180 29948 14908
rect 31334 14180 31544 14908
rect 29706 13938 31544 14180
rect 33706 14908 35544 15180
rect 33706 14180 33948 14908
rect 35334 14180 35544 14908
rect 33706 13938 35544 14180
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -27834 11740 -26806 13274
rect 17792 12068 19104 12262
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect -27834 9740 -26806 11274
rect 10308 11788 10394 11834
rect 17792 11788 18000 12068
rect 10308 11704 18000 11788
rect 10308 9980 10394 11704
rect 17792 11574 18000 11704
rect 18960 11574 19104 12068
rect 17792 11354 19104 11574
rect 10550 10144 11004 10158
rect 10550 10072 10564 10144
rect 10996 10072 11004 10144
rect 10550 9980 11004 10072
rect 10308 9908 11004 9980
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect 10550 9824 11004 9908
rect 10550 9752 10564 9824
rect 10996 9752 11004 9824
rect 10550 9736 11004 9752
rect 5354 9508 5812 9526
rect 5354 9434 5368 9508
rect 5800 9434 5812 9508
rect 5354 9416 5812 9434
rect 5498 9346 5564 9416
rect 5498 9278 6388 9346
rect -27834 7740 -26806 9274
rect 5354 9188 5814 9202
rect 5354 9114 5368 9188
rect 5800 9114 5814 9188
rect 5354 8994 5814 9114
rect 6324 8994 6388 9278
rect 5354 8930 6396 8994
rect 5354 8870 5814 8930
rect 5354 8794 5368 8870
rect 5802 8794 5814 8870
rect 5354 8776 5814 8794
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -27834 5740 -26806 7274
rect 6330 6190 6396 8930
rect 14836 8238 15290 8248
rect 17084 8238 17146 8240
rect 14836 8234 17206 8238
rect 14836 8164 14846 8234
rect 15278 8164 17206 8234
rect 14836 8162 17206 8164
rect 14836 8152 15290 8162
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 1280 5776 1374 6016
rect 1700 5776 1794 6016
rect 1280 5678 1794 5776
rect 6168 6094 6682 6190
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 6168 5756 6682 5854
rect 11480 5882 11994 5978
rect 17084 5920 17146 8162
rect 11480 5642 11574 5882
rect 11900 5642 11994 5882
rect 11480 5544 11994 5642
rect 16916 5824 17430 5920
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -96396 3740 -62544 3910
rect -27834 3846 -26806 5274
rect 16638 5108 16776 5136
rect 16638 5008 16664 5108
rect 16746 5008 16776 5108
rect 16638 4978 16776 5008
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -96396 2966 -62544 3274
rect -60278 3740 -26756 3846
rect 16228 3804 16448 3842
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect 10712 3772 10888 3786
rect 10712 3716 10738 3772
rect 10862 3762 10888 3772
rect 16228 3762 16256 3804
rect 10862 3716 16256 3762
rect 10712 3698 16256 3716
rect 16228 3686 16256 3698
rect 16414 3686 16448 3804
rect 16228 3656 16448 3686
rect -60278 3224 -26756 3274
rect -61896 2890 -61292 2894
rect -61896 2826 -61864 2890
rect -61800 2826 -61464 2890
rect -61400 2826 -61292 2890
rect -61896 2812 -61292 2826
rect 16676 2634 16742 4978
rect 26106 3638 26596 3676
rect 26106 3246 26138 3638
rect 26538 3246 26596 3638
rect 26106 3216 26596 3246
rect 16518 2632 16792 2634
rect 10754 2608 16792 2632
rect 10714 2598 16792 2608
rect 10714 2536 10728 2598
rect 10846 2546 16792 2598
rect 10846 2536 10860 2546
rect 16518 2544 16792 2546
rect 10714 2524 10860 2536
rect 26678 2264 26796 2282
rect 26678 2190 26690 2264
rect 26780 2260 26796 2264
rect 26780 2200 31382 2260
rect 26780 2190 26796 2200
rect 26678 2172 26796 2190
rect 31320 2090 31382 2200
rect 32364 2206 32976 2274
rect 31306 2074 31396 2090
rect 3316 1698 4628 1892
rect 17370 1832 18682 2026
rect 31306 2012 31320 2074
rect 31382 2012 31396 2074
rect 31306 1998 31396 2012
rect 3316 1204 3524 1698
rect 4484 1204 4628 1698
rect 3316 984 4628 1204
rect 10738 1514 12050 1708
rect 10738 1020 10946 1514
rect 11906 1020 12050 1514
rect 17370 1338 17578 1832
rect 18538 1338 18682 1832
rect 32364 1746 32424 2206
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 17370 1118 18682 1338
rect 10738 800 12050 1020
rect 8984 -8654 9262 -8635
rect 8984 -8967 9002 -8654
rect 9241 -8967 9262 -8654
rect 8984 -8986 9262 -8967
rect 16394 -8656 16700 -8641
rect 16394 -9006 16412 -8656
rect 16685 -9006 16700 -8656
rect 16394 -9018 16700 -9006
rect 7986 -11325 8500 -11247
rect 7986 -11549 8076 -11325
rect 8324 -11549 8500 -11325
rect 5190 -12769 7110 -12743
rect 5190 -13742 5237 -12769
rect 7037 -13742 7110 -12769
rect 7986 -25151 8500 -11549
rect 9950 -13161 10094 -13153
rect 9950 -13267 9970 -13161
rect 10076 -13267 10094 -13161
rect 9950 -13277 10094 -13267
rect 12616 -13161 12760 -13153
rect 12616 -13267 12634 -13161
rect 12740 -13267 12760 -13161
rect 12616 -13277 12760 -13267
rect 15277 -13161 15423 -13153
rect 15277 -13267 15296 -13161
rect 15402 -13267 15423 -13161
rect 15277 -13278 15423 -13267
rect 18889 -13305 20633 -13204
rect 18889 -14098 18999 -13305
rect 20398 -14098 20633 -13305
rect 8951 -14220 9229 -14206
rect 8951 -14525 8991 -14220
rect 9174 -14525 9229 -14220
rect 18889 -14247 20633 -14098
rect 8951 -14557 9229 -14525
rect 9942 -18880 10096 -18870
rect 9942 -18986 9964 -18880
rect 10070 -18986 10096 -18880
rect 9942 -18997 10096 -18986
rect 12626 -18885 12751 -18869
rect 12626 -18979 12640 -18885
rect 12732 -18979 12751 -18885
rect 12626 -18991 12751 -18979
rect 15290 -18885 15415 -18865
rect 15290 -18979 15306 -18885
rect 15398 -18979 15415 -18885
rect 15290 -18991 15415 -18979
rect 16191 -19562 16520 -19538
rect 16191 -19911 16230 -19562
rect 16476 -19911 16520 -19562
rect 16851 -19728 16995 -19714
rect 16851 -19839 16870 -19728
rect 16974 -19839 16995 -19728
rect 16851 -19853 16995 -19839
rect 16191 -19931 16520 -19911
rect 8922 -20129 9166 -20098
rect 8922 -20385 8952 -20129
rect 9133 -20385 9166 -20129
rect 8922 -20424 9166 -20385
rect 16498 -20399 16599 -20390
rect 16498 -20503 16510 -20399
rect 16589 -20503 16599 -20399
rect 16498 -20513 16599 -20503
rect 16886 -20400 16988 -20387
rect 16886 -20503 16900 -20400
rect 16974 -20503 16988 -20400
rect 16886 -20515 16988 -20503
rect 9942 -24781 10096 -24760
rect 9942 -24875 9972 -24781
rect 10064 -24875 10096 -24781
rect 9942 -24887 10096 -24875
rect 12616 -24781 12763 -24765
rect 12616 -24875 12642 -24781
rect 12734 -24875 12763 -24781
rect 12616 -24888 12763 -24875
rect 15284 -24781 15431 -24767
rect 15284 -24875 15308 -24781
rect 15400 -24875 15431 -24781
rect 15284 -24890 15431 -24875
rect 7986 -25413 8086 -25151
rect 8380 -25413 8500 -25151
rect 7986 -25567 8500 -25413
<< via3 >>
rect -18978 55462 -17592 56190
rect -14978 55462 -13592 56190
rect -10978 55462 -9592 56190
rect -6978 55462 -5592 56190
rect -2978 55462 -1592 56190
rect 1022 55462 2408 56190
rect 5022 55462 6408 56190
rect 9022 55462 10408 56190
rect 13022 55462 14408 56190
rect 17022 55462 18408 56190
rect 21022 55462 22408 56190
rect 25022 55462 26408 56190
rect 29022 55462 30408 56190
rect 33022 55462 34408 56190
rect 37022 55462 38408 56190
rect -20714 53298 -19328 54026
rect 37064 52260 38450 52988
rect -20714 49298 -19328 50026
rect -20714 45298 -19328 46026
rect -20714 41298 -19328 42026
rect -20714 37298 -19328 38026
rect -11578 36390 -11378 36624
rect -20714 33298 -19328 34026
rect -20714 29298 -19328 30026
rect -20714 25298 -19328 26026
rect 9172 28064 9526 28258
rect -8174 27104 -6984 27902
rect 37064 48260 38450 48988
rect 37064 44260 38450 44988
rect 37064 40260 38450 40988
rect 37064 36260 38450 36988
rect 37064 32260 38450 32988
rect 37064 28260 38450 28988
rect 37064 24260 38450 24988
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -96044 17274 -95512 17740
rect -96044 15274 -95512 15740
rect -96044 13274 -95512 13740
rect -96044 11274 -95512 11740
rect -96044 9274 -95512 9740
rect -96044 7274 -95512 7740
rect -96044 5274 -95512 5740
rect -20714 21298 -19328 22026
rect 37064 20260 38450 20988
rect -27644 19274 -27112 19740
rect -27644 17274 -27112 17740
rect 13138 18134 13424 18404
rect -20714 17298 -19328 18026
rect 37064 16260 38450 16988
rect -27644 15274 -27112 15740
rect -18052 14180 -16666 14908
rect -14052 14180 -12666 14908
rect -10052 14180 -8666 14908
rect -6052 14180 -4666 14908
rect -2052 14180 -666 14908
rect 1948 14180 3334 14908
rect 5948 14180 7334 14908
rect 9948 14180 11334 14908
rect 13948 14180 15334 14908
rect 17948 14180 19334 14908
rect 21948 14180 23334 14908
rect 25948 14180 27334 14908
rect 29948 14180 31334 14908
rect 33948 14180 35334 14908
rect -27644 13274 -27112 13740
rect -27644 11274 -27112 11740
rect 18000 11574 18960 12068
rect -27644 9274 -27112 9740
rect -27644 7274 -27112 7740
rect -27644 5274 -27112 5740
rect 1374 5776 1700 6016
rect 6262 5854 6588 6094
rect 11574 5642 11900 5882
rect 17010 5584 17336 5824
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect -61864 2882 -61800 2890
rect -61864 2826 -61806 2882
rect -61806 2826 -61800 2882
rect -61464 2882 -61400 2890
rect -61464 2826 -61406 2882
rect -61406 2826 -61400 2882
rect 26138 3246 26538 3638
rect 3524 1204 4484 1698
rect 10946 1020 11906 1514
rect 17578 1338 18538 1832
rect 32424 1746 32904 2206
rect 9002 -8967 9241 -8654
rect 16412 -9006 16685 -8656
rect 5237 -12920 7037 -12769
rect 5237 -13561 5392 -12920
rect 5392 -13561 6904 -12920
rect 6904 -13561 7037 -12920
rect 5237 -13742 7037 -13561
rect 9970 -13267 10076 -13161
rect 12634 -13267 12740 -13161
rect 15296 -13267 15402 -13161
rect 18999 -13362 20398 -13305
rect 18999 -14064 19119 -13362
rect 19119 -14064 20321 -13362
rect 20321 -14064 20398 -13362
rect 18999 -14098 20398 -14064
rect 8991 -14525 9174 -14220
rect 9964 -18986 10070 -18880
rect 12640 -18979 12732 -18885
rect 15306 -18979 15398 -18885
rect 16230 -19911 16476 -19562
rect 16870 -19839 16974 -19728
rect 8952 -20385 9133 -20129
rect 16510 -20503 16589 -20399
rect 16900 -20503 16974 -20400
rect 9972 -24875 10064 -24781
rect 12642 -24875 12734 -24781
rect 15308 -24875 15400 -24781
<< mimcap >>
rect -8656 48441 -3856 50174
rect -8656 46819 -8137 48441
rect -6873 46819 -3856 48441
rect -8656 45348 -3856 46819
rect -3076 48285 1724 50162
rect -3076 46823 -274 48285
rect 1121 46823 1724 48285
rect -3076 45342 1724 46823
rect 2424 48373 7224 50162
rect 2424 46911 5573 48373
rect 6968 46911 7224 48373
rect 2424 45342 7224 46911
rect 7924 48484 12724 50162
rect 7924 47022 10711 48484
rect 12106 47022 12724 48484
rect 7924 45342 12724 47022
rect 13424 48506 18224 50162
rect 13424 47044 16359 48506
rect 17754 47044 18224 48506
rect 13424 45342 18224 47044
rect 18924 48484 23724 50162
rect 18924 47022 21874 48484
rect 23269 47022 23724 48484
rect 18924 45342 23724 47022
rect 24424 48440 29224 50162
rect 24424 46978 24753 48440
rect 26148 46978 29224 48440
rect 24424 45342 29224 46978
rect -8656 42941 -3856 44674
rect -8656 41319 -8131 42941
rect -6873 41319 -3856 42941
rect -8656 39842 -3856 41319
rect -3076 42362 1724 44662
rect -3076 41284 -2580 42362
rect -1474 41284 1724 42362
rect -3076 39842 1724 41284
rect 2424 44000 7224 44662
rect 2424 43904 3174 44000
rect 2424 42386 4296 43904
rect 2424 42254 3174 42386
rect 4360 42254 7224 44000
rect 2424 39842 7224 42254
rect 7924 41646 12724 44662
rect 7924 40432 9000 41646
rect 10946 40432 12724 41646
rect 7924 39842 12724 40432
rect 13424 44296 18224 44662
rect 13424 42550 14250 44296
rect 15436 43970 18224 44296
rect 14316 42550 18224 43970
rect 13424 39842 18224 42550
rect 18924 42698 23724 44662
rect 18924 41748 19470 42698
rect 20756 41748 23724 42698
rect 18924 39842 23724 41748
rect 24424 41973 29224 44662
rect 24424 40511 24930 41973
rect 26325 40511 29224 41973
rect 24424 39842 29224 40511
rect -8656 37441 -3856 39162
rect -8656 35819 -8131 37441
rect -6873 35819 -3856 37441
rect -8656 34342 -3856 35819
rect -3076 38726 1724 39162
rect -3076 38662 -2464 38726
rect -3076 37208 -1308 38662
rect -3076 37144 -1342 37208
rect -1244 37144 1724 38726
rect -3076 36946 -2464 37144
rect -1278 36946 1724 37144
rect -3076 34342 1724 36946
rect 2424 38454 7224 39162
rect 2424 37104 3240 38454
rect 4206 37104 7224 38454
rect 2424 34342 7224 37104
rect 7924 38322 12724 39162
rect 7924 37108 8976 38322
rect 9076 37108 10618 38194
rect 10922 37108 12724 38322
rect 7924 34342 12724 37108
rect 13424 38682 18224 39162
rect 13424 37384 14362 38682
rect 15582 37384 18224 38682
rect 13424 34342 18224 37384
rect 18924 38956 23724 39162
rect 18924 37210 19888 38956
rect 21074 38826 23724 38956
rect 19954 37308 23724 38826
rect 21074 37210 23724 37308
rect 18924 34342 23724 37210
rect 24424 37344 29224 39162
rect 24424 35882 25019 37344
rect 26414 35882 29224 37344
rect 24424 34342 29224 35882
rect -8656 31941 -3856 33574
rect -8656 30319 -8131 31941
rect -6873 30319 -3856 31941
rect -8656 28748 -3856 30319
rect -3156 31941 1644 33574
rect -3156 30319 -2631 31941
rect -1373 30319 1644 31941
rect -3156 28748 1644 30319
rect 2344 31941 7144 33574
rect 2344 30319 2869 31941
rect 4127 30319 7144 31941
rect 2344 28748 7144 30319
rect 7844 31941 12644 33574
rect 7844 30319 8369 31941
rect 9627 30319 12644 31941
rect 7844 28748 12644 30319
rect 13344 31941 18144 33574
rect 13344 30319 13869 31941
rect 15127 30319 18144 31941
rect 13344 28748 18144 30319
rect 18844 31941 23644 33574
rect 18844 30319 19369 31941
rect 20627 30319 23644 31941
rect 18844 28748 23644 30319
rect 24344 31941 29144 33574
rect 24344 30319 24869 31941
rect 26127 30319 29144 31941
rect 24344 28748 29144 30319
<< mimcapcontact >>
rect -8137 46819 -6873 48441
rect -274 46823 1121 48285
rect 5573 46911 6968 48373
rect 10711 47022 12106 48484
rect 16359 47044 17754 48506
rect 21874 47022 23269 48484
rect 24753 46978 26148 48440
rect -8131 41319 -6873 42941
rect -2580 41284 -1474 42362
rect 3174 43904 4360 44000
rect 4296 42386 4360 43904
rect 3174 42254 4360 42386
rect 9000 40432 10946 41646
rect 14250 43970 15436 44296
rect 14250 42550 14316 43970
rect 19470 41748 20756 42698
rect 24930 40511 26325 41973
rect -8131 35819 -6873 37441
rect -2464 38662 -1244 38726
rect -1308 37208 -1244 38662
rect -1342 37144 -1244 37208
rect -2464 36946 -1278 37144
rect 3240 37104 4206 38454
rect 8976 38194 10922 38322
rect 8976 37108 9076 38194
rect 10618 37108 10922 38194
rect 14362 37384 15582 38682
rect 19888 38826 21074 38956
rect 19888 37308 19954 38826
rect 19888 37210 21074 37308
rect 25019 35882 26414 37344
rect -8131 30319 -6873 31941
rect -2631 30319 -1373 31941
rect 2869 30319 4127 31941
rect 8369 30319 9627 31941
rect 13869 30319 15127 31941
rect 19369 30319 20627 31941
rect 24869 30319 26127 31941
<< metal4 >>
rect -19220 56190 -17382 56450
rect -19220 55462 -18978 56190
rect -17592 55462 -17382 56190
rect -19220 55220 -17382 55462
rect -15220 56190 -13382 56450
rect -15220 55462 -14978 56190
rect -13592 55462 -13382 56190
rect -15220 55220 -13382 55462
rect -11220 56190 -9382 56450
rect -11220 55462 -10978 56190
rect -9592 55462 -9382 56190
rect -11220 55220 -9382 55462
rect -7220 56190 -5382 56450
rect -7220 55462 -6978 56190
rect -5592 55462 -5382 56190
rect -7220 55220 -5382 55462
rect -3220 56190 -1382 56450
rect -3220 55462 -2978 56190
rect -1592 55462 -1382 56190
rect -3220 55220 -1382 55462
rect 780 56190 2618 56450
rect 780 55462 1022 56190
rect 2408 55462 2618 56190
rect 780 55220 2618 55462
rect 4780 56190 6618 56450
rect 4780 55462 5022 56190
rect 6408 55462 6618 56190
rect 4780 55220 6618 55462
rect 8780 56190 10618 56450
rect 8780 55462 9022 56190
rect 10408 55462 10618 56190
rect 8780 55220 10618 55462
rect 12780 56190 14618 56450
rect 12780 55462 13022 56190
rect 14408 55462 14618 56190
rect 12780 55220 14618 55462
rect 16780 56190 18618 56450
rect 16780 55462 17022 56190
rect 18408 55462 18618 56190
rect 16780 55220 18618 55462
rect 20780 56190 22618 56450
rect 20780 55462 21022 56190
rect 22408 55462 22618 56190
rect 20780 55220 22618 55462
rect 24780 56190 26618 56450
rect 24780 55462 25022 56190
rect 26408 55462 26618 56190
rect 24780 55220 26618 55462
rect 28780 56190 30618 56450
rect 28780 55462 29022 56190
rect 30408 55462 30618 56190
rect 28780 55220 30618 55462
rect 32780 56190 34618 56450
rect 32780 55462 33022 56190
rect 34408 55462 34618 56190
rect 32780 55220 34618 55462
rect 36780 56190 38618 56450
rect 36780 55462 37022 56190
rect 38408 55462 38618 56190
rect 36780 55220 38618 55462
rect -20956 54026 -19118 54286
rect -20956 53298 -20714 54026
rect -19328 53298 -19118 54026
rect 28580 53656 35702 53680
rect -20956 53056 -19118 53298
rect 18990 53560 35702 53656
rect 18990 52822 19194 53560
rect 20672 52822 35702 53560
rect 18990 52656 35702 52822
rect 18990 52612 29220 52656
rect 32022 52564 35702 52656
rect 36822 52988 38660 53256
rect -11932 52000 -10624 52046
rect -11996 51779 4616 52000
rect -11996 51141 3367 51779
rect 4136 51141 4616 51779
rect -11996 50690 4616 51141
rect -20956 50026 -19118 50286
rect -20956 49298 -20714 50026
rect -19328 49298 -19118 50026
rect -20956 49056 -19118 49298
rect -20956 46026 -19118 46286
rect -20956 45298 -20714 46026
rect -19328 45298 -19118 46026
rect -20956 45056 -19118 45298
rect -20956 42026 -19118 42286
rect -20956 41298 -20714 42026
rect -19328 41298 -19118 42026
rect -20956 41056 -19118 41298
rect -20956 38026 -19118 38286
rect -20956 37298 -20714 38026
rect -19328 37298 -19118 38026
rect -20956 37056 -19118 37298
rect -11932 36624 -10624 50690
rect -11932 36390 -11578 36624
rect -11378 36390 -10624 36624
rect -20956 34026 -19118 34286
rect -20956 33298 -20714 34026
rect -19328 33298 -19118 34026
rect -20956 33056 -19118 33298
rect -20956 30026 -19118 30286
rect -20956 29298 -20714 30026
rect -19328 29298 -19118 30026
rect -20956 29056 -19118 29298
rect -20956 26026 -19118 26286
rect -20956 25298 -20714 26026
rect -19328 25298 -19118 26026
rect -20956 25056 -19118 25298
rect -11932 25128 -10624 36390
rect -8336 48806 -6680 48839
rect -8336 48773 26403 48806
rect -8336 48506 26469 48773
rect -8336 48484 16359 48506
rect -8336 48441 10711 48484
rect -8336 46819 -8137 48441
rect -6873 48373 10711 48441
rect -6873 48285 5573 48373
rect -6873 46823 -274 48285
rect 1121 46911 5573 48285
rect 6968 47022 10711 48373
rect 12106 47044 16359 48484
rect 17754 48484 26469 48506
rect 17754 47044 21874 48484
rect 12106 47022 21874 47044
rect 23269 48440 26469 48484
rect 23269 47022 24753 48440
rect 6968 46978 24753 47022
rect 26148 46978 26469 48440
rect 6968 46911 26469 46978
rect 1121 46823 26469 46911
rect -6873 46819 26469 46823
rect -8336 46554 26469 46819
rect -8336 42941 -6680 46554
rect -8336 41319 -8131 42941
rect -6873 41319 -6680 42941
rect -8336 37441 -6680 41319
rect -2888 43984 -1038 44446
rect 3048 44170 4531 44431
rect -2888 42878 -2504 43984
rect -1502 42878 -1038 43984
rect -2888 42362 -1038 42878
rect -2888 41284 -2580 42362
rect -1474 41284 -1038 42362
rect 2960 44000 4531 44170
rect 2960 43904 3174 44000
rect 2960 42386 3108 43904
rect 2960 42254 3174 42386
rect 4360 42254 4531 44000
rect 2960 41872 4531 42254
rect 14096 44296 15579 44373
rect 14096 42550 14250 44296
rect 15436 43970 15579 44296
rect 14096 42452 14316 42550
rect 15504 42452 15579 43970
rect 2960 41611 4443 41872
rect 8710 41646 11352 41912
rect 14096 41814 15579 42452
rect 19136 44164 21012 44678
rect 19136 43366 19702 44164
rect 20446 43366 21012 44164
rect 19136 42698 21012 43366
rect -2888 41054 -1038 41284
rect 8710 40432 9000 41646
rect 10946 40432 11352 41646
rect 19136 41748 19470 42698
rect 20756 41748 21012 42698
rect 19136 41130 21012 41748
rect 24648 41973 26469 46554
rect 8710 39640 11352 40432
rect 24648 40511 24930 41973
rect 26325 40511 26469 41973
rect 8710 39256 11198 39640
rect -8336 35819 -8131 37441
rect -6873 35819 -6680 37441
rect -3024 38726 -650 39156
rect 8710 38968 11352 39256
rect -3024 38662 -2464 38726
rect -3024 37144 -2496 38662
rect -1244 37144 -650 38726
rect -3024 36946 -2464 37144
rect -1278 36946 -650 37144
rect 2984 38454 4766 38936
rect 8710 38790 11176 38968
rect 2984 37104 3240 38454
rect 4206 37104 4766 38454
rect -2651 36377 -1168 36946
rect 2984 36874 4766 37104
rect 2934 36774 4766 36874
rect 8658 38322 11176 38790
rect 8658 37108 8976 38322
rect 8658 36868 9076 37108
rect 10922 37108 11176 38322
rect 10618 36868 11176 37108
rect -8336 32281 -6680 35819
rect 2934 35858 4716 36774
rect 8658 36470 11176 36868
rect 14004 38682 15990 38962
rect 14004 37384 14362 38682
rect 15582 37384 15990 38682
rect 2934 34966 3392 35858
rect 4054 34966 4716 35858
rect 2934 34712 4716 34966
rect 14004 36088 15990 37384
rect 19492 38956 21866 38990
rect 19492 37210 19888 38956
rect 21074 38826 21866 38956
rect 21142 37308 21866 38826
rect 21074 37210 21866 37308
rect 19492 36780 21866 37210
rect 24648 37344 26469 40511
rect 19766 36319 21249 36780
rect 14004 35196 14336 36088
rect 14998 35196 15990 36088
rect 14004 34916 15990 35196
rect 24648 35882 25019 37344
rect 26414 35882 26469 37344
rect 24648 32281 26469 35882
rect -8402 31941 26634 32281
rect -8402 30319 -8131 31941
rect -6873 30319 -2631 31941
rect -1373 30319 2869 31941
rect 4127 30319 8369 31941
rect 9627 30319 13869 31941
rect 15127 30319 19369 31941
rect 20627 30319 24869 31941
rect 26127 30319 26634 31941
rect -8402 29930 26634 30319
rect -8402 27902 -6746 29930
rect 24648 29830 26469 29930
rect 8960 28300 9880 28336
rect 8960 28064 9172 28300
rect 9526 28064 9880 28300
rect 8960 28032 9880 28064
rect -8402 27104 -8174 27902
rect -6984 27104 -6746 27902
rect -8402 26890 -6746 27104
rect 2998 27028 4580 27260
rect 2998 25912 3278 27028
rect 4440 25912 4580 27028
rect 2998 25540 4580 25912
rect -12226 23460 -10522 25128
rect -4056 23906 -946 24186
rect -4056 23460 -2162 23906
rect -12226 22970 -2162 23460
rect -1134 22970 -946 23906
rect -12226 22738 -946 22970
rect -20956 22026 -19118 22286
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -96266 13740 -95320 15274
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -96266 4182 -95320 5274
rect -27834 19740 -26806 21200
rect -20956 21298 -20714 22026
rect -19328 21298 -19118 22026
rect -12226 21628 -10522 22738
rect -20956 21056 -19118 21298
rect 2998 20656 4486 25540
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -27834 17740 -26806 19274
rect 2812 19308 4486 20656
rect 33324 19308 35650 52564
rect 36822 52260 37064 52988
rect 38450 52260 38660 52988
rect 36822 52018 38660 52260
rect 36822 48988 38660 49256
rect 36822 48260 37064 48988
rect 38450 48260 38660 48988
rect 36822 48018 38660 48260
rect 36822 44988 38660 45256
rect 36822 44260 37064 44988
rect 38450 44260 38660 44988
rect 36822 44018 38660 44260
rect 36822 40988 38660 41256
rect 36822 40260 37064 40988
rect 38450 40260 38660 40988
rect 36822 40018 38660 40260
rect 36822 36988 38660 37256
rect 36822 36260 37064 36988
rect 38450 36260 38660 36988
rect 36822 36018 38660 36260
rect 36822 32988 38660 33256
rect 36822 32260 37064 32988
rect 38450 32260 38660 32988
rect 36822 32018 38660 32260
rect 36822 28988 38660 29256
rect 36822 28260 37064 28988
rect 38450 28260 38660 28988
rect 36822 28018 38660 28260
rect 36822 24988 38660 25256
rect 36822 24260 37064 24988
rect 38450 24260 38660 24988
rect 36822 24018 38660 24260
rect 36822 20988 38660 21256
rect 36822 20260 37064 20988
rect 38450 20260 38660 20988
rect 36822 20018 38660 20260
rect 2812 18404 35650 19308
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -27834 15740 -26806 17274
rect -20956 18026 -19118 18286
rect -20956 17298 -20714 18026
rect -19328 17298 -19118 18026
rect 2812 18134 13138 18404
rect 13424 18134 35650 18404
rect 2812 17632 35650 18134
rect 33324 17494 35650 17632
rect -20956 17056 -19118 17298
rect 36822 16988 38660 17256
rect 36822 16260 37064 16988
rect 38450 16260 38660 16988
rect 36822 16018 38660 16260
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -27834 13740 -26806 15274
rect -18294 14908 -16456 15184
rect -18294 14180 -18052 14908
rect -16666 14180 -16456 14908
rect -18294 13938 -16456 14180
rect -14294 15084 -14106 15180
rect -13566 15084 -12456 15180
rect -14294 14908 -12456 15084
rect -14294 14180 -14052 14908
rect -12666 14180 -12456 14908
rect -14294 13938 -12456 14180
rect -10294 14908 -8456 15180
rect -10294 14180 -10052 14908
rect -8666 14180 -8456 14908
rect -10294 13938 -8456 14180
rect -6294 14908 -4456 15180
rect -6294 14180 -6052 14908
rect -4666 14180 -4456 14908
rect -6294 13938 -4456 14180
rect -2294 14908 -456 15180
rect -2294 14180 -2052 14908
rect -666 14180 -456 14908
rect -2294 13938 -456 14180
rect 1706 14908 3544 15180
rect 1706 14180 1948 14908
rect 3334 14180 3544 14908
rect 1706 13938 3544 14180
rect 5706 14908 7544 15180
rect 5706 14180 5948 14908
rect 7334 14180 7544 14908
rect 5706 13938 7544 14180
rect 9706 14908 11544 15180
rect 9706 14180 9948 14908
rect 11334 14180 11544 14908
rect 9706 13938 11544 14180
rect 13706 14908 15544 15180
rect 13706 14180 13948 14908
rect 15334 14180 15544 14908
rect 13706 13938 15544 14180
rect 17706 14908 19544 15180
rect 17706 14180 17948 14908
rect 19334 14180 19544 14908
rect 17706 13938 19544 14180
rect 21706 14908 23544 15180
rect 21706 14180 21948 14908
rect 23334 14180 23544 14908
rect 21706 13938 23544 14180
rect 25706 14908 27544 15180
rect 25706 14180 25948 14908
rect 27334 14180 27544 14908
rect 25706 13938 27544 14180
rect 29706 14908 31544 15180
rect 29706 14180 29948 14908
rect 31334 14180 31544 14908
rect 29706 13938 31544 14180
rect 33706 14908 35544 15180
rect 33706 14180 33948 14908
rect 35334 14180 35544 14908
rect 33706 13938 35544 14180
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -27834 11740 -26806 13274
rect 17792 12068 19104 12262
rect 17792 11828 18000 12068
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect 17786 11574 18000 11828
rect 18960 11574 19104 12068
rect 17786 11534 19104 11574
rect 17792 11354 19104 11534
rect -27834 9740 -26806 11274
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect -27834 7740 -26806 9274
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -27834 5740 -26806 7274
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6016 1794 6112
rect 1280 5776 1374 6016
rect 1700 5776 1794 6016
rect 1280 5678 1794 5776
rect 6168 6094 6682 6190
rect 6168 5854 6262 6094
rect 6588 5854 6682 6094
rect 6168 5756 6682 5854
rect 11480 5882 11994 5978
rect 11480 5642 11574 5882
rect 11900 5642 11994 5882
rect 11480 5544 11994 5642
rect 16916 5824 17430 5920
rect 16916 5584 17010 5824
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect -96266 4178 -95322 4182
rect -96396 3910 -95322 4178
rect -96396 3740 -62544 3910
rect -27834 3846 -26806 5274
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -96396 2966 -62544 3274
rect -60278 3740 -26756 3846
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect -60278 3224 -26756 3274
rect -61896 2890 -61292 2894
rect -61896 2826 -61864 2890
rect -61800 2826 -61464 2890
rect -61400 2826 -61292 2890
rect -61896 2812 -61292 2826
rect 18322 2026 18670 11354
rect 26106 3638 26596 3676
rect 26106 3246 26138 3638
rect 26538 3246 26596 3638
rect 26106 3216 26596 3246
rect 32364 2206 32976 2274
rect 3316 1698 4628 1892
rect 17370 1832 18682 2026
rect 3316 1204 3524 1698
rect 4484 1592 4628 1698
rect 10738 1592 12050 1708
rect 17370 1592 17578 1832
rect 4484 1514 17578 1592
rect 4484 1298 10946 1514
rect 4484 1204 4628 1298
rect 3316 984 4628 1204
rect 10738 1020 10946 1298
rect 11906 1338 17578 1514
rect 18538 1338 18682 1832
rect 32364 1746 32424 2206
rect 32904 1746 32976 2206
rect 32364 1676 32976 1746
rect 11906 1298 18682 1338
rect 11906 1020 12050 1298
rect 17370 1118 18682 1298
rect 10738 800 12050 1020
rect 8984 -8654 9262 -8635
rect 8984 -8967 9002 -8654
rect 9241 -8967 9262 -8654
rect 8984 -8986 9262 -8967
rect 16394 -8656 16700 -8641
rect 16394 -9006 16412 -8656
rect 16685 -9006 16700 -8656
rect 16394 -9018 16700 -9006
rect 5173 -12769 10124 -12730
rect 5173 -13742 5237 -12769
rect 7037 -13109 10124 -12769
rect 7037 -13140 10452 -13109
rect 15135 -13140 20792 -13136
rect 7037 -13161 20792 -13140
rect 7037 -13267 9970 -13161
rect 10076 -13267 12634 -13161
rect 12740 -13267 15296 -13161
rect 15402 -13267 20792 -13161
rect 7037 -13305 20792 -13267
rect 7037 -13327 18999 -13305
rect 7037 -13333 10452 -13327
rect 7037 -13742 10124 -13333
rect 12616 -13552 12760 -13327
rect 5173 -13875 10124 -13742
rect 5173 -13880 10129 -13875
rect 8935 -14220 9259 -14190
rect 8935 -14525 8991 -14220
rect 9227 -14525 9259 -14220
rect 8935 -14550 9259 -14525
rect 8951 -14557 9229 -14550
rect 9942 -15040 10129 -13880
rect 12611 -15020 12765 -13552
rect 15135 -14098 18999 -13327
rect 20398 -14098 20792 -13305
rect 15135 -14178 20792 -14098
rect 15137 -14367 20792 -14178
rect 15137 -14451 16245 -14367
rect 15137 -15016 16143 -14451
rect 9942 -18852 10096 -15040
rect 12616 -18852 12760 -15020
rect 15285 -17370 15429 -15016
rect 15285 -17618 15430 -17370
rect 15285 -18852 15429 -17618
rect 9876 -18880 15431 -18852
rect 9876 -18986 9964 -18880
rect 10070 -18885 15431 -18880
rect 10070 -18979 12640 -18885
rect 12732 -18979 15306 -18885
rect 15398 -18979 15431 -18885
rect 10070 -18986 15431 -18979
rect 9876 -19039 15431 -18986
rect 8913 -20129 9211 -20096
rect 8913 -20132 8952 -20129
rect 9133 -20132 9211 -20129
rect 8913 -20406 8947 -20132
rect 9183 -20406 9211 -20132
rect 8913 -20436 9211 -20406
rect 9942 -24744 10096 -19039
rect 12616 -24744 12760 -19039
rect 15285 -20387 15429 -19039
rect 16191 -19558 16520 -19538
rect 16191 -19916 16220 -19558
rect 16484 -19916 16520 -19558
rect 16191 -19931 16520 -19916
rect 15285 -20399 16995 -20387
rect 15285 -20503 16510 -20399
rect 16589 -20400 16995 -20399
rect 16589 -20503 16900 -20400
rect 16974 -20503 16995 -20400
rect 15285 -20520 16995 -20503
rect 15285 -24744 15429 -20520
rect 9888 -24781 15443 -24744
rect 9888 -24875 9972 -24781
rect 10064 -24875 12642 -24781
rect 12734 -24875 15308 -24781
rect 15400 -24875 15443 -24781
rect 9888 -24931 15443 -24875
rect 9942 -24933 10096 -24931
<< via4 >>
rect 19194 52822 20672 53560
rect 3367 51141 4136 51779
rect -2504 42878 -1502 43984
rect 3108 42386 4296 43904
rect 14316 42452 15504 43970
rect 19702 43366 20446 44164
rect -2496 37208 -1308 38662
rect -2496 37144 -1342 37208
rect 9076 36868 10618 38194
rect 3392 34966 4054 35858
rect 19954 37308 21142 38826
rect 14336 35196 14998 36088
rect 9172 28258 9526 28300
rect 9172 28064 9526 28258
rect 3278 25912 4440 27028
rect -2162 22970 -1134 23906
rect -96044 21274 -95512 21740
rect -94044 21274 -93512 21740
rect -92044 21274 -91512 21740
rect -90044 21274 -89512 21740
rect -88044 21274 -87512 21740
rect -86044 21274 -85512 21740
rect -84044 21274 -83512 21740
rect -82044 21274 -81512 21740
rect -80044 21274 -79512 21740
rect -78044 21274 -77512 21740
rect -76044 21274 -75512 21740
rect -74044 21274 -73512 21740
rect -72044 21274 -71512 21740
rect -70044 21274 -69512 21740
rect -68044 21274 -67512 21740
rect -66044 21274 -65512 21740
rect -64044 21274 -63512 21740
rect -62044 21274 -61512 21740
rect -60044 21274 -59512 21740
rect -58044 21274 -57512 21740
rect -56044 21274 -55512 21740
rect -54044 21274 -53512 21740
rect -52044 21274 -51512 21740
rect -50044 21274 -49512 21740
rect -48044 21274 -47512 21740
rect -46044 21274 -45512 21740
rect -44044 21274 -43512 21740
rect -42044 21274 -41512 21740
rect -40044 21274 -39512 21740
rect -38044 21274 -37512 21740
rect -36044 21274 -35512 21740
rect -34044 21274 -33512 21740
rect -32044 21274 -31512 21740
rect -30044 21274 -29512 21740
rect -27644 21274 -27112 21740
rect -96044 19274 -95512 19740
rect -96044 17274 -95512 17740
rect -96044 15274 -95512 15740
rect -96044 13274 -95512 13740
rect -96044 11274 -95512 11740
rect -96044 9274 -95512 9740
rect -96044 7274 -95512 7740
rect -96044 5274 -95512 5740
rect -27644 19274 -27112 19740
rect -27644 17274 -27112 17740
rect -27644 15274 -27112 15740
rect -27644 13274 -27112 13740
rect -27644 11274 -27112 11740
rect -27644 9274 -27112 9740
rect -27644 7274 -27112 7740
rect -27644 5274 -27112 5740
rect 1374 5776 1700 6016
rect 6262 5854 6588 6094
rect 11574 5642 11900 5882
rect 17010 5584 17336 5824
rect -95644 3274 -95112 3740
rect -93644 3274 -93112 3740
rect -91644 3274 -91112 3740
rect -89644 3274 -89112 3740
rect -87644 3274 -87112 3740
rect -85644 3274 -85112 3740
rect -83644 3274 -83112 3740
rect -81644 3274 -81112 3740
rect -79644 3274 -79112 3740
rect -77644 3274 -77112 3740
rect -75644 3274 -75112 3740
rect -73644 3274 -73112 3740
rect -71644 3274 -71112 3740
rect -69644 3274 -69112 3740
rect -67644 3274 -67112 3740
rect -65644 3274 -65112 3740
rect -63644 3274 -63112 3740
rect -59644 3274 -59112 3740
rect -57644 3274 -57112 3740
rect -55644 3274 -55112 3740
rect -53644 3274 -53112 3740
rect -51644 3274 -51112 3740
rect -49644 3274 -49112 3740
rect -47644 3274 -47112 3740
rect -45644 3274 -45112 3740
rect -43644 3274 -43112 3740
rect -41644 3274 -41112 3740
rect -39644 3274 -39112 3740
rect -37644 3274 -37112 3740
rect -35644 3274 -35112 3740
rect -33644 3274 -33112 3740
rect -31644 3274 -31112 3740
rect -29644 3274 -29112 3740
rect -27644 3274 -27112 3740
rect 9002 -8967 9241 -8654
rect 16412 -9006 16685 -8656
rect 8991 -14525 9174 -14220
rect 9174 -14525 9227 -14220
rect 8947 -20385 8952 -20132
rect 8952 -20385 9133 -20132
rect 9133 -20385 9183 -20132
rect 8947 -20406 9183 -20385
rect 16220 -19562 16484 -19558
rect 16220 -19911 16230 -19562
rect 16230 -19911 16476 -19562
rect 16476 -19911 16484 -19562
rect 16220 -19916 16484 -19911
rect 16846 -19728 17083 -19624
rect 16846 -19839 16870 -19728
rect 16870 -19839 16974 -19728
rect 16974 -19839 17083 -19728
rect 16846 -19862 17083 -19839
<< metal5 >>
rect -2626 53560 20854 53816
rect -2626 52822 19194 53560
rect 20672 52850 20854 53560
rect 20672 52822 20882 52850
rect -2626 52442 20882 52822
rect -2592 45062 -1290 52442
rect 3040 51846 15292 52024
rect 3040 51779 15472 51846
rect 3040 51141 3367 51779
rect 4136 51141 15472 51779
rect 3040 50966 15472 51141
rect 3124 50944 4488 50966
rect -2734 43984 -1168 45062
rect 3124 44431 4316 50944
rect 3048 44258 4531 44431
rect 14280 44373 15472 50966
rect 19580 46914 20882 52442
rect 19136 46580 20882 46914
rect -2734 42878 -2504 43984
rect -1502 42878 -1168 43984
rect -2734 42544 -1168 42878
rect 2890 43904 4702 44258
rect 2890 42386 3108 43904
rect 4296 42386 4702 43904
rect 2890 42284 4702 42386
rect 14096 43970 15579 44373
rect 14096 42452 14316 43970
rect 15504 42452 15579 43970
rect 19136 44164 20832 46580
rect 19136 43366 19702 44164
rect 20446 43366 20832 44164
rect 19136 43186 20832 43366
rect 3048 41872 4531 42284
rect 14096 41814 15579 42452
rect -2651 38906 -1168 38936
rect -2812 38662 -1000 38906
rect -2812 37144 -2496 38662
rect -1308 37208 -1000 38662
rect 19732 38826 21544 39064
rect -1342 37144 -1000 37208
rect -2812 36932 -1000 37144
rect 8684 38194 10720 38448
rect -2651 36377 -1168 36932
rect 8684 36868 9076 38194
rect 10618 36868 10720 38194
rect 19732 37308 19954 38826
rect 21142 37308 21544 38826
rect 19732 37090 21544 37308
rect -2602 26346 -1182 36377
rect 8684 36256 10720 36868
rect 19766 36638 21249 37090
rect 19754 36319 21249 36638
rect 3170 35858 4384 35990
rect 8684 35882 10264 36256
rect 3170 34966 3392 35858
rect 4054 34966 4384 35858
rect 8672 35256 10264 35882
rect 14136 36088 15396 36270
rect 3170 27404 4384 34966
rect 8734 28406 10174 35256
rect 14136 35216 14336 36088
rect 14166 35196 14336 35216
rect 14998 35216 15396 36088
rect 14998 35196 15380 35216
rect 8722 28300 10184 28406
rect 8722 28064 9172 28300
rect 9526 28064 10184 28300
rect 8722 27962 10184 28064
rect 14166 27404 15380 35196
rect 3102 27028 15426 27404
rect -2602 25412 -1168 26346
rect 3102 25912 3278 27028
rect 4440 25912 15426 27028
rect 3102 25526 15426 25912
rect 19754 25682 21174 36319
rect -2570 24210 -1168 25412
rect 19728 25458 21174 25682
rect 19728 24210 21130 25458
rect -2570 23906 21246 24210
rect -2570 22970 -2162 23906
rect -1134 22970 21246 23906
rect -2570 22944 21246 22970
rect -2524 22898 21246 22944
rect 19728 22876 21130 22898
rect -96266 21946 -94632 21968
rect -96266 21906 -26824 21946
rect -96266 21740 -26806 21906
rect -96266 21274 -96044 21740
rect -95512 21274 -94044 21740
rect -93512 21274 -92044 21740
rect -91512 21274 -90044 21740
rect -89512 21274 -88044 21740
rect -87512 21274 -86044 21740
rect -85512 21274 -84044 21740
rect -83512 21274 -82044 21740
rect -81512 21274 -80044 21740
rect -79512 21274 -78044 21740
rect -77512 21274 -76044 21740
rect -75512 21274 -74044 21740
rect -73512 21274 -72044 21740
rect -71512 21274 -70044 21740
rect -69512 21274 -68044 21740
rect -67512 21274 -66044 21740
rect -65512 21274 -64044 21740
rect -63512 21274 -62044 21740
rect -61512 21274 -60044 21740
rect -59512 21274 -58044 21740
rect -57512 21274 -56044 21740
rect -55512 21274 -54044 21740
rect -53512 21274 -52044 21740
rect -51512 21274 -50044 21740
rect -49512 21274 -48044 21740
rect -47512 21274 -46044 21740
rect -45512 21274 -44044 21740
rect -43512 21274 -42044 21740
rect -41512 21274 -40044 21740
rect -39512 21274 -38044 21740
rect -37512 21274 -36044 21740
rect -35512 21274 -34044 21740
rect -33512 21274 -32044 21740
rect -31512 21274 -30044 21740
rect -29512 21274 -27644 21740
rect -27112 21274 -26806 21740
rect -96266 21200 -26806 21274
rect -96266 21172 -94632 21200
rect -96266 21170 -95308 21172
rect -96266 19740 -95320 21170
rect -96266 19274 -96044 19740
rect -95512 19274 -95320 19740
rect -96266 17740 -95320 19274
rect -96266 17274 -96044 17740
rect -95512 17274 -95320 17740
rect -96266 15740 -95320 17274
rect -96266 15274 -96044 15740
rect -95512 15274 -95320 15740
rect -96266 13740 -95320 15274
rect -96266 13274 -96044 13740
rect -95512 13274 -95320 13740
rect -96266 11740 -95320 13274
rect -96266 11274 -96044 11740
rect -95512 11274 -95320 11740
rect -96266 9740 -95320 11274
rect -96266 9274 -96044 9740
rect -95512 9274 -95320 9740
rect -96266 7740 -95320 9274
rect -96266 7274 -96044 7740
rect -95512 7274 -95320 7740
rect -96266 5740 -95320 7274
rect -96266 5274 -96044 5740
rect -95512 5274 -95320 5740
rect -96266 4178 -95320 5274
rect -96396 3910 -95320 4178
rect -27834 19740 -26806 21200
rect -27834 19274 -27644 19740
rect -27112 19274 -26806 19740
rect -27834 17740 -26806 19274
rect -27834 17274 -27644 17740
rect -27112 17274 -26806 17740
rect -27834 15740 -26806 17274
rect -27834 15274 -27644 15740
rect -27112 15274 -26806 15740
rect -27834 13740 -26806 15274
rect -27834 13274 -27644 13740
rect -27112 13274 -26806 13740
rect -27834 11740 -26806 13274
rect -27834 11274 -27644 11740
rect -27112 11274 -26806 11740
rect -27834 9740 -26806 11274
rect -27834 9274 -27644 9740
rect -27112 9274 -26806 9740
rect -27834 7740 -26806 9274
rect -27834 7274 -27644 7740
rect -27112 7274 -26806 7740
rect -27834 5740 -26806 7274
rect -27834 5274 -27644 5740
rect -27112 5274 -26806 5740
rect 1280 6098 1794 6112
rect 6168 6098 6682 6190
rect 1280 6094 17234 6098
rect 1280 6016 6262 6094
rect 1280 5776 1374 6016
rect 1700 5854 6262 6016
rect 6588 5920 17234 6094
rect 6588 5882 17430 5920
rect 6588 5854 11574 5882
rect 1700 5776 11574 5854
rect 1280 5724 11574 5776
rect 1280 5678 1794 5724
rect 11480 5642 11574 5724
rect 11900 5824 17430 5882
rect 11900 5724 17010 5824
rect 11900 5642 11994 5724
rect 11480 5544 11994 5642
rect 16916 5584 17010 5724
rect 17336 5584 17430 5824
rect 16916 5486 17430 5584
rect -96396 3740 -62544 3910
rect -27834 3846 -26806 5274
rect -96396 3274 -95644 3740
rect -95112 3274 -93644 3740
rect -93112 3274 -91644 3740
rect -91112 3274 -89644 3740
rect -89112 3274 -87644 3740
rect -87112 3274 -85644 3740
rect -85112 3274 -83644 3740
rect -83112 3274 -81644 3740
rect -81112 3274 -79644 3740
rect -79112 3274 -77644 3740
rect -77112 3274 -75644 3740
rect -75112 3274 -73644 3740
rect -73112 3274 -71644 3740
rect -71112 3274 -69644 3740
rect -69112 3274 -67644 3740
rect -67112 3274 -65644 3740
rect -65112 3274 -63644 3740
rect -63112 3274 -62544 3740
rect -96396 2966 -62544 3274
rect -60278 3740 -26756 3846
rect -60278 3274 -59644 3740
rect -59112 3274 -57644 3740
rect -57112 3274 -55644 3740
rect -55112 3274 -53644 3740
rect -53112 3274 -51644 3740
rect -51112 3274 -49644 3740
rect -49112 3274 -47644 3740
rect -47112 3274 -45644 3740
rect -45112 3274 -43644 3740
rect -43112 3274 -41644 3740
rect -41112 3274 -39644 3740
rect -39112 3274 -37644 3740
rect -37112 3274 -35644 3740
rect -35112 3274 -33644 3740
rect -33112 3274 -31644 3740
rect -31112 3274 -29644 3740
rect -29112 3274 -27644 3740
rect -27112 3274 -26756 3740
rect -60278 3224 -26756 3274
rect 26106 3216 26596 3676
rect 8943 -8654 9310 -8619
rect 8943 -8967 9002 -8654
rect 9241 -8967 9310 -8654
rect 8943 -14199 9310 -8967
rect 8938 -14220 9310 -14199
rect 16360 -8656 16760 -8611
rect 16360 -9006 16412 -8656
rect 16685 -9006 16760 -8656
rect 16360 -11055 16760 -9006
rect 16360 -11375 18228 -11055
rect 16360 -14211 16760 -11375
rect 8938 -14525 8991 -14220
rect 9227 -14525 9310 -14220
rect 8938 -14527 9310 -14525
rect 8938 -19309 9312 -14527
rect 16208 -14626 16760 -14211
rect 8741 -19311 9320 -19309
rect 16208 -19311 16758 -14626
rect 8741 -19381 16758 -19311
rect 8741 -19558 17398 -19381
rect 8741 -19916 16220 -19558
rect 16484 -19624 17398 -19558
rect 16484 -19862 16846 -19624
rect 17083 -19862 17398 -19624
rect 16484 -19916 17398 -19862
rect 8741 -19990 17398 -19916
rect 8741 -19991 16758 -19990
rect 8741 -19998 16513 -19991
rect 17078 -19992 17398 -19990
rect 8741 -20097 9320 -19998
rect 8738 -20125 9320 -20097
rect 8738 -20132 9313 -20125
rect 8738 -20406 8947 -20132
rect 9183 -20406 9313 -20132
rect 8738 -20518 9313 -20406
rect 8938 -20519 9312 -20518
<< res0p35 >>
rect -16258 44520 -16184 49250
rect -15940 44520 -15866 49250
rect -15622 44520 -15548 49250
rect -15304 44520 -15230 49250
rect -16206 37242 -16132 41972
rect -15850 37224 -15776 41954
rect -15532 37224 -15458 41954
rect -15134 37206 -15060 41936
rect -16214 30742 -16140 35472
rect -15876 30762 -15802 35492
rect -15558 30762 -15484 35492
rect -15188 30760 -15114 35490
rect -16192 23990 -16118 28720
rect -15874 23990 -15800 28720
rect -15556 23990 -15482 28720
rect -15238 23990 -15164 28720
rect 554 10730 4408 10804
rect 5784 10730 9638 10804
rect 11014 10730 14868 10804
rect 16244 10730 20098 10804
rect 554 10410 4408 10484
rect 5784 10410 9638 10484
rect 11014 10410 14868 10484
rect 16244 10410 20098 10484
rect 554 10090 4408 10164
rect 5798 10068 9652 10142
rect 10994 10070 14848 10144
rect 16244 10090 20098 10164
rect 554 9770 4408 9844
rect 5798 9750 9652 9824
rect 10994 9752 14848 9826
rect 16244 9770 20098 9844
rect 554 9450 4408 9524
rect 5798 9432 9652 9506
rect 10994 9434 14848 9508
rect 16244 9450 20098 9524
rect 554 9130 4408 9204
rect 5798 9114 9652 9188
rect 10994 9116 14848 9190
rect 16244 9130 20098 9204
rect 554 8810 4408 8884
rect 5798 8796 9652 8870
rect 10994 8798 14848 8872
rect 16244 8810 20098 8884
rect 554 8490 4408 8564
rect 5798 8478 9652 8552
rect 10994 8480 14848 8554
rect 16244 8490 20098 8564
rect 554 8170 4408 8244
rect 5798 8160 9652 8234
rect 10994 8162 14848 8236
rect 16244 8170 20098 8244
rect 554 7850 4408 7924
rect 5798 7842 9652 7916
rect 10994 7844 14848 7918
rect 16244 7850 20098 7924
rect 554 7530 4408 7604
rect 5798 7524 9652 7598
rect 10994 7526 14848 7600
rect 16244 7530 20098 7604
rect 554 7210 4408 7284
rect 5818 7178 9672 7252
rect 11014 7208 14868 7282
rect 16244 7210 20098 7284
rect 554 6890 4408 6964
rect 5818 6858 9672 6932
rect 11014 6890 14868 6964
rect 16244 6890 20098 6964
<< labels >>
flabel metal4 17676 -13705 17676 -13705 0 FreeSans 1600 0 0 0 ring_changed_0/GND
flabel metal5 17698 -11225 17698 -11225 0 FreeSans 1600 0 0 0 ring_changed_0/VDD
flabel metal2 17378 -7765 17378 -7765 0 FreeSans 1600 0 0 0 ring_changed_0/Vinit
flabel metal2 8226 -7773 8226 -7773 0 FreeSans 1600 0 0 0 ring_changed_0/Vctrl
flabel metal1 17564 -20195 17564 -20195 0 FreeSans 1600 0 0 0 ring_changed_0/FvcoBUF
flabel metal1 16984 -20827 16984 -20827 0 FreeSans 1600 0 0 0 ring_changed_0/Fvco
flabel locali 11446 -9417 11446 -9417 0 FreeSans 1600 0 0 0 ring_changed_0/Vso1
flabel locali 14364 -9417 14364 -9417 0 FreeSans 1600 0 0 0 ring_changed_0/Vso2
flabel locali 16146 -9411 16146 -9411 0 FreeSans 1600 0 0 0 ring_changed_0/Vso3
flabel locali 10944 -21023 10944 -21023 0 FreeSans 1600 0 0 0 ring_changed_0/Vso7
flabel locali 14064 -21035 14064 -21035 0 FreeSans 1600 0 0 0 ring_changed_0/Vso8
flabel locali 12616 -7119 12616 -7119 0 FreeSans 1600 0 0 0 ring_changed_0/Vst
flabel locali 14698 -15115 14698 -15115 0 FreeSans 1600 0 0 0 ring_changed_0/Vso4
flabel locali 12166 -15141 12166 -15141 0 FreeSans 1600 0 0 0 ring_changed_0/Vso5
flabel locali 9580 -15101 9580 -15101 0 FreeSans 1600 0 0 0 ring_changed_0/Vso6
flabel locali -7677 -4636 -7643 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
flabel locali -9128 -4568 -9094 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/CLK
rlabel viali -7677 -4636 -7643 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel locali -7677 -4662 -7629 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel locali -7737 -4582 -7629 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -7689 -4642 -7631 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -7749 -4596 -7691 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -7749 -4605 -7631 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -8409 -4605 -8279 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -8409 -4633 -7631 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
rlabel metal1 -8409 -4642 -8279 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/RESET_B
flabel locali -7404 -4571 -7375 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/Q
flabel locali -7102 -4568 -7080 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/Q_N
flabel locali -9128 -4500 -9094 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/CLK
flabel locali -8853 -4500 -8819 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/D
rlabel viali -9129 -4262 -9095 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/VPWR
rlabel viali -9037 -4262 -9003 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/VPB
rlabel viali -9129 -4806 -9095 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/VGND
rlabel viali -9037 -4806 -9003 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[0]/VNB
flabel locali -5561 -4636 -5527 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
flabel locali -7012 -4568 -6978 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/CLK
rlabel viali -5561 -4636 -5527 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel locali -5561 -4662 -5513 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel locali -5621 -4582 -5513 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -5573 -4642 -5515 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -5633 -4596 -5575 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -5633 -4605 -5515 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -6293 -4605 -6163 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -6293 -4633 -5515 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
rlabel metal1 -6293 -4642 -6163 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/RESET_B
flabel locali -5288 -4571 -5259 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/Q
flabel locali -4986 -4568 -4964 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/Q_N
flabel locali -7012 -4500 -6978 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/CLK
flabel locali -6737 -4500 -6703 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/D
rlabel viali -7013 -4262 -6979 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/VPWR
rlabel viali -6921 -4262 -6887 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/VPB
rlabel viali -7013 -4806 -6979 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/VGND
rlabel viali -6921 -4806 -6887 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[1]/VNB
flabel locali -3445 -4636 -3411 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
flabel locali -4896 -4568 -4862 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/CLK
rlabel viali -3445 -4636 -3411 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel locali -3445 -4662 -3397 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel locali -3505 -4582 -3397 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -3457 -4642 -3399 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -3517 -4596 -3459 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -3517 -4605 -3399 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -4177 -4605 -4047 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -4177 -4633 -3399 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
rlabel metal1 -4177 -4642 -4047 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/RESET_B
flabel locali -3172 -4571 -3143 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/Q
flabel locali -2870 -4568 -2848 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/Q_N
flabel locali -4896 -4500 -4862 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/CLK
flabel locali -4621 -4500 -4587 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/D
rlabel viali -4897 -4262 -4863 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/VPWR
rlabel viali -4805 -4262 -4771 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/VPB
rlabel viali -4897 -4806 -4863 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/VGND
rlabel viali -4805 -4806 -4771 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[2]/VNB
flabel locali -1329 -4636 -1295 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
flabel locali -2780 -4568 -2746 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/CLK
rlabel viali -1329 -4636 -1295 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel locali -1329 -4662 -1281 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel locali -1389 -4582 -1281 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -1341 -4642 -1283 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -1401 -4596 -1343 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -1401 -4605 -1283 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -2061 -4605 -1931 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -2061 -4633 -1283 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
rlabel metal1 -2061 -4642 -1931 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/RESET_B
flabel locali -1056 -4571 -1027 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/Q
flabel locali -754 -4568 -732 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/Q_N
flabel locali -2780 -4500 -2746 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/CLK
flabel locali -2505 -4500 -2471 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/D
rlabel viali -2781 -4262 -2747 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/VPWR
rlabel viali -2689 -4262 -2655 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/VPB
rlabel viali -2781 -4806 -2747 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/VGND
rlabel viali -2689 -4806 -2655 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[3]/VNB
flabel locali 787 -4636 821 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
flabel locali -664 -4568 -630 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/CLK
rlabel viali 787 -4636 821 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel locali 787 -4662 835 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel locali 727 -4582 835 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 775 -4642 833 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 715 -4596 773 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 715 -4605 833 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 55 -4605 185 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 55 -4633 833 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
rlabel metal1 55 -4642 185 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/RESET_B
flabel locali 1060 -4571 1089 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/Q
flabel locali 1362 -4568 1384 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/Q_N
flabel locali -664 -4500 -630 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/CLK
flabel locali -389 -4500 -355 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/D
rlabel viali -665 -4262 -631 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/VPWR
rlabel viali -573 -4262 -539 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/VPB
rlabel viali -665 -4806 -631 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/VGND
rlabel viali -573 -4806 -539 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[4]/VNB
flabel locali 2903 -4636 2937 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
flabel locali 1452 -4568 1486 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/CLK
rlabel viali 2903 -4636 2937 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel locali 2903 -4662 2951 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel locali 2843 -4582 2951 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2891 -4642 2949 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2831 -4596 2889 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2831 -4605 2949 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2171 -4605 2301 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2171 -4633 2949 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
rlabel metal1 2171 -4642 2301 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/RESET_B
flabel locali 3176 -4571 3205 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/Q
flabel locali 3478 -4568 3500 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/Q_N
flabel locali 1452 -4500 1486 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/CLK
flabel locali 1727 -4500 1761 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/D
rlabel viali 1451 -4262 1485 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/VPWR
rlabel viali 1543 -4262 1577 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/VPB
rlabel viali 1451 -4806 1485 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/VGND
rlabel viali 1543 -4806 1577 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[5]/VNB
flabel locali 5019 -4636 5053 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
flabel locali 3568 -4568 3602 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/CLK
rlabel viali 5019 -4636 5053 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel locali 5019 -4662 5067 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel locali 4959 -4582 5067 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 5007 -4642 5065 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 4947 -4596 5005 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 4947 -4605 5065 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 4287 -4605 4417 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 4287 -4633 5065 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
rlabel metal1 4287 -4642 4417 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/RESET_B
flabel locali 5292 -4571 5321 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/Q
flabel locali 5594 -4568 5616 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/Q_N
flabel locali 3568 -4500 3602 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/CLK
flabel locali 3843 -4500 3877 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/D
rlabel viali 3567 -4262 3601 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/VPWR
rlabel viali 3659 -4262 3693 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/VPB
rlabel viali 3567 -4806 3601 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/VGND
rlabel viali 3659 -4806 3693 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[6]/VNB
flabel locali 7135 -4636 7169 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
flabel locali 5684 -4568 5718 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/CLK
rlabel viali 7135 -4636 7169 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel locali 7135 -4662 7183 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel locali 7075 -4582 7183 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 7123 -4642 7181 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 7063 -4596 7121 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 7063 -4605 7181 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 6403 -4605 6533 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 6403 -4633 7181 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
rlabel metal1 6403 -4642 6533 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/RESET_B
flabel locali 7408 -4571 7437 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/Q
flabel locali 7710 -4568 7732 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/Q_N
flabel locali 5684 -4500 5718 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/CLK
flabel locali 5959 -4500 5993 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/D
rlabel viali 5683 -4262 5717 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/VPWR
rlabel viali 5775 -4262 5809 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/VPB
rlabel viali 5683 -4806 5717 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/VGND
rlabel viali 5775 -4806 5809 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[7]/VNB
flabel locali 9251 -4636 9285 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
flabel locali 7800 -4568 7834 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/CLK
rlabel viali 9251 -4636 9285 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel locali 9251 -4662 9299 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel locali 9191 -4582 9299 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 9239 -4642 9297 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 9179 -4596 9237 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 9179 -4605 9297 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 8519 -4605 8649 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 8519 -4633 9297 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
rlabel metal1 8519 -4642 8649 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/RESET_B
flabel locali 9524 -4571 9553 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/Q
flabel locali 9826 -4568 9848 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/Q_N
flabel locali 7800 -4500 7834 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/CLK
flabel locali 8075 -4500 8109 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/D
rlabel viali 7799 -4262 7833 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/VPWR
rlabel viali 7891 -4262 7925 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/VPB
rlabel viali 7799 -4806 7833 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/VGND
rlabel viali 7891 -4806 7925 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[8]/VNB
flabel locali 11367 -4636 11401 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
flabel locali 9916 -4568 9950 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/CLK
rlabel viali 11367 -4636 11401 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel locali 11367 -4662 11415 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel locali 11307 -4582 11415 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 11355 -4642 11413 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 11295 -4596 11353 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 11295 -4605 11413 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 10635 -4605 10765 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 10635 -4633 11413 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
rlabel metal1 10635 -4642 10765 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
flabel locali 11640 -4571 11669 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/Q
flabel locali 11942 -4568 11964 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/Q_N
flabel locali 9916 -4500 9950 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/CLK
flabel locali 10191 -4500 10225 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/D
rlabel viali 9915 -4262 9949 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/VPWR
rlabel viali 10007 -4262 10041 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/VPB
rlabel viali 9915 -4806 9949 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/VGND
rlabel viali 10007 -4806 10041 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[9]/VNB
flabel locali 13483 -4636 13517 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
flabel locali 12032 -4568 12066 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/CLK
rlabel viali 13483 -4636 13517 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel locali 13483 -4662 13531 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel locali 13423 -4582 13531 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 13471 -4642 13529 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 13411 -4596 13469 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 13411 -4605 13529 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 12751 -4605 12881 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 12751 -4633 13529 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
rlabel metal1 12751 -4642 12881 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/RESET_B
flabel locali 13756 -4571 13785 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/Q
flabel locali 14058 -4568 14080 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/Q_N
flabel locali 12032 -4500 12066 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/CLK
flabel locali 12307 -4500 12341 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/D
rlabel viali 12031 -4262 12065 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/VPWR
rlabel viali 12123 -4262 12157 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/VPB
rlabel viali 12031 -4806 12065 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/VGND
rlabel viali 12123 -4806 12157 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[10]/VNB
flabel locali 15599 -4636 15633 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
flabel locali 14148 -4568 14182 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/CLK
rlabel viali 15599 -4636 15633 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel locali 15599 -4662 15647 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel locali 15539 -4582 15647 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 15587 -4642 15645 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 15527 -4596 15585 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 15527 -4605 15645 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 14867 -4605 14997 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 14867 -4633 15645 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
rlabel metal1 14867 -4642 14997 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/RESET_B
flabel locali 15872 -4571 15901 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/Q
flabel locali 16174 -4568 16196 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/Q_N
flabel locali 14148 -4500 14182 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/CLK
flabel locali 14423 -4500 14457 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/D
rlabel viali 14147 -4262 14181 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/VPWR
rlabel viali 14239 -4262 14273 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/VPB
rlabel viali 14147 -4806 14181 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/VGND
rlabel viali 14239 -4806 14273 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[11]/VNB
flabel locali 17715 -4636 17749 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
flabel locali 16264 -4568 16298 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/CLK
rlabel viali 17715 -4636 17749 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel locali 17715 -4662 17763 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel locali 17655 -4582 17763 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 17703 -4642 17761 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 17643 -4596 17701 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 17643 -4605 17761 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 16983 -4605 17113 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 16983 -4633 17761 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
rlabel metal1 16983 -4642 17113 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/RESET_B
flabel locali 17988 -4571 18017 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/Q
flabel locali 18290 -4568 18312 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/Q_N
flabel locali 16264 -4500 16298 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/CLK
flabel locali 16539 -4500 16573 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/D
rlabel viali 16263 -4262 16297 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/VPWR
rlabel viali 16355 -4262 16389 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/VPB
rlabel viali 16263 -4806 16297 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/VGND
rlabel viali 16355 -4806 16389 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[12]/VNB
flabel locali 19831 -4636 19865 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
flabel locali 18380 -4568 18414 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/CLK
rlabel viali 19831 -4636 19865 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel locali 19831 -4662 19879 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel locali 19771 -4582 19879 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19819 -4642 19877 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19759 -4596 19817 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19759 -4605 19877 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19099 -4605 19229 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19099 -4633 19877 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
rlabel metal1 19099 -4642 19229 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/RESET_B
flabel locali 20104 -4571 20133 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/Q
flabel locali 20406 -4568 20428 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/Q_N
flabel locali 18380 -4500 18414 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/CLK
flabel locali 18655 -4500 18689 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/D
rlabel viali 18379 -4262 18413 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/VPWR
rlabel viali 18471 -4262 18505 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/VPB
rlabel viali 18379 -4806 18413 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/VGND
rlabel viali 18471 -4806 18505 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[13]/VNB
flabel locali 21947 -4636 21981 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
flabel locali 20496 -4568 20530 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/CLK
rlabel viali 21947 -4636 21981 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel locali 21947 -4662 21995 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel locali 21887 -4582 21995 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21935 -4642 21993 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21875 -4596 21933 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21875 -4605 21993 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21215 -4605 21345 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21215 -4633 21993 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
rlabel metal1 21215 -4642 21345 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/RESET_B
flabel locali 22220 -4571 22249 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/Q
flabel locali 22522 -4568 22544 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/Q_N
flabel locali 20496 -4500 20530 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/CLK
flabel locali 20771 -4500 20805 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/D
rlabel viali 20495 -4262 20529 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/VPWR
rlabel viali 20587 -4262 20621 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/VPB
rlabel viali 20495 -4806 20529 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/VGND
rlabel viali 20587 -4806 20621 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[14]/VNB
flabel locali 24063 -4636 24097 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
flabel locali 22612 -4568 22646 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/CLK
rlabel viali 24063 -4636 24097 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel locali 24063 -4662 24111 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel locali 24003 -4582 24111 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 24051 -4642 24109 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 23991 -4596 24049 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 23991 -4605 24109 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 23331 -4605 23461 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 23331 -4633 24109 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
rlabel metal1 23331 -4642 23461 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/RESET_B
flabel locali 24336 -4571 24365 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/Q
flabel locali 24638 -4568 24660 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/Q_N
flabel locali 22612 -4500 22646 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/CLK
flabel locali 22887 -4500 22921 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/D
rlabel viali 22611 -4262 22645 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/VPWR
rlabel viali 22703 -4262 22737 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/VPB
rlabel viali 22611 -4806 22645 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/VGND
rlabel viali 22703 -4806 22737 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[15]/VNB
flabel locali 26179 -4636 26213 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
flabel locali 24728 -4568 24762 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/CLK
rlabel viali 26179 -4636 26213 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel locali 26179 -4662 26227 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel locali 26119 -4582 26227 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 26167 -4642 26225 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 26107 -4596 26165 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 26107 -4605 26225 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 25447 -4605 25577 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 25447 -4633 26225 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
rlabel metal1 25447 -4642 25577 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/RESET_B
flabel locali 26452 -4571 26481 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/Q
flabel locali 26754 -4568 26776 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/Q_N
flabel locali 24728 -4500 24762 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/CLK
flabel locali 25003 -4500 25037 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/D
rlabel viali 24727 -4262 24761 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/VPWR
rlabel viali 24819 -4262 24853 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/VPB
rlabel viali 24727 -4806 24761 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/VGND
rlabel viali 24819 -4806 24853 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[16]/VNB
flabel locali 28295 -4636 28329 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
flabel locali 26844 -4568 26878 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/CLK
rlabel viali 28295 -4636 28329 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel locali 28295 -4662 28343 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel locali 28235 -4582 28343 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 28283 -4642 28341 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 28223 -4596 28281 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 28223 -4605 28341 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 27563 -4605 27693 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 27563 -4633 28341 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
rlabel metal1 27563 -4642 27693 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/RESET_B
flabel locali 28568 -4571 28597 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/Q
flabel locali 28870 -4568 28892 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/Q_N
flabel locali 26844 -4500 26878 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/CLK
flabel locali 27119 -4500 27153 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/D
rlabel viali 26843 -4262 26877 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/VPWR
rlabel viali 26935 -4262 26969 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/VPB
rlabel viali 26843 -4806 26877 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/VGND
rlabel viali 26935 -4806 26969 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[17]/VNB
flabel locali 30411 -4636 30445 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
flabel locali 28960 -4568 28994 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/CLK
rlabel viali 30411 -4636 30445 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel locali 30411 -4662 30459 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel locali 30351 -4582 30459 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 30399 -4642 30457 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 30339 -4596 30397 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 30339 -4605 30457 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 29679 -4605 29809 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 29679 -4633 30457 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
rlabel metal1 29679 -4642 29809 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/RESET_B
flabel locali 30684 -4571 30713 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/Q
flabel locali 30986 -4568 31008 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/Q_N
flabel locali 28960 -4500 28994 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/CLK
flabel locali 29235 -4500 29269 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/D
rlabel viali 28959 -4262 28993 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/VPWR
rlabel viali 29051 -4262 29085 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/VPB
rlabel viali 28959 -4806 28993 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/VGND
rlabel viali 29051 -4806 29085 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[18]/VNB
flabel locali 32527 -4636 32561 -4602 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
flabel locali 31076 -4568 31110 -4534 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/CLK
rlabel viali 32527 -4636 32561 -4602 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel locali 32527 -4662 32575 -4582 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel locali 32467 -4582 32575 -4508 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 32515 -4642 32573 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 32455 -4596 32513 -4533 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 32455 -4605 32573 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 31795 -4605 31925 -4596 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 31795 -4633 32573 -4605 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
rlabel metal1 31795 -4642 31925 -4633 1 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/RESET_B
flabel locali 32800 -4571 32829 -4536 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/Q
flabel locali 33102 -4568 33124 -4535 0 FreeSans 200 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/Q_N
flabel locali 31076 -4500 31110 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/CLK
flabel locali 31351 -4500 31385 -4466 0 FreeSans 400 0 0 0 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/D
rlabel viali 31075 -4262 31109 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/VPWR
rlabel viali 31167 -4262 31201 -4228 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/VPB
rlabel viali 31075 -4806 31109 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/VGND
rlabel viali 31167 -4806 31201 -4772 3 20bitCounter_flat_0/sky130_fd_sc_hd__dfrbp_1_0[19]/VNB
flabel locali 12954 -1301 12983 -1266 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/Q
flabel locali 13256 -1298 13278 -1265 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/Q_N
flabel locali 12681 -1366 12715 -1332 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 11505 -1230 11539 -1196 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/D
flabel locali 11230 -1230 11264 -1196 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 11230 -1298 11264 -1264 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/CLK
flabel locali 12681 -1298 12715 -1264 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel metal1 11229 -1536 11263 -1502 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/VGND
flabel metal1 11229 -992 11263 -958 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/VPWR
flabel nwell 11229 -992 11263 -958 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/VPB
flabel pwell 11229 -1536 11263 -1502 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/VNB
rlabel comment 11200 -1519 11200 -1519 4 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/dfrbp_1
rlabel viali 12681 -1366 12715 -1332 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel viali 12621 -1303 12655 -1269 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 12681 -1392 12729 -1312 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel locali 12621 -1312 12729 -1238 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 12669 -1372 12727 -1363 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 12609 -1326 12667 -1263 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 12609 -1335 12727 -1326 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 11949 -1335 12079 -1326 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 11949 -1363 12727 -1335 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
rlabel metal1 11949 -1372 12079 -1363 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_1/RESET_B
flabel locali 10488 -1301 10517 -1266 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/Q
flabel locali 10790 -1298 10812 -1265 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/Q_N
flabel locali 10215 -1366 10249 -1332 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 9039 -1230 9073 -1196 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/D
flabel locali 8764 -1230 8798 -1196 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 8764 -1298 8798 -1264 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/CLK
flabel locali 10215 -1298 10249 -1264 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel metal1 8763 -1536 8797 -1502 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/VGND
flabel metal1 8763 -992 8797 -958 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/VPWR
flabel nwell 8763 -992 8797 -958 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/VPB
flabel pwell 8763 -1536 8797 -1502 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/VNB
rlabel comment 8734 -1519 8734 -1519 4 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/dfrbp_1
rlabel viali 10215 -1366 10249 -1332 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel viali 10155 -1303 10189 -1269 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 10215 -1392 10263 -1312 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel locali 10155 -1312 10263 -1238 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 10203 -1372 10261 -1363 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 10143 -1326 10201 -1263 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 10143 -1335 10261 -1326 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 9483 -1335 9613 -1326 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 9483 -1363 10261 -1335 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
rlabel metal1 9483 -1372 9613 -1363 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_0/RESET_B
flabel locali 12954 -2103 12983 -2068 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/Q
flabel locali 13256 -2100 13278 -2067 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/Q_N
flabel locali 12681 -2168 12715 -2134 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
flabel locali 11505 -2032 11539 -1998 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/D
flabel locali 11230 -2032 11264 -1998 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/CLK
flabel locali 11230 -2100 11264 -2066 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/CLK
flabel locali 12681 -2100 12715 -2066 0 FreeSans 400 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
flabel metal1 11229 -2338 11263 -2304 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/VGND
flabel metal1 11229 -1794 11263 -1760 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/VPWR
flabel nwell 11229 -1794 11263 -1760 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/VPB
flabel pwell 11229 -2338 11263 -2304 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/VNB
rlabel comment 11200 -2321 11200 -2321 4 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/dfrbp_1
rlabel viali 12681 -2168 12715 -2134 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel viali 12621 -2105 12655 -2071 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel locali 12681 -2194 12729 -2114 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel locali 12621 -2114 12729 -2040 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 12669 -2174 12727 -2165 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 12609 -2128 12667 -2065 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 12609 -2137 12727 -2128 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 11949 -2137 12079 -2128 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 11949 -2165 12727 -2137 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
rlabel metal1 11949 -2174 12079 -2165 1 static_freqDiv_0/sky130_fd_sc_hd__dfrbp_1_2/RESET_B
flabel locali 10181 -2100 10215 -2066 0 FreeSans 340 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/A
flabel locali 10273 -2168 10307 -2134 0 FreeSans 340 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/Y
flabel locali 10273 -2032 10307 -1998 0 FreeSans 340 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/Y
flabel locali 10273 -2100 10307 -2066 0 FreeSans 340 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/Y
flabel nwell 10181 -1794 10215 -1760 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/VPB
flabel pwell 10181 -2338 10215 -2304 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/VNB
flabel metal1 10181 -1794 10215 -1760 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/VPWR
flabel metal1 10181 -2338 10215 -2304 0 FreeSans 200 0 0 0 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/VGND
rlabel comment 10152 -2321 10152 -2321 4 static_freqDiv_0/sky130_fd_sc_hd__inv_2_0/inv_2
flabel locali -60736 4140 -60736 4140 0 FreeSans 320 0 0 0 extract1_0/net2
flabel locali -62234 4164 -62234 4164 0 FreeSans 320 0 0 0 extract1_0/net1
flabel metal1 -61750 3344 -61750 3344 0 FreeSans 320 0 0 0 extract1_0/in
flabel metal1 -61542 3358 -61542 3358 0 FreeSans 320 0 0 0 extract1_0/out
flabel locali -61318 3298 -61318 3298 0 FreeSans 480 0 0 0 extract1_0/clkb_in
flabel locali -61880 3000 -61880 3000 0 FreeSans 480 0 0 0 extract1_0/cl_in
flabel metal1 -15484 42578 -15484 42578 0 FreeSans 1600 0 0 0 wb_flat_0/vbias1
flabel metal1 -15820 42508 -15820 42508 0 FreeSans 1600 0 0 0 wb_flat_0/vbias2
flabel psubdiff -15328 14500 -15328 14500 0 FreeSans 1600 0 0 0 wb_flat_0/gnd
flabel metal3 31426 27128 31426 27128 0 FreeSans 1600 0 0 0 wb_flat_0/Bot_2
flabel metal4 34358 26184 34358 26184 0 FreeSans 1600 0 0 0 wb_flat_0/Top_2
flabel metal3 -13786 34218 -13786 34218 0 FreeSans 1600 0 0 0 wb_flat_0/Bot_1
flabel metal4 -11238 34274 -11238 34274 0 FreeSans 1600 0 0 0 wb_flat_0/Top_1
flabel metal1 -14810 30044 -14810 30044 0 FreeSans 1600 0 0 0 wb_flat_0/vinp2
flabel metal1 -16564 30024 -16564 30024 0 FreeSans 1600 0 0 0 wb_flat_0/vinp1
flabel metal4 6784 1400 6784 1400 0 FreeSans 1600 0 0 0 buff_final_flat_0/GND
flabel metal5 2090 5904 2090 5904 0 FreeSans 1600 0 0 0 buff_final_flat_0/VDD
flabel metal1 7550 4964 7550 4964 0 FreeSans 800 0 0 0 buff_final_flat_0/vinp1
flabel metal1 7466 4316 7466 4316 0 FreeSans 800 0 0 0 buff_final_flat_0/vinpch2
flabel metal2 7112 5578 7112 5580 0 FreeSans 800 0 0 0 buff_final_flat_0/outp1
flabel metal2 7098 5378 7098 5380 0 FreeSans 800 0 0 0 buff_final_flat_0/outp2
flabel locali 10324 3934 10324 3934 0 FreeSans 800 0 0 0 buff_final_flat_0/Bout
flabel locali 9148 3972 9148 3972 0 FreeSans 800 0 0 0 buff_final_flat_0/Bout_mirror
flabel metal3 11548 2598 11548 2598 0 FreeSans 800 0 0 0 buff_final_flat_0/outn1
flabel metal3 11508 3736 11508 3736 0 FreeSans 800 0 0 0 buff_final_flat_0/outn2
flabel locali 11204 3108 11204 3108 0 FreeSans 800 0 0 0 buff_final_flat_0/vinn1
flabel locali 11352 3204 11352 3204 0 FreeSans 800 0 0 0 buff_final_flat_0/vinnch1
flabel locali 11588 2146 11588 2146 0 FreeSans 800 0 0 0 buff_final_flat_0/vinnch2
flabel metal1 11630 2490 11630 2490 0 FreeSans 800 0 0 0 buff_final_flat_0/vinn2
flabel locali 3968 3412 3968 3412 0 FreeSans 800 0 0 0 buff_final_flat_0/outpch1
flabel locali 4944 3392 4944 3392 0 FreeSans 800 0 0 0 buff_final_flat_0/outpch2
flabel metal1 14492 6140 14492 6140 0 FreeSans 800 0 0 0 buff_final_flat_0/vbiasob
flabel metal1 5600 2896 5600 2896 0 FreeSans 800 0 0 0 buff_final_flat_0/vbiasot
flabel locali 11442 5200 11442 5200 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH_bar
flabel locali 6220 5198 6220 5198 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH_bar
flabel locali 952 5182 952 5182 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH_bar
flabel locali 1030 4460 1030 4460 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH
flabel locali 6186 4472 6186 4472 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH
flabel locali 11448 4488 11448 4488 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH
flabel locali 14658 3994 14658 3994 0 FreeSans 400 0 0 0 buff_final_flat_0/outnch1
flabel locali 15264 4002 15264 4002 0 FreeSans 400 0 0 0 buff_final_flat_0/outnch2
flabel metal1 7524 3964 7524 3964 0 FreeSans 400 0 0 0 buff_final_flat_0/vinp2
flabel metal2 7460 4762 7460 4762 0 FreeSans 400 0 0 0 buff_final_flat_0/vinpch1
flabel metal1 10754 5690 10754 5690 0 FreeSans 400 0 0 0 buff_final_flat_0/vbiaschopper
flabel locali 17082 5004 17082 5004 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH
flabel locali 17052 4272 17052 4272 0 FreeSans 400 0 0 0 buff_final_flat_0/Fvco_By4_QPH_bar
flabel via3 32624 1940 32624 1940 0 FreeSans 1600 0 0 0 edge_0/GND!
flabel viali 26732 2242 26732 2242 0 FreeSans 400 0 0 0 edge_0/n1
flabel locali 26994 2126 26994 2126 0 FreeSans 400 0 0 0 edge_0/net9
flabel locali 27606 2132 27606 2132 0 FreeSans 400 0 0 0 edge_0/net8
flabel locali 28190 2128 28190 2128 0 FreeSans 400 0 0 0 edge_0/net7
flabel locali 27286 2334 27286 2334 0 FreeSans 400 0 0 0 edge_0/n2
flabel locali 27864 2332 27864 2332 0 FreeSans 400 0 0 0 edge_0/n3
flabel locali 28442 2334 28442 2334 0 FreeSans 400 0 0 0 edge_0/n4
flabel locali 29040 2346 29040 2346 0 FreeSans 400 0 0 0 edge_0/n5
flabel locali 29618 2348 29618 2348 0 FreeSans 400 0 0 0 edge_0/n6
flabel locali 30186 2356 30186 2356 0 FreeSans 400 0 0 0 edge_0/n7
flabel locali 30770 2348 30770 2348 0 FreeSans 400 0 0 0 edge_0/n8
flabel locali 31354 2342 31354 2342 0 FreeSans 400 0 0 0 edge_0/n9
flabel locali 28766 2136 28766 2136 0 FreeSans 400 0 0 0 edge_0/net1
flabel locali 29340 2140 29340 2140 0 FreeSans 400 0 0 0 edge_0/net2
flabel locali 29916 2138 29916 2138 0 FreeSans 400 0 0 0 edge_0/net3
flabel locali 30498 2134 30498 2134 0 FreeSans 400 0 0 0 edge_0/net4
flabel locali 31084 2128 31084 2128 0 FreeSans 400 0 0 0 edge_0/net5
flabel locali 31644 2134 31644 2134 0 FreeSans 400 0 0 0 edge_0/net6
flabel metal1 27196 2152 27196 2152 0 FreeSans 400 0 0 0 edge_0/v1!
flabel metal1 27810 2158 27810 2158 0 FreeSans 400 0 0 0 edge_0/v2!
flabel metal1 28394 2154 28394 2154 0 FreeSans 400 0 0 0 edge_0/v3!
flabel metal1 28960 2160 28960 2160 0 FreeSans 400 0 0 0 edge_0/v4!
flabel metal1 30700 2158 30700 2158 0 FreeSans 400 0 0 0 edge_0/v7!
flabel metal1 31272 2166 31272 2166 0 FreeSans 400 0 0 0 edge_0/v8!
flabel metal1 31844 2170 31844 2170 0 FreeSans 400 0 0 0 edge_0/v9!
flabel metal1 30112 2164 30112 2164 0 FreeSans 400 0 0 0 edge_0/v6!
flabel metal1 29546 2160 29546 2160 0 FreeSans 400 0 0 0 edge_0/v5!
flabel locali 25918 3390 25918 3390 0 FreeSans 1600 0 0 0 edge_0/VDD
flabel metal1 28870 262 28870 262 0 FreeSans 400 0 0 0 edge_0/vout
flabel locali 28230 -198 28230 -198 0 FreeSans 400 0 0 0 edge_0/v1!
flabel locali 28742 -204 28742 -204 0 FreeSans 400 0 0 0 edge_0/v3!
flabel locali 28544 -122 28544 -122 0 FreeSans 400 0 0 0 edge_0/v4!
flabel locali 28352 306 28352 306 0 FreeSans 400 0 0 0 edge_0/v5!
flabel locali 28738 310 28738 310 0 FreeSans 400 0 0 0 edge_0/v6!
flabel locali 28546 382 28546 382 0 FreeSans 400 0 0 0 edge_0/v7!
flabel locali 29776 -328 29776 -328 0 FreeSans 400 0 0 0 edge_0/v1!
flabel locali 29676 426 29676 426 0 FreeSans 400 0 0 0 edge_0/v2!
flabel locali 29490 428 29490 428 0 FreeSans 400 0 0 0 edge_0/v4!
flabel locali 29290 422 29290 422 0 FreeSans 400 0 0 0 edge_0/v6!
flabel locali 29104 426 29104 426 0 FreeSans 400 0 0 0 edge_0/v8!
flabel locali 29586 -338 29586 -338 0 FreeSans 400 0 0 0 edge_0/v3!
flabel locali 29200 -336 29200 -336 0 FreeSans 400 0 0 0 edge_0/v7!
flabel locali 29004 -338 29004 -338 0 FreeSans 400 0 0 0 edge_0/v9!
flabel locali 29388 -334 29388 -334 0 FreeSans 400 0 0 0 edge_0/v5!
flabel locali 29054 128 29054 128 0 FreeSans 400 0 0 0 edge_0/net17!
flabel locali 29150 60 29150 60 0 FreeSans 400 0 0 0 edge_0/net16!
flabel locali 29244 120 29244 120 0 FreeSans 400 0 0 0 edge_0/net15!
flabel locali 29326 42 29326 42 0 FreeSans 400 0 0 0 edge_0/net14!
flabel locali 29418 106 29418 106 0 FreeSans 400 0 0 0 edge_0/net13!
flabel locali 29524 30 29524 30 0 FreeSans 400 0 0 0 edge_0/net12!
flabel locali 29614 98 29614 98 0 FreeSans 400 0 0 0 edge_0/net11!
flabel locali 29716 46 29716 46 0 FreeSans 400 0 0 0 edge_0/net10!
flabel locali 28718 800 28718 800 0 FreeSans 400 0 0 0 edge_0/v9!
flabel locali 28312 810 28312 810 0 FreeSans 400 0 0 0 edge_0/v8!
flabel locali 28554 -644 28554 -644 0 FreeSans 400 0 0 0 edge_0/v2!
<< end >>
