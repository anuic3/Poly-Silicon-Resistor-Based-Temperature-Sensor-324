magic
tech sky130A
magscale 1 2
timestamp 1634293258
<< viali >>
rect 2076 240 2114 274
rect 4192 240 4230 274
rect 6308 240 6346 274
rect 8424 240 8462 274
rect 10540 240 10578 274
rect 12656 240 12694 274
rect 14772 240 14810 274
rect 16888 240 16926 274
rect 19004 240 19042 274
rect 21120 240 21158 274
rect 23236 240 23274 274
rect 25352 240 25390 274
rect 27468 240 27506 274
rect 29584 240 29622 274
rect 31700 240 31738 274
rect 33816 240 33854 274
rect 35932 240 35970 274
rect 38048 240 38086 274
rect 40164 240 40202 274
rect 42280 240 42318 274
<< metal1 >>
rect 1409 294 1529 300
rect 1409 242 1433 294
rect 1485 242 1529 294
rect 1409 184 1529 242
rect 2045 282 2138 309
rect 2045 230 2069 282
rect 2121 230 2138 282
rect 2045 208 2138 230
rect 3525 294 3645 300
rect 3525 242 3549 294
rect 3601 242 3645 294
rect 3525 184 3645 242
rect 4161 282 4254 309
rect 4161 230 4185 282
rect 4237 230 4254 282
rect 4161 208 4254 230
rect 5641 294 5761 300
rect 5641 242 5665 294
rect 5717 242 5761 294
rect 5641 184 5761 242
rect 6277 282 6370 309
rect 6277 230 6301 282
rect 6353 230 6370 282
rect 6277 208 6370 230
rect 7757 294 7877 300
rect 7757 242 7781 294
rect 7833 242 7877 294
rect 7757 184 7877 242
rect 8393 282 8486 309
rect 8393 230 8417 282
rect 8469 230 8486 282
rect 8393 208 8486 230
rect 9873 294 9993 300
rect 9873 242 9897 294
rect 9949 242 9993 294
rect 9873 184 9993 242
rect 10509 282 10602 309
rect 10509 230 10533 282
rect 10585 230 10602 282
rect 10509 208 10602 230
rect 11989 294 12109 300
rect 11989 242 12013 294
rect 12065 242 12109 294
rect 11989 184 12109 242
rect 12625 282 12718 309
rect 12625 230 12649 282
rect 12701 230 12718 282
rect 12625 208 12718 230
rect 14105 294 14225 300
rect 14105 242 14129 294
rect 14181 242 14225 294
rect 14105 184 14225 242
rect 14741 282 14834 309
rect 14741 230 14765 282
rect 14817 230 14834 282
rect 14741 208 14834 230
rect 16221 294 16341 300
rect 16221 242 16245 294
rect 16297 242 16341 294
rect 16221 184 16341 242
rect 16857 282 16950 309
rect 16857 230 16881 282
rect 16933 230 16950 282
rect 16857 208 16950 230
rect 18337 294 18457 300
rect 18337 242 18361 294
rect 18413 242 18457 294
rect 18337 184 18457 242
rect 18973 282 19066 309
rect 18973 230 18997 282
rect 19049 230 19066 282
rect 18973 208 19066 230
rect 20453 294 20573 300
rect 20453 242 20477 294
rect 20529 242 20573 294
rect 20453 184 20573 242
rect 21089 282 21182 309
rect 21089 230 21113 282
rect 21165 230 21182 282
rect 21089 208 21182 230
rect 22569 294 22689 300
rect 22569 242 22593 294
rect 22645 242 22689 294
rect 22569 184 22689 242
rect 23205 282 23298 309
rect 23205 230 23229 282
rect 23281 230 23298 282
rect 23205 208 23298 230
rect 24685 294 24805 300
rect 24685 242 24709 294
rect 24761 242 24805 294
rect 24685 184 24805 242
rect 25321 282 25414 309
rect 25321 230 25345 282
rect 25397 230 25414 282
rect 25321 208 25414 230
rect 26801 294 26921 300
rect 26801 242 26825 294
rect 26877 242 26921 294
rect 26801 184 26921 242
rect 27437 282 27530 309
rect 27437 230 27461 282
rect 27513 230 27530 282
rect 27437 208 27530 230
rect 28917 294 29037 300
rect 28917 242 28941 294
rect 28993 242 29037 294
rect 28917 184 29037 242
rect 29553 282 29646 309
rect 29553 230 29577 282
rect 29629 230 29646 282
rect 29553 208 29646 230
rect 31033 294 31153 300
rect 31033 242 31057 294
rect 31109 242 31153 294
rect 31033 184 31153 242
rect 31669 282 31762 309
rect 31669 230 31693 282
rect 31745 230 31762 282
rect 31669 208 31762 230
rect 33149 294 33269 300
rect 33149 242 33173 294
rect 33225 242 33269 294
rect 33149 184 33269 242
rect 33785 282 33878 309
rect 33785 230 33809 282
rect 33861 230 33878 282
rect 33785 208 33878 230
rect 35265 294 35385 300
rect 35265 242 35289 294
rect 35341 242 35385 294
rect 35265 184 35385 242
rect 35901 282 35994 309
rect 35901 230 35925 282
rect 35977 230 35994 282
rect 35901 208 35994 230
rect 37381 294 37501 300
rect 37381 242 37405 294
rect 37457 242 37501 294
rect 37381 184 37501 242
rect 38017 282 38110 309
rect 38017 230 38041 282
rect 38093 230 38110 282
rect 38017 208 38110 230
rect 39497 294 39617 300
rect 39497 242 39521 294
rect 39573 242 39617 294
rect 39497 184 39617 242
rect 40133 282 40226 309
rect 40133 230 40157 282
rect 40209 230 40226 282
rect 40133 208 40226 230
rect 41613 294 41733 300
rect 41613 242 41637 294
rect 41689 242 41733 294
rect 41613 184 41733 242
rect 42249 282 42342 309
rect 42249 230 42273 282
rect 42325 230 42342 282
rect 42249 208 42342 230
<< via1 >>
rect 1433 242 1485 294
rect 2069 274 2121 282
rect 2069 240 2076 274
rect 2076 240 2114 274
rect 2114 240 2121 274
rect 2069 230 2121 240
rect 3549 242 3601 294
rect 4185 274 4237 282
rect 4185 240 4192 274
rect 4192 240 4230 274
rect 4230 240 4237 274
rect 4185 230 4237 240
rect 5665 242 5717 294
rect 6301 274 6353 282
rect 6301 240 6308 274
rect 6308 240 6346 274
rect 6346 240 6353 274
rect 6301 230 6353 240
rect 7781 242 7833 294
rect 8417 274 8469 282
rect 8417 240 8424 274
rect 8424 240 8462 274
rect 8462 240 8469 274
rect 8417 230 8469 240
rect 9897 242 9949 294
rect 10533 274 10585 282
rect 10533 240 10540 274
rect 10540 240 10578 274
rect 10578 240 10585 274
rect 10533 230 10585 240
rect 12013 242 12065 294
rect 12649 274 12701 282
rect 12649 240 12656 274
rect 12656 240 12694 274
rect 12694 240 12701 274
rect 12649 230 12701 240
rect 14129 242 14181 294
rect 14765 274 14817 282
rect 14765 240 14772 274
rect 14772 240 14810 274
rect 14810 240 14817 274
rect 14765 230 14817 240
rect 16245 242 16297 294
rect 16881 274 16933 282
rect 16881 240 16888 274
rect 16888 240 16926 274
rect 16926 240 16933 274
rect 16881 230 16933 240
rect 18361 242 18413 294
rect 18997 274 19049 282
rect 18997 240 19004 274
rect 19004 240 19042 274
rect 19042 240 19049 274
rect 18997 230 19049 240
rect 20477 242 20529 294
rect 21113 274 21165 282
rect 21113 240 21120 274
rect 21120 240 21158 274
rect 21158 240 21165 274
rect 21113 230 21165 240
rect 22593 242 22645 294
rect 23229 274 23281 282
rect 23229 240 23236 274
rect 23236 240 23274 274
rect 23274 240 23281 274
rect 23229 230 23281 240
rect 24709 242 24761 294
rect 25345 274 25397 282
rect 25345 240 25352 274
rect 25352 240 25390 274
rect 25390 240 25397 274
rect 25345 230 25397 240
rect 26825 242 26877 294
rect 27461 274 27513 282
rect 27461 240 27468 274
rect 27468 240 27506 274
rect 27506 240 27513 274
rect 27461 230 27513 240
rect 28941 242 28993 294
rect 29577 274 29629 282
rect 29577 240 29584 274
rect 29584 240 29622 274
rect 29622 240 29629 274
rect 29577 230 29629 240
rect 31057 242 31109 294
rect 31693 274 31745 282
rect 31693 240 31700 274
rect 31700 240 31738 274
rect 31738 240 31745 274
rect 31693 230 31745 240
rect 33173 242 33225 294
rect 33809 274 33861 282
rect 33809 240 33816 274
rect 33816 240 33854 274
rect 33854 240 33861 274
rect 33809 230 33861 240
rect 35289 242 35341 294
rect 35925 274 35977 282
rect 35925 240 35932 274
rect 35932 240 35970 274
rect 35970 240 35977 274
rect 35925 230 35977 240
rect 37405 242 37457 294
rect 38041 274 38093 282
rect 38041 240 38048 274
rect 38048 240 38086 274
rect 38086 240 38093 274
rect 38041 230 38093 240
rect 39521 242 39573 294
rect 40157 274 40209 282
rect 40157 240 40164 274
rect 40164 240 40202 274
rect 40202 240 40209 274
rect 40157 230 40209 240
rect 41637 242 41689 294
rect 42273 274 42325 282
rect 42273 240 42280 274
rect 42280 240 42318 274
rect 42318 240 42325 274
rect 42273 230 42325 240
rect 300 131 352 183
rect 2416 131 2468 183
rect 4532 131 4584 183
rect 6648 131 6700 183
rect 8764 131 8816 183
rect 10880 131 10932 183
rect 12996 131 13048 183
rect 15112 131 15164 183
rect 17228 131 17280 183
rect 19344 131 19396 183
rect 21460 131 21512 183
rect 23576 131 23628 183
rect 25692 131 25744 183
rect 27808 131 27860 183
rect 29924 131 29976 183
rect 32040 131 32092 183
rect 34156 131 34208 183
rect 36272 131 36324 183
rect 38388 131 38440 183
rect 40504 131 40556 183
<< metal2 >>
rect 1409 357 41733 426
rect 1409 294 1529 357
rect 1409 242 1433 294
rect 1485 242 1529 294
rect 1409 220 1529 242
rect 2045 282 2138 325
rect 2045 230 2069 282
rect 2121 230 2138 282
rect 2045 191 2138 230
rect 3525 294 3645 357
rect 3525 242 3549 294
rect 3601 242 3645 294
rect 3525 220 3645 242
rect 4161 282 4254 325
rect 4161 230 4185 282
rect 4237 230 4254 282
rect 4161 191 4254 230
rect 5641 294 5761 357
rect 5641 242 5665 294
rect 5717 242 5761 294
rect 5641 220 5761 242
rect 6277 282 6370 325
rect 6277 230 6301 282
rect 6353 230 6370 282
rect 6277 191 6370 230
rect 7757 294 7877 357
rect 7757 242 7781 294
rect 7833 242 7877 294
rect 7757 220 7877 242
rect 8393 282 8486 325
rect 8393 230 8417 282
rect 8469 230 8486 282
rect 8393 191 8486 230
rect 9873 294 9993 357
rect 9873 242 9897 294
rect 9949 242 9993 294
rect 9873 220 9993 242
rect 10509 282 10602 325
rect 10509 230 10533 282
rect 10585 230 10602 282
rect 10509 191 10602 230
rect 11989 294 12109 357
rect 11989 242 12013 294
rect 12065 242 12109 294
rect 11989 220 12109 242
rect 12625 282 12718 325
rect 12625 230 12649 282
rect 12701 230 12718 282
rect 12625 191 12718 230
rect 14105 294 14225 357
rect 14105 242 14129 294
rect 14181 242 14225 294
rect 14105 220 14225 242
rect 14741 282 14834 325
rect 14741 230 14765 282
rect 14817 230 14834 282
rect 14741 191 14834 230
rect 16221 294 16341 357
rect 16221 242 16245 294
rect 16297 242 16341 294
rect 16221 220 16341 242
rect 16857 282 16950 325
rect 16857 230 16881 282
rect 16933 230 16950 282
rect 16857 191 16950 230
rect 18337 294 18457 357
rect 18337 242 18361 294
rect 18413 242 18457 294
rect 18337 220 18457 242
rect 18973 282 19066 325
rect 18973 230 18997 282
rect 19049 230 19066 282
rect 18973 191 19066 230
rect 20453 294 20573 357
rect 20453 242 20477 294
rect 20529 242 20573 294
rect 20453 220 20573 242
rect 21089 282 21182 325
rect 21089 230 21113 282
rect 21165 230 21182 282
rect 21089 191 21182 230
rect 22569 294 22689 357
rect 22569 242 22593 294
rect 22645 242 22689 294
rect 22569 220 22689 242
rect 23205 282 23298 325
rect 23205 230 23229 282
rect 23281 230 23298 282
rect 23205 191 23298 230
rect 24685 294 24805 357
rect 24685 242 24709 294
rect 24761 242 24805 294
rect 24685 220 24805 242
rect 25321 282 25414 325
rect 25321 230 25345 282
rect 25397 230 25414 282
rect 25321 191 25414 230
rect 26801 294 26921 357
rect 26801 242 26825 294
rect 26877 242 26921 294
rect 26801 220 26921 242
rect 27437 282 27530 325
rect 27437 230 27461 282
rect 27513 230 27530 282
rect 27437 191 27530 230
rect 28917 294 29037 357
rect 28917 242 28941 294
rect 28993 242 29037 294
rect 28917 220 29037 242
rect 29553 282 29646 325
rect 29553 230 29577 282
rect 29629 230 29646 282
rect 29553 191 29646 230
rect 31033 294 31153 357
rect 31033 242 31057 294
rect 31109 242 31153 294
rect 31033 220 31153 242
rect 31669 282 31762 325
rect 31669 230 31693 282
rect 31745 230 31762 282
rect 31669 191 31762 230
rect 33149 294 33269 357
rect 33149 242 33173 294
rect 33225 242 33269 294
rect 33149 220 33269 242
rect 33785 282 33878 325
rect 33785 230 33809 282
rect 33861 230 33878 282
rect 33785 191 33878 230
rect 35265 294 35385 357
rect 35265 242 35289 294
rect 35341 242 35385 294
rect 35265 220 35385 242
rect 35901 282 35994 325
rect 35901 230 35925 282
rect 35977 230 35994 282
rect 35901 191 35994 230
rect 37381 294 37501 357
rect 37381 242 37405 294
rect 37457 242 37501 294
rect 37381 220 37501 242
rect 38017 282 38110 325
rect 38017 230 38041 282
rect 38093 230 38110 282
rect 38017 191 38110 230
rect 39497 294 39617 357
rect 39497 242 39521 294
rect 39573 242 39617 294
rect 39497 220 39617 242
rect 40133 282 40226 325
rect 40133 230 40157 282
rect 40209 230 40226 282
rect 40133 191 40226 230
rect 41613 294 41733 357
rect 41613 242 41637 294
rect 41689 242 41733 294
rect 41613 220 41733 242
rect 42249 282 42342 325
rect 42249 230 42273 282
rect 42325 230 42342 282
rect 42249 191 42342 230
rect 249 183 2138 191
rect 249 131 300 183
rect 352 131 2138 183
rect 249 122 2138 131
rect 2365 183 4254 191
rect 2365 131 2416 183
rect 2468 131 4254 183
rect 2365 122 4254 131
rect 4481 183 6370 191
rect 4481 131 4532 183
rect 4584 131 6370 183
rect 4481 122 6370 131
rect 6597 183 8486 191
rect 6597 131 6648 183
rect 6700 131 8486 183
rect 6597 122 8486 131
rect 8713 183 10602 191
rect 8713 131 8764 183
rect 8816 131 10602 183
rect 8713 122 10602 131
rect 10829 183 12718 191
rect 10829 131 10880 183
rect 10932 131 12718 183
rect 10829 122 12718 131
rect 12945 183 14834 191
rect 12945 131 12996 183
rect 13048 131 14834 183
rect 12945 122 14834 131
rect 15061 183 16950 191
rect 15061 131 15112 183
rect 15164 131 16950 183
rect 15061 122 16950 131
rect 17177 183 19066 191
rect 17177 131 17228 183
rect 17280 131 19066 183
rect 17177 122 19066 131
rect 19293 183 21182 191
rect 19293 131 19344 183
rect 19396 131 21182 183
rect 19293 122 21182 131
rect 21409 183 23298 191
rect 21409 131 21460 183
rect 21512 131 23298 183
rect 21409 122 23298 131
rect 23525 183 25414 191
rect 23525 131 23576 183
rect 23628 131 25414 183
rect 23525 122 25414 131
rect 25641 183 27530 191
rect 25641 131 25692 183
rect 25744 131 27530 183
rect 25641 122 27530 131
rect 27757 183 29646 191
rect 27757 131 27808 183
rect 27860 131 29646 183
rect 27757 122 29646 131
rect 29873 183 31762 191
rect 29873 131 29924 183
rect 29976 131 31762 183
rect 29873 122 31762 131
rect 31989 183 33878 191
rect 31989 131 32040 183
rect 32092 131 33878 183
rect 31989 122 33878 131
rect 34105 183 35994 191
rect 34105 131 34156 183
rect 34208 131 35994 183
rect 34105 122 35994 131
rect 36221 183 38110 191
rect 36221 131 36272 183
rect 36324 131 38110 183
rect 36221 122 38110 131
rect 38337 183 40226 191
rect 38337 131 38388 183
rect 38440 131 40226 183
rect 38337 122 40226 131
rect 40453 183 42342 191
rect 40453 131 40504 183
rect 40556 131 42342 183
rect 40453 122 42342 131
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
array 0 19 2116 0 0 640
timestamp 1634293258
transform 1 0 0 0 1 0
box -38 -77 2154 621
<< end >>
