magic
tech sky130A
magscale 1 2
timestamp 1634876261
<< psubdiff >>
rect -5852 39628 -4018 39714
rect -6540 39592 -4018 39628
rect -6540 39046 53570 39592
rect -6540 38318 -4336 39046
rect -2950 38318 -336 39046
rect 1050 38318 3664 39046
rect 5050 38318 7664 39046
rect 9050 38318 11664 39046
rect 13050 38318 15664 39046
rect 17050 38318 19664 39046
rect 21050 38318 23664 39046
rect 25050 38318 27664 39046
rect 29050 38318 31664 39046
rect 33050 38318 35664 39046
rect 37050 38318 39664 39046
rect 41050 38318 43664 39046
rect 45050 38318 47664 39046
rect 49050 38318 51664 39046
rect 53050 38318 53570 39046
rect -6540 37696 53570 38318
rect -6540 36882 -4018 37696
rect -6540 36154 -6072 36882
rect -4686 36154 -4018 36882
rect -6540 32882 -4018 36154
rect -6540 32154 -6072 32882
rect -4686 32154 -4018 32882
rect 51308 35844 53508 37696
rect 51308 35116 51706 35844
rect 53092 35116 53508 35844
rect -6540 28882 -4018 32154
rect -6540 28154 -6072 28882
rect -4686 28154 -4018 28882
rect -6540 24882 -4018 28154
rect 51308 31844 53508 35116
rect 51308 31116 51706 31844
rect 53092 31116 53508 31844
rect 51308 27844 53508 31116
rect 51308 27116 51706 27844
rect 53092 27116 53508 27844
rect -6540 24154 -6072 24882
rect -4686 24154 -4018 24882
rect -6540 20882 -4018 24154
rect -6540 20154 -6072 20882
rect -4686 20154 -4018 20882
rect -6540 16882 -4018 20154
rect 51308 23844 53508 27116
rect 51308 23116 51706 23844
rect 53092 23116 53508 23844
rect 51308 19844 53508 23116
rect 51308 19116 51706 19844
rect 53092 19116 53508 19844
rect -6540 16154 -6072 16882
rect -4686 16154 -4018 16882
rect -6540 12882 -4018 16154
rect 51308 15844 53508 19116
rect 51308 15116 51706 15844
rect 53092 15116 53508 15844
rect -6540 12154 -6072 12882
rect -4686 12154 -4018 12882
rect -6540 8882 -4018 12154
rect -6540 8154 -6072 8882
rect -4686 8154 -4018 8882
rect -6540 4882 -4018 8154
rect 51308 11844 53508 15116
rect 51308 11116 51706 11844
rect 53092 11116 53508 11844
rect 51308 7844 53508 11116
rect 51308 7116 51706 7844
rect 53092 7116 53508 7844
rect -6540 4154 -6072 4882
rect -4686 4154 -4018 4882
rect -6540 882 -4018 4154
rect -6540 154 -6072 882
rect -4686 154 -4018 882
rect -6540 -1734 -4018 154
rect 51308 3844 53508 7116
rect 51308 3116 51706 3844
rect 53092 3116 53508 3844
rect 51308 -156 53508 3116
rect 51308 -884 51706 -156
rect 53092 -884 53508 -156
rect 51308 -1734 53508 -884
rect -6540 -2236 53508 -1734
rect -6540 -2964 -3410 -2236
rect -2024 -2964 590 -2236
rect 1976 -2964 4590 -2236
rect 5976 -2964 8590 -2236
rect 9976 -2964 12590 -2236
rect 13976 -2964 16590 -2236
rect 17976 -2964 20590 -2236
rect 21976 -2964 24590 -2236
rect 25976 -2964 28590 -2236
rect 29976 -2964 32590 -2236
rect 33976 -2964 36590 -2236
rect 37976 -2964 40590 -2236
rect 41976 -2964 44590 -2236
rect 45976 -2964 48590 -2236
rect 49976 -2964 53508 -2236
rect -6540 -3386 53508 -2964
rect -6540 -3478 -4018 -3386
rect 51308 -3446 53508 -3386
rect -5852 -3568 -4018 -3478
<< psubdiffcont >>
rect -4336 38318 -2950 39046
rect -336 38318 1050 39046
rect 3664 38318 5050 39046
rect 7664 38318 9050 39046
rect 11664 38318 13050 39046
rect 15664 38318 17050 39046
rect 19664 38318 21050 39046
rect 23664 38318 25050 39046
rect 27664 38318 29050 39046
rect 31664 38318 33050 39046
rect 35664 38318 37050 39046
rect 39664 38318 41050 39046
rect 43664 38318 45050 39046
rect 47664 38318 49050 39046
rect 51664 38318 53050 39046
rect -6072 36154 -4686 36882
rect -6072 32154 -4686 32882
rect 51706 35116 53092 35844
rect -6072 28154 -4686 28882
rect 51706 31116 53092 31844
rect 51706 27116 53092 27844
rect -6072 24154 -4686 24882
rect -6072 20154 -4686 20882
rect 51706 23116 53092 23844
rect 51706 19116 53092 19844
rect -6072 16154 -4686 16882
rect 51706 15116 53092 15844
rect -6072 12154 -4686 12882
rect -6072 8154 -4686 8882
rect 51706 11116 53092 11844
rect 51706 7116 53092 7844
rect -6072 4154 -4686 4882
rect -6072 154 -4686 882
rect 51706 3116 53092 3844
rect 51706 -884 53092 -156
rect -3410 -2964 -2024 -2236
rect 590 -2964 1976 -2236
rect 4590 -2964 5976 -2236
rect 8590 -2964 9976 -2236
rect 12590 -2964 13976 -2236
rect 16590 -2964 17976 -2236
rect 20590 -2964 21976 -2236
rect 24590 -2964 25976 -2236
rect 28590 -2964 29976 -2236
rect 32590 -2964 33976 -2236
rect 36590 -2964 37976 -2236
rect 40590 -2964 41976 -2236
rect 44590 -2964 45976 -2236
rect 48590 -2964 49976 -2236
<< xpolycontact >>
rect -1614 32104 -1544 32536
rect -1614 26946 -1544 27378
rect -1296 32104 -1226 32536
rect -1296 26946 -1226 27378
rect -978 32104 -908 32536
rect -978 26946 -908 27378
rect -660 32104 -590 32536
rect -660 26946 -590 27378
rect -1562 24826 -1492 25258
rect -1562 19668 -1492 20100
rect -1206 24808 -1136 25240
rect -1206 19650 -1136 20082
rect -888 24808 -818 25240
rect -888 19650 -818 20082
rect -490 24790 -420 25222
rect -490 19632 -420 20064
rect -1570 18326 -1500 18758
rect -1570 13168 -1500 13600
rect -1232 18346 -1162 18778
rect -1232 13188 -1162 13620
rect -914 18346 -844 18778
rect -914 13188 -844 13620
rect -544 18344 -474 18776
rect -544 13186 -474 13618
rect -1548 11574 -1478 12006
rect -1548 6416 -1478 6848
rect -1230 11574 -1160 12006
rect -1230 6416 -1160 6848
rect -912 11574 -842 12006
rect -912 6416 -842 6848
rect -594 11574 -524 12006
rect -594 6416 -524 6848
<< xpolyres >>
rect -1614 27378 -1544 32104
rect -1296 27378 -1226 32104
rect -978 27378 -908 32104
rect -660 27378 -590 32104
rect -1562 20100 -1492 24826
rect -1206 20082 -1136 24808
rect -888 20082 -818 24808
rect -490 20064 -420 24790
rect -1570 13600 -1500 18326
rect -1232 13620 -1162 18346
rect -914 13620 -844 18346
rect -544 13618 -474 18344
rect -1548 6848 -1478 11574
rect -1230 6848 -1160 11574
rect -912 6848 -842 11574
rect -594 6848 -524 11574
<< locali >>
rect -4578 39046 -2740 39306
rect -4578 38318 -4336 39046
rect -2950 38318 -2740 39046
rect -4578 38076 -2740 38318
rect -578 39046 1260 39306
rect -578 38318 -336 39046
rect 1050 38318 1260 39046
rect -578 38076 1260 38318
rect 3422 39046 5260 39306
rect 3422 38318 3664 39046
rect 5050 38318 5260 39046
rect 3422 38076 5260 38318
rect 7422 39046 9260 39306
rect 7422 38318 7664 39046
rect 9050 38318 9260 39046
rect 7422 38076 9260 38318
rect 11422 39046 13260 39306
rect 11422 38318 11664 39046
rect 13050 38318 13260 39046
rect 11422 38076 13260 38318
rect 15422 39046 17260 39306
rect 15422 38318 15664 39046
rect 17050 38318 17260 39046
rect 15422 38076 17260 38318
rect 19422 39046 21260 39306
rect 19422 38318 19664 39046
rect 21050 38318 21260 39046
rect 19422 38076 21260 38318
rect 23422 39046 25260 39306
rect 23422 38318 23664 39046
rect 25050 38318 25260 39046
rect 23422 38076 25260 38318
rect 27422 39046 29260 39306
rect 27422 38318 27664 39046
rect 29050 38318 29260 39046
rect 27422 38076 29260 38318
rect 31422 39046 33260 39306
rect 31422 38318 31664 39046
rect 33050 38318 33260 39046
rect 31422 38076 33260 38318
rect 35422 39046 37260 39306
rect 35422 38318 35664 39046
rect 37050 38318 37260 39046
rect 35422 38076 37260 38318
rect 39422 39046 41260 39306
rect 39422 38318 39664 39046
rect 41050 38318 41260 39046
rect 39422 38076 41260 38318
rect 43422 39046 45260 39306
rect 43422 38318 43664 39046
rect 45050 38318 45260 39046
rect 43422 38076 45260 38318
rect 47422 39046 49260 39306
rect 47422 38318 47664 39046
rect 49050 38318 49260 39046
rect 47422 38076 49260 38318
rect 51422 39046 53260 39306
rect 51422 38318 51664 39046
rect 53050 38318 53260 39046
rect 51422 38076 53260 38318
rect -6314 36882 -4476 37142
rect -6314 36154 -6072 36882
rect -4686 36154 -4476 36882
rect -6314 35912 -4476 36154
rect 51464 35844 53302 36112
rect 51464 35116 51706 35844
rect 53092 35116 53302 35844
rect 51464 34874 53302 35116
rect -6314 32882 -4476 33142
rect -6314 32154 -6072 32882
rect -4686 32154 -4476 32882
rect -6314 31912 -4476 32154
rect 51464 31844 53302 32112
rect 51464 31116 51706 31844
rect 53092 31116 53302 31844
rect 51464 30874 53302 31116
rect -6314 28882 -4476 29142
rect -6314 28154 -6072 28882
rect -4686 28154 -4476 28882
rect -6314 27912 -4476 28154
rect 51464 27844 53302 28112
rect 51464 27116 51706 27844
rect 53092 27116 53302 27844
rect 51464 26874 53302 27116
rect -6314 24882 -4476 25142
rect -6314 24154 -6072 24882
rect -4686 24154 -4476 24882
rect -6314 23912 -4476 24154
rect 51464 23844 53302 24112
rect 51464 23116 51706 23844
rect 53092 23116 53302 23844
rect 51464 22874 53302 23116
rect -6314 20882 -4476 21142
rect -6314 20154 -6072 20882
rect -4686 20154 -4476 20882
rect -6314 19912 -4476 20154
rect 51464 19844 53302 20112
rect 51464 19116 51706 19844
rect 53092 19116 53302 19844
rect 51464 18874 53302 19116
rect -6314 16882 -4476 17142
rect -6314 16154 -6072 16882
rect -4686 16154 -4476 16882
rect -6314 15912 -4476 16154
rect 51464 15844 53302 16112
rect 51464 15116 51706 15844
rect 53092 15116 53302 15844
rect 51464 14874 53302 15116
rect -6314 12882 -4476 13142
rect -6314 12154 -6072 12882
rect -4686 12154 -4476 12882
rect -6314 11912 -4476 12154
rect 51464 11844 53302 12112
rect 51464 11116 51706 11844
rect 53092 11116 53302 11844
rect 51464 10874 53302 11116
rect -6314 8882 -4476 9142
rect -6314 8154 -6072 8882
rect -4686 8154 -4476 8882
rect -6314 7912 -4476 8154
rect 51464 7844 53302 8112
rect 51464 7116 51706 7844
rect 53092 7116 53302 7844
rect 51464 6874 53302 7116
rect -6314 4882 -4476 5142
rect -6314 4154 -6072 4882
rect -4686 4154 -4476 4882
rect -6314 3912 -4476 4154
rect 51464 3844 53302 4112
rect 51464 3116 51706 3844
rect 53092 3116 53302 3844
rect 51464 2874 53302 3116
rect -6314 882 -4476 1142
rect -6314 154 -6072 882
rect -4686 154 -4476 882
rect -6314 -88 -4476 154
rect 51464 -156 53302 112
rect 51464 -884 51706 -156
rect 53092 -884 53302 -156
rect 51464 -1126 53302 -884
rect -3652 -2236 -1814 -1960
rect -3652 -2964 -3410 -2236
rect -2024 -2964 -1814 -2236
rect -3652 -3206 -1814 -2964
rect 348 -2060 536 -1964
rect 1076 -2060 2186 -1964
rect 348 -2236 2186 -2060
rect 348 -2964 590 -2236
rect 1976 -2964 2186 -2236
rect 348 -3206 2186 -2964
rect 4348 -2236 6186 -1964
rect 4348 -2964 4590 -2236
rect 5976 -2964 6186 -2236
rect 4348 -3206 6186 -2964
rect 8348 -2236 10186 -1964
rect 8348 -2964 8590 -2236
rect 9976 -2964 10186 -2236
rect 8348 -3206 10186 -2964
rect 12348 -2236 14186 -1964
rect 12348 -2964 12590 -2236
rect 13976 -2964 14186 -2236
rect 12348 -3206 14186 -2964
rect 16348 -2236 18186 -1964
rect 16348 -2964 16590 -2236
rect 17976 -2964 18186 -2236
rect 16348 -3206 18186 -2964
rect 20348 -2236 22186 -1964
rect 20348 -2964 20590 -2236
rect 21976 -2964 22186 -2236
rect 20348 -3206 22186 -2964
rect 24348 -2236 26186 -1964
rect 24348 -2964 24590 -2236
rect 25976 -2964 26186 -2236
rect 24348 -3206 26186 -2964
rect 28348 -2236 30186 -1964
rect 28348 -2964 28590 -2236
rect 29976 -2964 30186 -2236
rect 28348 -3206 30186 -2964
rect 32348 -2236 34186 -1964
rect 32348 -2964 32590 -2236
rect 33976 -2964 34186 -2236
rect 32348 -3206 34186 -2964
rect 36348 -2236 38186 -1964
rect 36348 -2964 36590 -2236
rect 37976 -2964 38186 -2236
rect 36348 -3206 38186 -2964
rect 40348 -2236 42186 -1964
rect 40348 -2964 40590 -2236
rect 41976 -2964 42186 -2236
rect 40348 -3206 42186 -2964
rect 44348 -2236 46186 -1964
rect 44348 -2964 44590 -2236
rect 45976 -2964 46186 -2236
rect 44348 -3206 46186 -2964
rect 48348 -2236 50186 -1964
rect 48348 -2964 48590 -2236
rect 49976 -2964 50186 -2236
rect 48348 -3206 50186 -2964
<< viali >>
rect -4336 38318 -2950 39046
rect -336 38318 1050 39046
rect 3664 38318 5050 39046
rect 7664 38318 9050 39046
rect 11664 38318 13050 39046
rect 15664 38318 17050 39046
rect 19664 38318 21050 39046
rect 23664 38318 25050 39046
rect 27664 38318 29050 39046
rect 31664 38318 33050 39046
rect 35664 38318 37050 39046
rect 39664 38318 41050 39046
rect 43664 38318 45050 39046
rect 47664 38318 49050 39046
rect 51664 38318 53050 39046
rect -6072 36154 -4686 36882
rect 51706 35116 53092 35844
rect -6072 32154 -4686 32882
rect -1598 32121 -1560 32518
rect -1280 32121 -1242 32518
rect -962 32121 -924 32518
rect -644 32121 -606 32518
rect 51706 31116 53092 31844
rect -6072 28154 -4686 28882
rect -1598 26964 -1560 27361
rect -1280 26964 -1242 27361
rect -962 26964 -924 27361
rect -644 26964 -606 27361
rect 51706 27116 53092 27844
rect -888 25240 -816 25242
rect -6072 24154 -4686 24882
rect -1546 24843 -1508 25240
rect -1210 24808 -1206 25240
rect -1206 24808 -1138 25240
rect -888 24810 -818 25240
rect -818 24810 -816 25240
rect -474 24807 -436 25204
rect 51706 23116 53092 23844
rect -6072 20154 -4686 20882
rect -1546 19686 -1508 20083
rect -1208 19650 -1206 20082
rect -1206 19650 -1136 20082
rect -890 19650 -888 20078
rect -888 19650 -818 20078
rect -890 19646 -818 19650
rect -474 19650 -436 20047
rect 51706 19116 53092 19844
rect -1554 18343 -1516 18740
rect -1234 18346 -1232 18778
rect -1232 18346 -1162 18778
rect -914 18346 -844 18778
rect -844 18346 -842 18778
rect -528 18361 -490 18758
rect -6072 16154 -4686 16882
rect 51706 15116 53092 15844
rect -1554 13186 -1516 13583
rect -1234 13188 -1232 13620
rect -1232 13188 -1162 13620
rect -1162 13188 -1160 13620
rect -1234 13186 -1160 13188
rect -916 13188 -914 13620
rect -914 13188 -844 13620
rect -844 13188 -842 13620
rect -916 13186 -842 13188
rect -528 13204 -490 13601
rect -6072 12154 -4686 12882
rect -1532 11591 -1494 11988
rect -1214 11591 -1176 11988
rect -896 11591 -858 11988
rect -578 11591 -540 11988
rect 51706 11116 53092 11844
rect -6072 8154 -4686 8882
rect 51706 7116 53092 7844
rect -1532 6434 -1494 6831
rect -1214 6434 -1176 6831
rect -896 6434 -858 6831
rect -578 6434 -540 6831
rect -6072 4154 -4686 4882
rect 51706 3116 53092 3844
rect -6072 154 -4686 882
rect 51706 -884 53092 -156
rect -3410 -2964 -2024 -2236
rect 590 -2964 1976 -2236
rect 4590 -2964 5976 -2236
rect 8590 -2964 9976 -2236
rect 12590 -2964 13976 -2236
rect 16590 -2964 17976 -2236
rect 20590 -2964 21976 -2236
rect 24590 -2964 25976 -2236
rect 28590 -2964 29976 -2236
rect 32590 -2964 33976 -2236
rect 36590 -2964 37976 -2236
rect 40590 -2964 41976 -2236
rect 44590 -2964 45976 -2236
rect 48590 -2964 49976 -2236
<< metal1 >>
rect -4578 39046 -2740 39306
rect -4578 38318 -4336 39046
rect -2950 38318 -2740 39046
rect -4578 38076 -2740 38318
rect -578 39046 1260 39306
rect -578 38318 -336 39046
rect 1050 38318 1260 39046
rect -578 38076 1260 38318
rect 3422 39046 5260 39306
rect 3422 38318 3664 39046
rect 5050 38318 5260 39046
rect 3422 38076 5260 38318
rect 7422 39046 9260 39306
rect 7422 38318 7664 39046
rect 9050 38318 9260 39046
rect 7422 38076 9260 38318
rect 11422 39046 13260 39306
rect 11422 38318 11664 39046
rect 13050 38318 13260 39046
rect 11422 38076 13260 38318
rect 15422 39046 17260 39306
rect 15422 38318 15664 39046
rect 17050 38318 17260 39046
rect 15422 38076 17260 38318
rect 19422 39046 21260 39306
rect 19422 38318 19664 39046
rect 21050 38318 21260 39046
rect 19422 38076 21260 38318
rect 23422 39046 25260 39306
rect 23422 38318 23664 39046
rect 25050 38318 25260 39046
rect 23422 38076 25260 38318
rect 27422 39046 29260 39306
rect 27422 38318 27664 39046
rect 29050 38318 29260 39046
rect 27422 38076 29260 38318
rect 31422 39046 33260 39306
rect 31422 38318 31664 39046
rect 33050 38318 33260 39046
rect 31422 38076 33260 38318
rect 35422 39046 37260 39306
rect 35422 38318 35664 39046
rect 37050 38318 37260 39046
rect 35422 38076 37260 38318
rect 39422 39046 41260 39306
rect 39422 38318 39664 39046
rect 41050 38318 41260 39046
rect 39422 38076 41260 38318
rect 43422 39046 45260 39306
rect 43422 38318 43664 39046
rect 45050 38318 45260 39046
rect 43422 38076 45260 38318
rect 47422 39046 49260 39306
rect 47422 38318 47664 39046
rect 49050 38318 49260 39046
rect 47422 38076 49260 38318
rect 51422 39046 53260 39306
rect 51422 38318 51664 39046
rect 53050 38318 53260 39046
rect 51422 38076 53260 38318
rect -6314 36882 -4476 37142
rect -6314 36154 -6072 36882
rect -4686 36154 -4476 36882
rect -6314 35912 -4476 36154
rect 51464 35844 53302 36112
rect 51464 35116 51706 35844
rect 53092 35116 53302 35844
rect 51464 34874 53302 35116
rect -6314 32882 -4476 33142
rect -6314 32154 -6072 32882
rect -4686 32154 -4476 32882
rect -6314 31912 -4476 32154
rect -1634 32540 -566 32552
rect -1634 32104 -1618 32540
rect -1542 32104 -1298 32540
rect -1222 32104 -982 32540
rect -906 32104 -662 32540
rect -586 32104 -566 32540
rect -1634 32086 -566 32104
rect 51464 31844 53302 32112
rect 51464 31116 51706 31844
rect 53092 31116 53302 31844
rect 51464 30874 53302 31116
rect -6314 28882 -4476 29142
rect -6314 28154 -6072 28882
rect -4686 28154 -4476 28882
rect -6314 27912 -4476 28154
rect 51464 27844 53302 28112
rect -1636 27378 -568 27386
rect -1636 26946 -1614 27378
rect -1542 26946 -1298 27378
rect -1226 26946 -978 27378
rect -906 26946 -662 27378
rect -590 26946 -568 27378
rect -1636 26920 -568 26946
rect 51464 27116 51706 27844
rect 53092 27116 53302 27844
rect 51464 26874 53302 27116
rect -1578 25256 -1472 25272
rect -6314 24882 -4476 25142
rect -6314 24154 -6072 24882
rect -4686 24154 -4476 24882
rect -1578 24824 -1562 25256
rect -1490 24824 -1472 25256
rect -1230 25240 -1120 25556
rect -1230 25180 -1210 25240
rect -1578 24814 -1472 24824
rect -1226 24808 -1210 25180
rect -1138 24808 -1120 25240
rect -908 25242 -798 25576
rect -908 25200 -888 25242
rect -1226 24800 -1120 24808
rect -904 24810 -888 25200
rect -816 24810 -798 25242
rect -904 24800 -798 24810
rect -510 25228 -404 25238
rect -510 24796 -492 25228
rect -420 24796 -404 25228
rect -510 24780 -404 24796
rect -6314 23912 -4476 24154
rect 51464 23844 53302 24112
rect 51464 23116 51706 23844
rect 53092 23116 53302 23844
rect 51464 22874 53302 23116
rect -6314 20882 -4476 21142
rect -6314 20154 -6072 20882
rect -4686 20154 -4476 20882
rect -6314 19912 -4476 20154
rect -1578 20100 -1472 20112
rect -1578 19668 -1564 20100
rect -1490 19668 -1472 20100
rect -1220 20090 -1134 20094
rect -1220 20082 -1124 20090
rect -1220 20060 -1208 20082
rect -1578 19654 -1472 19668
rect -1218 19650 -1208 20060
rect -1136 19650 -1124 20082
rect -1218 19336 -1124 19650
rect -908 20078 -802 20094
rect -908 19646 -890 20078
rect -818 19646 -802 20078
rect -908 19408 -802 19646
rect -508 20060 -402 20074
rect -508 19628 -492 20060
rect -418 19628 -402 20060
rect -508 19616 -402 19628
rect 51464 19844 53302 20112
rect 3026 19480 3308 19568
rect 3026 19408 3064 19480
rect -908 19364 3064 19408
rect -908 19358 -248 19364
rect -908 19354 -802 19358
rect -1858 19328 -1124 19336
rect -2926 19276 -1124 19328
rect -218 19314 -176 19316
rect -218 19284 994 19314
rect -218 19282 264 19284
rect -2924 18916 -2844 19276
rect -1858 19274 -1136 19276
rect -6314 16882 -4476 17142
rect -2922 16938 -2844 18916
rect -2762 18858 -1852 18864
rect -1244 18858 -1152 18862
rect -2762 18814 -1152 18858
rect -2762 18796 -1650 18814
rect -1418 18796 -1152 18814
rect -2762 18794 -1852 18796
rect -2762 18778 -2126 18794
rect -1244 18778 -1152 18796
rect -6314 16154 -6072 16882
rect -4686 16154 -4476 16882
rect -6314 15912 -4476 16154
rect -2926 16812 -2844 16938
rect -2926 14294 -2852 16812
rect -2926 14254 -2848 14294
rect -6314 12882 -4476 13142
rect -6314 12154 -6072 12882
rect -4686 12154 -4476 12882
rect -6314 11912 -4476 12154
rect -2922 11714 -2848 14254
rect -2922 11610 -2842 11714
rect -2916 9142 -2842 11610
rect -6314 8882 -4476 9142
rect -6314 8154 -6072 8882
rect -4686 8154 -4476 8882
rect -6314 7912 -4476 8154
rect -2922 9030 -2842 9142
rect -2922 6458 -2848 9030
rect -2758 6594 -2652 18778
rect -1592 18764 -1480 18772
rect -1592 18332 -1572 18764
rect -1498 18332 -1480 18764
rect -1592 18312 -1480 18332
rect -1244 18346 -1234 18778
rect -1162 18346 -1152 18778
rect -1244 18330 -1152 18346
rect -926 18850 -830 18852
rect -218 18850 -176 19282
rect 716 19194 994 19284
rect 716 19018 766 19194
rect 954 19018 994 19194
rect 3026 19246 3064 19364
rect 3264 19246 3308 19480
rect 3026 19166 3308 19246
rect 716 18928 994 19018
rect 51464 19116 51706 19844
rect 53092 19116 53302 19844
rect 51464 18874 53302 19116
rect -926 18816 -140 18850
rect -926 18810 -604 18816
rect -422 18810 -140 18816
rect -926 18778 -830 18810
rect -926 18346 -914 18778
rect -842 18346 -830 18778
rect -926 18332 -830 18346
rect -572 18774 -450 18788
rect -572 18342 -548 18774
rect -474 18342 -450 18774
rect -572 18322 -450 18342
rect 25738 17086 26516 17138
rect 25738 16990 26014 17086
rect 26278 16990 26516 17086
rect 25738 16862 26516 16990
rect -1598 13600 -1472 13624
rect -1598 13166 -1570 13600
rect -1500 13166 -1472 13600
rect -1250 13620 -1146 13630
rect -1250 13186 -1234 13620
rect -1160 13186 -1146 13620
rect -1250 13168 -1146 13186
rect -930 13620 -826 13634
rect -930 13186 -916 13620
rect -842 13186 -826 13620
rect -930 13172 -826 13186
rect -566 13620 -440 13640
rect -566 13186 -544 13620
rect -474 13186 -440 13620
rect -1598 13138 -1472 13166
rect -1234 12904 -1154 13168
rect -918 12926 -838 13172
rect -566 13158 -440 13186
rect -1986 12850 -1148 12904
rect -918 12872 -78 12926
rect -1602 12016 -478 12060
rect -1602 12012 -912 12016
rect -1602 11574 -1550 12012
rect -1478 11574 -1224 12012
rect -1152 11578 -912 12012
rect -840 12008 -478 12016
rect -840 11578 -594 12008
rect -1152 11574 -594 11578
rect -1602 11570 -594 11574
rect -522 11570 -478 12008
rect -1602 11546 -478 11570
rect 23640 11114 24348 11166
rect 23640 10920 23814 11114
rect 24168 10920 24348 11114
rect 23640 10638 24348 10920
rect 23632 10594 24348 10638
rect 23638 10438 24348 10594
rect -1612 6854 -398 6888
rect -1612 6848 -594 6854
rect -2758 6484 -2650 6594
rect -2912 5644 -2852 6458
rect -2916 5440 -2852 5644
rect -6314 4882 -4476 5142
rect -6314 4154 -6072 4882
rect -4686 4154 -4476 4882
rect -6314 3912 -4476 4154
rect -2916 3946 -2856 5440
rect -2920 3760 -2856 3946
rect -2920 2494 -2860 3760
rect -2926 2062 -2860 2494
rect -2926 1506 -2866 2062
rect -2744 1896 -2650 6484
rect -1612 6410 -1550 6848
rect -1478 6410 -1234 6848
rect -1162 6410 -910 6848
rect -838 6446 -594 6848
rect -522 6446 -398 6854
rect -838 6434 -578 6446
rect -540 6434 -398 6446
rect -838 6410 -398 6434
rect -1612 6364 -398 6410
rect -2758 1708 -2650 1896
rect 23638 3916 24326 10438
rect 25740 5700 26512 16862
rect 51464 15844 53302 16112
rect 51464 15116 51706 15844
rect 53092 15116 53302 15844
rect 51464 14874 53302 15116
rect 51464 11844 53302 12112
rect 51464 11116 51706 11844
rect 53092 11116 53302 11844
rect 51464 10874 53302 11116
rect 51464 7844 53302 8112
rect 51464 7116 51706 7844
rect 53092 7116 53302 7844
rect 51464 6874 53302 7116
rect 23638 3648 23860 3916
rect 24124 3648 24326 3916
rect -6314 882 -4476 1142
rect -6314 154 -6072 882
rect -4686 154 -4476 882
rect -6314 -88 -4476 154
rect -2934 -998 -2862 1506
rect -2758 -404 -2664 1708
rect 23638 0 24326 3648
rect 26006 3658 26512 5700
rect 51464 3844 53302 4112
rect 31082 3716 31478 3820
rect 31082 3658 31166 3716
rect 26006 3616 31166 3658
rect 26006 0 26512 3616
rect 31082 3474 31166 3616
rect 31396 3474 31478 3716
rect 31082 3384 31478 3474
rect 51464 3116 51706 3844
rect 53092 3116 53302 3844
rect 51464 2874 53302 3116
rect 27708 1260 28132 1332
rect 27708 990 27780 1260
rect 28066 990 28132 1260
rect 27708 908 28132 990
rect -2766 -408 126 -404
rect 20652 -408 23544 -404
rect 26234 -408 26278 0
rect -2766 -412 4766 -408
rect 17860 -412 26280 -408
rect -2766 -416 7302 -412
rect 12342 -416 26280 -412
rect -2766 -458 26280 -416
rect -2758 -460 -2664 -458
rect -690 -462 20752 -458
rect 23388 -462 26280 -458
rect 498 -464 1172 -462
rect 4410 -466 17924 -462
rect 6816 -470 12456 -466
rect 27838 -998 28000 908
rect -2934 -1190 28000 -998
rect 51464 -156 53302 112
rect 51464 -884 51706 -156
rect 53092 -884 53302 -156
rect 51464 -1126 53302 -884
rect -2934 -1198 27984 -1190
rect -2934 -1200 536 -1198
rect 1076 -1200 27984 -1198
rect -3652 -2236 -1814 -1960
rect -3652 -2964 -3410 -2236
rect -2024 -2964 -1814 -2236
rect -3652 -3206 -1814 -2964
rect 348 -2060 536 -1964
rect 1076 -2060 2186 -1964
rect 348 -2236 2186 -2060
rect 348 -2964 590 -2236
rect 1976 -2964 2186 -2236
rect 348 -3206 2186 -2964
rect 4348 -2236 6186 -1964
rect 4348 -2964 4590 -2236
rect 5976 -2964 6186 -2236
rect 4348 -3206 6186 -2964
rect 8348 -2236 10186 -1964
rect 8348 -2964 8590 -2236
rect 9976 -2964 10186 -2236
rect 8348 -3206 10186 -2964
rect 12348 -2236 14186 -1964
rect 12348 -2964 12590 -2236
rect 13976 -2964 14186 -2236
rect 12348 -3206 14186 -2964
rect 16348 -2236 18186 -1964
rect 16348 -2964 16590 -2236
rect 17976 -2964 18186 -2236
rect 16348 -3206 18186 -2964
rect 20348 -2236 22186 -1964
rect 20348 -2964 20590 -2236
rect 21976 -2964 22186 -2236
rect 20348 -3206 22186 -2964
rect 24348 -2236 26186 -1964
rect 24348 -2964 24590 -2236
rect 25976 -2964 26186 -2236
rect 24348 -3206 26186 -2964
rect 28348 -2236 30186 -1964
rect 28348 -2964 28590 -2236
rect 29976 -2964 30186 -2236
rect 28348 -3206 30186 -2964
rect 32348 -2236 34186 -1964
rect 32348 -2964 32590 -2236
rect 33976 -2964 34186 -2236
rect 32348 -3206 34186 -2964
rect 36348 -2236 38186 -1964
rect 36348 -2964 36590 -2236
rect 37976 -2964 38186 -2236
rect 36348 -3206 38186 -2964
rect 40348 -2236 42186 -1964
rect 40348 -2964 40590 -2236
rect 41976 -2964 42186 -2236
rect 40348 -3206 42186 -2964
rect 44348 -2236 46186 -1964
rect 44348 -2964 44590 -2236
rect 45976 -2964 46186 -2236
rect 44348 -3206 46186 -2964
rect 48348 -2236 50186 -1964
rect 48348 -2964 48590 -2236
rect 49976 -2964 50186 -2236
rect 48348 -3206 50186 -2964
<< via1 >>
rect -4336 38318 -2950 39046
rect -336 38318 1050 39046
rect 3664 38318 5050 39046
rect 7664 38318 9050 39046
rect 11664 38318 13050 39046
rect 15664 38318 17050 39046
rect 19664 38318 21050 39046
rect 23664 38318 25050 39046
rect 27664 38318 29050 39046
rect 31664 38318 33050 39046
rect 35664 38318 37050 39046
rect 39664 38318 41050 39046
rect 43664 38318 45050 39046
rect 47664 38318 49050 39046
rect 51664 38318 53050 39046
rect -6072 36154 -4686 36882
rect 51706 35116 53092 35844
rect -6072 32154 -4686 32882
rect -1618 32518 -1542 32540
rect -1618 32121 -1598 32518
rect -1598 32121 -1560 32518
rect -1560 32121 -1542 32518
rect -1618 32104 -1542 32121
rect -1298 32518 -1222 32540
rect -1298 32121 -1280 32518
rect -1280 32121 -1242 32518
rect -1242 32121 -1222 32518
rect -1298 32104 -1222 32121
rect -982 32518 -906 32540
rect -982 32121 -962 32518
rect -962 32121 -924 32518
rect -924 32121 -906 32518
rect -982 32104 -906 32121
rect -662 32518 -586 32540
rect -662 32121 -644 32518
rect -644 32121 -606 32518
rect -606 32121 -586 32518
rect -662 32104 -586 32121
rect 51706 31116 53092 31844
rect -6072 28154 -4686 28882
rect -1614 27361 -1542 27378
rect -1614 26964 -1598 27361
rect -1598 26964 -1560 27361
rect -1560 26964 -1542 27361
rect -1614 26946 -1542 26964
rect -1298 27361 -1226 27378
rect -1298 26964 -1280 27361
rect -1280 26964 -1242 27361
rect -1242 26964 -1226 27361
rect -1298 26946 -1226 26964
rect -978 27361 -906 27378
rect -978 26964 -962 27361
rect -962 26964 -924 27361
rect -924 26964 -906 27361
rect -978 26946 -906 26964
rect -662 27361 -590 27378
rect -662 26964 -644 27361
rect -644 26964 -606 27361
rect -606 26964 -590 27361
rect -662 26946 -590 26964
rect 51706 27116 53092 27844
rect -6072 24154 -4686 24882
rect -1562 25240 -1490 25256
rect -1562 24843 -1546 25240
rect -1546 24843 -1508 25240
rect -1508 24843 -1490 25240
rect -1562 24824 -1490 24843
rect -492 25204 -420 25228
rect -492 24807 -474 25204
rect -474 24807 -436 25204
rect -436 24807 -420 25204
rect -492 24796 -420 24807
rect 51706 23116 53092 23844
rect -6072 20154 -4686 20882
rect -1564 20083 -1490 20100
rect -1564 19686 -1546 20083
rect -1546 19686 -1508 20083
rect -1508 19686 -1490 20083
rect -1564 19668 -1490 19686
rect -492 20047 -418 20060
rect -492 19650 -474 20047
rect -474 19650 -436 20047
rect -436 19650 -418 20047
rect -492 19628 -418 19650
rect -6072 16154 -4686 16882
rect -6072 12154 -4686 12882
rect -6072 8154 -4686 8882
rect -1572 18740 -1498 18764
rect -1572 18343 -1554 18740
rect -1554 18343 -1516 18740
rect -1516 18343 -1498 18740
rect -1572 18332 -1498 18343
rect 766 19018 954 19194
rect 3064 19246 3264 19480
rect 51706 19116 53092 19844
rect -548 18758 -474 18774
rect -548 18361 -528 18758
rect -528 18361 -490 18758
rect -490 18361 -474 18758
rect -548 18342 -474 18361
rect 26014 16990 26278 17086
rect -1570 13583 -1500 13600
rect -1570 13186 -1554 13583
rect -1554 13186 -1516 13583
rect -1516 13186 -1500 13583
rect -1570 13166 -1500 13186
rect -544 13601 -474 13620
rect -544 13204 -528 13601
rect -528 13204 -490 13601
rect -490 13204 -474 13601
rect -544 13186 -474 13204
rect -1550 11988 -1478 12012
rect -1550 11591 -1532 11988
rect -1532 11591 -1494 11988
rect -1494 11591 -1478 11988
rect -1550 11574 -1478 11591
rect -1224 11988 -1152 12012
rect -1224 11591 -1214 11988
rect -1214 11591 -1176 11988
rect -1176 11591 -1152 11988
rect -1224 11574 -1152 11591
rect -912 11988 -840 12016
rect -912 11591 -896 11988
rect -896 11591 -858 11988
rect -858 11591 -840 11988
rect -912 11578 -840 11591
rect -594 11988 -522 12008
rect -594 11591 -578 11988
rect -578 11591 -540 11988
rect -540 11591 -522 11988
rect -594 11570 -522 11591
rect 23814 10920 24168 11114
rect -6072 4154 -4686 4882
rect -1550 6831 -1478 6848
rect -1550 6434 -1532 6831
rect -1532 6434 -1494 6831
rect -1494 6434 -1478 6831
rect -1550 6410 -1478 6434
rect -1234 6831 -1162 6848
rect -1234 6434 -1214 6831
rect -1214 6434 -1176 6831
rect -1176 6434 -1162 6831
rect -1234 6410 -1162 6434
rect -910 6831 -838 6848
rect -910 6434 -896 6831
rect -896 6434 -858 6831
rect -858 6434 -838 6831
rect -594 6831 -522 6854
rect -594 6446 -578 6831
rect -578 6446 -540 6831
rect -540 6446 -522 6831
rect -910 6410 -838 6434
rect 51706 15116 53092 15844
rect 51706 11116 53092 11844
rect 51706 7116 53092 7844
rect 23860 3648 24124 3916
rect -6072 154 -4686 882
rect 31166 3474 31396 3716
rect 51706 3116 53092 3844
rect 27780 990 28066 1260
rect 51706 -884 53092 -156
rect -3410 -2964 -2024 -2236
rect 590 -2964 1976 -2236
rect 4590 -2964 5976 -2236
rect 8590 -2964 9976 -2236
rect 12590 -2964 13976 -2236
rect 16590 -2964 17976 -2236
rect 20590 -2964 21976 -2236
rect 24590 -2964 25976 -2236
rect 28590 -2964 29976 -2236
rect 32590 -2964 33976 -2236
rect 36590 -2964 37976 -2236
rect 40590 -2964 41976 -2236
rect 44590 -2964 45976 -2236
rect 48590 -2964 49976 -2236
<< metal2 >>
rect -4578 39046 -2740 39306
rect -4578 38318 -4336 39046
rect -2950 38318 -2740 39046
rect -4578 38076 -2740 38318
rect -578 39046 1260 39306
rect -578 38318 -336 39046
rect 1050 38318 1260 39046
rect -578 38076 1260 38318
rect 3422 39046 5260 39306
rect 3422 38318 3664 39046
rect 5050 38318 5260 39046
rect 3422 38076 5260 38318
rect 7422 39046 9260 39306
rect 7422 38318 7664 39046
rect 9050 38318 9260 39046
rect 7422 38076 9260 38318
rect 11422 39046 13260 39306
rect 11422 38318 11664 39046
rect 13050 38318 13260 39046
rect 11422 38076 13260 38318
rect 15422 39046 17260 39306
rect 15422 38318 15664 39046
rect 17050 38318 17260 39046
rect 15422 38076 17260 38318
rect 19422 39046 21260 39306
rect 19422 38318 19664 39046
rect 21050 38318 21260 39046
rect 19422 38076 21260 38318
rect 23422 39046 25260 39306
rect 23422 38318 23664 39046
rect 25050 38318 25260 39046
rect 23422 38076 25260 38318
rect 27422 39046 29260 39306
rect 27422 38318 27664 39046
rect 29050 38318 29260 39046
rect 27422 38076 29260 38318
rect 31422 39046 33260 39306
rect 31422 38318 31664 39046
rect 33050 38318 33260 39046
rect 31422 38076 33260 38318
rect 35422 39046 37260 39306
rect 35422 38318 35664 39046
rect 37050 38318 37260 39046
rect 35422 38076 37260 38318
rect 39422 39046 41260 39306
rect 39422 38318 39664 39046
rect 41050 38318 41260 39046
rect 39422 38076 41260 38318
rect 43422 39046 45260 39306
rect 43422 38318 43664 39046
rect 45050 38318 45260 39046
rect 43422 38076 45260 38318
rect 47422 39046 49260 39306
rect 47422 38318 47664 39046
rect 49050 38318 49260 39046
rect 47422 38076 49260 38318
rect 51422 39046 53260 39306
rect 51422 38318 51664 39046
rect 53050 38318 53260 39046
rect 51422 38076 53260 38318
rect -6314 36882 -4476 37142
rect -6314 36154 -6072 36882
rect -4686 36154 -4476 36882
rect -6314 35912 -4476 36154
rect 14330 35820 37810 36672
rect 51464 35844 53302 36112
rect 14330 35298 37902 35820
rect -6314 32882 -4476 33142
rect -6314 32154 -6072 32882
rect -4686 32154 -4476 32882
rect -6314 31912 -4476 32154
rect -1820 32540 -252 32556
rect -1820 32104 -1618 32540
rect -1542 32104 -1298 32540
rect -1222 32104 -982 32540
rect -906 32104 -662 32540
rect -586 32104 -252 32540
rect -6314 28882 -4476 29142
rect -6314 28154 -6072 28882
rect -4686 28154 -4476 28882
rect -6314 27912 -4476 28154
rect -1820 27378 -252 32104
rect -1820 26946 -1614 27378
rect -1542 26946 -1298 27378
rect -1226 26946 -978 27378
rect -906 26946 -662 27378
rect -590 26946 -252 27378
rect -1820 25256 -252 26946
rect -6314 24882 -4476 25142
rect -6314 24154 -6072 24882
rect -4686 24154 -4476 24882
rect -6314 23912 -4476 24154
rect -1820 24824 -1562 25256
rect -1490 25228 -252 25256
rect 14382 27834 15684 35298
rect 36600 34958 37902 35298
rect 20486 34724 32738 34858
rect 20486 33932 31362 34724
rect 32478 33932 32738 34724
rect 20486 33800 32738 33932
rect 36600 34170 36834 34958
rect 37692 34170 37902 34958
rect 51464 35116 51706 35844
rect 53092 35116 53302 35844
rect 51464 34874 53302 35116
rect 20492 27852 21684 33800
rect 14382 27814 15686 27834
rect 14382 27742 15030 27814
rect 15192 27742 15686 27814
rect 14382 26378 15686 27742
rect 20492 27780 20926 27852
rect 21088 27780 21684 27852
rect 20492 27740 21684 27780
rect 31304 27860 32496 33800
rect 31304 27788 31818 27860
rect 31980 27788 32496 27860
rect 14382 25626 14628 26378
rect 15310 25626 15686 26378
rect 14382 25416 15686 25626
rect 20418 26050 21694 27740
rect 20418 25836 20920 26050
rect 21178 25836 21694 26050
rect 14382 25238 15684 25416
rect 20418 25322 21694 25836
rect 31304 26908 32496 27788
rect 31304 25444 31502 26908
rect 32464 25444 32496 26908
rect -1490 24824 -492 25228
rect -1820 24796 -492 24824
rect -420 24796 -252 25228
rect 20492 25104 21684 25322
rect 31304 25058 32496 25444
rect 36600 27784 37902 34170
rect 51464 31844 53302 32112
rect 51464 31116 51706 31844
rect 53092 31116 53302 31844
rect 51464 30874 53302 31116
rect 36600 27712 37088 27784
rect 37250 27712 37902 27784
rect 36600 27160 37902 27712
rect 36600 25696 36784 27160
rect 37746 25696 37902 27160
rect 51464 27844 53302 28112
rect 51464 27116 51706 27844
rect 53092 27116 53302 27844
rect 51464 26874 53302 27116
rect 36600 25306 37902 25696
rect -6314 20882 -4476 21142
rect -6314 20154 -6072 20882
rect -4686 20154 -4476 20882
rect -6314 19912 -4476 20154
rect -1820 20100 -252 24796
rect 51464 23844 53302 24112
rect 51464 23116 51706 23844
rect 53092 23116 53302 23844
rect 51464 22874 53302 23116
rect -1820 19668 -1564 20100
rect -1490 20060 -252 20100
rect -1490 19668 -492 20060
rect -1820 19628 -492 19668
rect -418 19628 -252 20060
rect -1820 18774 -252 19628
rect 14398 21696 15818 21966
rect 14398 20232 14588 21696
rect 15550 20232 15818 21696
rect 28398 21692 31114 21868
rect 20118 21330 20766 21554
rect 3028 19480 3308 19568
rect 718 19194 996 19296
rect 718 19018 766 19194
rect 954 19018 996 19194
rect 3028 19246 3064 19480
rect 3264 19246 3308 19480
rect 3028 19170 3308 19246
rect 718 18930 996 19018
rect -1820 18764 -548 18774
rect -1820 18332 -1572 18764
rect -1498 18342 -548 18764
rect -474 18342 -252 18774
rect -1498 18332 -252 18342
rect -6314 16882 -4476 17142
rect -6314 16154 -6072 16882
rect -4686 16154 -4476 16882
rect -6314 15912 -4476 16154
rect -1820 13620 -252 18332
rect -1820 13600 -544 13620
rect -1820 13166 -1570 13600
rect -1500 13186 -544 13600
rect -474 13186 -252 13620
rect -1500 13166 -252 13186
rect -6314 12882 -4476 13142
rect -6314 12154 -6072 12882
rect -4686 12154 -4476 12882
rect -6314 11912 -4476 12154
rect -1820 12016 -252 13166
rect -1820 12012 -912 12016
rect -1820 11574 -1550 12012
rect -1478 11574 -1224 12012
rect -1152 11578 -912 12012
rect -840 12008 -252 12016
rect -840 11578 -594 12008
rect -1152 11574 -594 11578
rect -1820 11570 -594 11574
rect -522 11570 -252 12008
rect -6314 8882 -4476 9142
rect -6314 8154 -6072 8882
rect -4686 8154 -4476 8882
rect -6314 7912 -4476 8154
rect -1820 6854 -252 11570
rect 14398 17050 15818 20232
rect 20624 19866 20766 21330
rect 20118 18846 20766 19866
rect 28398 21422 31968 21692
rect 28398 19958 31114 21422
rect 31848 19958 31968 21422
rect 28398 19126 31968 19958
rect 14398 16978 15150 17050
rect 15312 16978 15818 17050
rect 6252 10758 7870 11032
rect 6252 9960 6468 10758
rect 7658 9960 7870 10758
rect 6252 9744 7870 9960
rect -1820 6848 -594 6854
rect -1820 6410 -1550 6848
rect -1478 6410 -1234 6848
rect -1162 6410 -910 6848
rect -838 6446 -594 6848
rect -522 6446 -252 6854
rect -838 6410 -252 6446
rect -1820 5540 -252 6410
rect 6378 6592 6454 9744
rect 14398 9112 15818 16978
rect 19552 17120 20766 18846
rect 19552 17048 20076 17120
rect 20238 17048 20766 17120
rect 19552 10306 20766 17048
rect 25966 17086 26342 17130
rect 25966 16990 26014 17086
rect 26278 16990 26342 17086
rect 25966 16962 26342 16990
rect 30754 16972 31968 19126
rect 30754 16900 31346 16972
rect 31508 16900 31968 16972
rect 23602 11114 24522 11192
rect 23602 10920 23814 11114
rect 24168 10920 24522 11114
rect 23602 10888 24522 10920
rect 30754 10306 31968 16900
rect 36344 21606 37764 21874
rect 36344 20142 36508 21606
rect 37470 20142 37764 21606
rect 36344 17060 37764 20142
rect 51464 19844 53302 20112
rect 51464 19116 51706 19844
rect 53092 19116 53302 19844
rect 51464 18874 53302 19116
rect 36344 16988 36870 17060
rect 37032 16988 37764 17060
rect 14394 8906 15818 9112
rect 14394 7974 14662 8906
rect 15370 8588 15818 8906
rect 19530 9884 32060 10306
rect 19530 8768 30570 9884
rect 31732 8768 32060 9884
rect 15370 7974 15796 8588
rect 19530 8520 32060 8768
rect 36344 8998 37764 16988
rect 51464 15844 53302 16112
rect 51464 15116 51706 15844
rect 53092 15116 53302 15844
rect 51464 14874 53302 15116
rect 51464 11844 53302 12112
rect 51464 11116 51706 11844
rect 53092 11116 53302 11844
rect 51464 10874 53302 11116
rect 36344 8496 37796 8998
rect 14394 7572 15796 7974
rect 36394 7572 37796 8496
rect 51464 7844 53302 8112
rect -6314 4882 -4476 5142
rect -6314 4154 -6072 4882
rect -4686 4154 -4476 4882
rect -6314 3912 -4476 4154
rect -6314 882 -4476 1142
rect -6314 154 -6072 882
rect -4686 154 -4476 882
rect -6314 -88 -4476 154
rect -3652 -2236 -1814 -1960
rect -3652 -2964 -3410 -2236
rect -2024 -2538 -1814 -2236
rect -1672 -2538 -1500 5540
rect 6378 4684 6450 6592
rect 14188 6260 37958 7572
rect 51464 7116 51706 7844
rect 53092 7116 53302 7844
rect 51464 6874 53302 7116
rect 36394 6192 37796 6260
rect 6378 4618 6452 4684
rect 6380 3644 6452 4618
rect 23778 3916 24190 3986
rect 23778 3648 23860 3916
rect 24124 3648 24190 3916
rect 51464 3844 53302 4112
rect 6380 3586 6454 3644
rect 6382 2634 6454 3586
rect 23778 3582 24190 3648
rect 31082 3716 31478 3820
rect 31082 3474 31166 3716
rect 31396 3474 31478 3716
rect 31082 3384 31478 3474
rect 51464 3116 51706 3844
rect 53092 3116 53302 3844
rect 51464 2874 53302 3116
rect 6382 2546 6458 2634
rect 6386 -508 6458 2546
rect 27708 1260 28132 1332
rect 27708 990 27780 1260
rect 28066 990 28132 1260
rect 27708 908 28132 990
rect 6384 -564 6458 -508
rect 51464 -156 53302 112
rect 6384 -1534 6456 -564
rect 51464 -884 51706 -156
rect 53092 -884 53302 -156
rect 51464 -1126 53302 -884
rect 6384 -1606 6460 -1534
rect -2024 -2608 -1500 -2538
rect -2024 -2964 -1814 -2608
rect -1672 -2636 -1500 -2608
rect 348 -2060 536 -1964
rect 1076 -2060 2186 -1964
rect 348 -2236 2186 -2060
rect -3652 -3206 -1814 -2964
rect 348 -2964 590 -2236
rect 1976 -2964 2186 -2236
rect 348 -3206 2186 -2964
rect 4348 -2236 6186 -1964
rect 4348 -2964 4590 -2236
rect 5976 -2562 6186 -2236
rect 6388 -2562 6460 -1606
rect 8348 -2236 10186 -1964
rect 5976 -2620 6466 -2562
rect 5976 -2964 6186 -2620
rect 6388 -2632 6460 -2620
rect 4348 -3206 6186 -2964
rect 8348 -2964 8590 -2236
rect 9976 -2964 10186 -2236
rect 8348 -3206 10186 -2964
rect 12348 -2236 14186 -1964
rect 12348 -2964 12590 -2236
rect 13976 -2964 14186 -2236
rect 12348 -3206 14186 -2964
rect 16348 -2236 18186 -1964
rect 16348 -2964 16590 -2236
rect 17976 -2964 18186 -2236
rect 16348 -3206 18186 -2964
rect 20348 -2236 22186 -1964
rect 20348 -2964 20590 -2236
rect 21976 -2964 22186 -2236
rect 20348 -3206 22186 -2964
rect 24348 -2236 26186 -1964
rect 24348 -2964 24590 -2236
rect 25976 -2964 26186 -2236
rect 24348 -3206 26186 -2964
rect 28348 -2236 30186 -1964
rect 28348 -2964 28590 -2236
rect 29976 -2964 30186 -2236
rect 28348 -3206 30186 -2964
rect 32348 -2236 34186 -1964
rect 32348 -2964 32590 -2236
rect 33976 -2964 34186 -2236
rect 32348 -3206 34186 -2964
rect 36348 -2236 38186 -1964
rect 36348 -2964 36590 -2236
rect 37976 -2964 38186 -2236
rect 36348 -3206 38186 -2964
rect 40348 -2236 42186 -1964
rect 40348 -2964 40590 -2236
rect 41976 -2964 42186 -2236
rect 40348 -3206 42186 -2964
rect 44348 -2236 46186 -1964
rect 44348 -2964 44590 -2236
rect 45976 -2964 46186 -2236
rect 44348 -3206 46186 -2964
rect 48348 -2236 50186 -1964
rect 48348 -2964 48590 -2236
rect 49976 -2964 50186 -2236
rect 48348 -3206 50186 -2964
<< via2 >>
rect -4336 38318 -2950 39046
rect -336 38318 1050 39046
rect 3664 38318 5050 39046
rect 7664 38318 9050 39046
rect 11664 38318 13050 39046
rect 15664 38318 17050 39046
rect 19664 38318 21050 39046
rect 23664 38318 25050 39046
rect 27664 38318 29050 39046
rect 31664 38318 33050 39046
rect 35664 38318 37050 39046
rect 39664 38318 41050 39046
rect 43664 38318 45050 39046
rect 47664 38318 49050 39046
rect 51664 38318 53050 39046
rect -6072 36154 -4686 36882
rect -6072 32154 -4686 32882
rect -6072 28154 -4686 28882
rect -6072 24154 -4686 24882
rect 31362 33932 32478 34724
rect 36834 34170 37692 34958
rect 51706 35116 53092 35844
rect 15030 27742 15192 27814
rect 20926 27780 21088 27852
rect 31818 27788 31980 27860
rect 51706 31116 53092 31844
rect 37088 27712 37250 27784
rect 51706 27116 53092 27844
rect -6072 20154 -4686 20882
rect 51706 23116 53092 23844
rect 766 19018 954 19194
rect 3064 19246 3264 19480
rect -6072 16154 -4686 16882
rect -6072 12154 -4686 12882
rect -6072 8154 -4686 8882
rect 15150 16978 15312 17050
rect 6468 9960 7658 10758
rect 20076 17048 20238 17120
rect 26014 16990 26278 17086
rect 31346 16900 31508 16972
rect 23814 10920 24168 11114
rect 51706 19116 53092 19844
rect 36870 16988 37032 17060
rect 14662 7974 15370 8906
rect 30570 8768 31732 9884
rect 51706 15116 53092 15844
rect 51706 11116 53092 11844
rect -6072 4154 -4686 4882
rect -6072 154 -4686 882
rect -3410 -2964 -2024 -2236
rect 51706 7116 53092 7844
rect 23860 3648 24124 3916
rect 31166 3474 31396 3716
rect 51706 3116 53092 3844
rect 27780 990 28066 1260
rect 51706 -884 53092 -156
rect 590 -2964 1976 -2236
rect 4590 -2964 5976 -2236
rect 8590 -2964 9976 -2236
rect 12590 -2964 13976 -2236
rect 16590 -2964 17976 -2236
rect 20590 -2964 21976 -2236
rect 24590 -2964 25976 -2236
rect 28590 -2964 29976 -2236
rect 32590 -2964 33976 -2236
rect 36590 -2964 37976 -2236
rect 40590 -2964 41976 -2236
rect 44590 -2964 45976 -2236
rect 48590 -2964 49976 -2236
<< metal3 >>
rect -4578 39046 -2740 39306
rect -4578 38318 -4336 39046
rect -2950 38318 -2740 39046
rect -4578 38076 -2740 38318
rect -578 39046 1260 39306
rect -578 38318 -336 39046
rect 1050 38318 1260 39046
rect -578 38076 1260 38318
rect 3422 39046 5260 39306
rect 3422 38318 3664 39046
rect 5050 38318 5260 39046
rect 3422 38076 5260 38318
rect 7422 39046 9260 39306
rect 7422 38318 7664 39046
rect 9050 38318 9260 39046
rect 7422 38076 9260 38318
rect 11422 39046 13260 39306
rect 11422 38318 11664 39046
rect 13050 38318 13260 39046
rect 11422 38076 13260 38318
rect 15422 39046 17260 39306
rect 15422 38318 15664 39046
rect 17050 38318 17260 39046
rect 15422 38076 17260 38318
rect 19422 39046 21260 39306
rect 19422 38318 19664 39046
rect 21050 38318 21260 39046
rect 19422 38076 21260 38318
rect 23422 39046 25260 39306
rect 23422 38318 23664 39046
rect 25050 38318 25260 39046
rect 23422 38076 25260 38318
rect 27422 39046 29260 39306
rect 27422 38318 27664 39046
rect 29050 38318 29260 39046
rect 27422 38076 29260 38318
rect 31422 39046 33260 39306
rect 31422 38318 31664 39046
rect 33050 38318 33260 39046
rect 31422 38076 33260 38318
rect 35422 39046 37260 39306
rect 35422 38318 35664 39046
rect 37050 38318 37260 39046
rect 35422 38076 37260 38318
rect 39422 39046 41260 39306
rect 39422 38318 39664 39046
rect 41050 38318 41260 39046
rect 39422 38076 41260 38318
rect 43422 39046 45260 39306
rect 43422 38318 43664 39046
rect 45050 38318 45260 39046
rect 43422 38076 45260 38318
rect 47422 39046 49260 39306
rect 47422 38318 47664 39046
rect 49050 38318 49260 39046
rect 47422 38076 49260 38318
rect 51422 39046 53260 39306
rect 51422 38318 51664 39046
rect 53050 38318 53260 39046
rect 51422 38076 53260 38318
rect -6314 36882 -4476 37142
rect -6314 36154 -6072 36882
rect -4686 36154 -4476 36882
rect -6314 35912 -4476 36154
rect 51464 35844 53302 36112
rect 36672 35094 46902 35120
rect 51464 35116 51706 35844
rect 53092 35116 53302 35844
rect 36672 34958 46990 35094
rect 0 34724 33188 34856
rect 0 33932 31362 34724
rect 32478 33932 33188 34724
rect 36672 34170 36834 34958
rect 37692 34170 46990 34958
rect 51464 34874 53302 35116
rect 36672 34076 46990 34170
rect 0 33594 33188 33932
rect -6314 32882 -4476 33142
rect -6314 32154 -6072 32882
rect -4686 32154 -4476 32882
rect -6314 31912 -4476 32154
rect -6314 28882 -4476 29142
rect -6314 28154 -6072 28882
rect -4686 28154 -4476 28882
rect -6314 27912 -4476 28154
rect -6314 24882 -4476 25142
rect -6314 24154 -6072 24882
rect -4686 24154 -4476 24882
rect -6314 23912 -4476 24154
rect -6314 20882 -4476 21142
rect -6314 20154 -6072 20882
rect -4686 20154 -4476 20882
rect -6314 19912 -4476 20154
rect 280 19194 1588 33594
rect 5807 28154 44028 33272
rect 5807 28152 31194 28154
rect 5807 28122 20600 28152
rect 5807 28000 14682 28122
rect 15572 28000 20600 28122
rect 21502 28000 31194 28152
rect 32828 28102 44028 28154
rect 32828 28000 36796 28102
rect 37708 28000 44028 28102
rect 280 19018 766 19194
rect 954 19018 1588 19194
rect 3028 19480 3308 19568
rect 3028 19246 3064 19480
rect 3264 19246 3308 19480
rect 3028 19170 3308 19246
rect -6314 16882 -4476 17142
rect -6314 16154 -6072 16882
rect -4686 16154 -4476 16882
rect -6314 15912 -4476 16154
rect -6314 12882 -4476 13142
rect -6314 12154 -6072 12882
rect -4686 12154 -4476 12882
rect -6314 11912 -4476 12154
rect -6314 8882 -4476 9142
rect -6314 8154 -6072 8882
rect -4686 8154 -4476 8882
rect -6314 7912 -4476 8154
rect 280 5452 1588 19018
rect 5840 16566 10947 28000
rect 20902 27852 21120 27882
rect 15006 27814 15224 27844
rect 20902 27824 20926 27852
rect 15006 27786 15030 27814
rect 15004 27742 15030 27786
rect 15192 27742 15224 27814
rect 15004 27684 15224 27742
rect 20900 27780 20926 27824
rect 21088 27780 21120 27852
rect 31794 27860 32012 27890
rect 31794 27832 31818 27860
rect 20900 27684 21120 27780
rect 31792 27788 31818 27832
rect 31980 27788 32012 27860
rect 31792 27724 32012 27788
rect 37064 27784 37282 27814
rect 37064 27756 37088 27784
rect 11344 27546 16390 27684
rect 11344 22670 16394 27546
rect 16868 27530 21914 27684
rect 16868 24252 21928 27530
rect 11344 22566 16390 22670
rect 16868 22566 21914 24252
rect 22373 22566 27419 27684
rect 27857 22606 32903 27724
rect 37062 27712 37088 27756
rect 37250 27712 37282 27784
rect 37062 27684 37282 27712
rect 38789 27684 43896 28000
rect 33382 22566 38428 27684
rect 38789 22566 43928 27684
rect 22414 22148 27388 22566
rect 16850 22095 21836 22108
rect 11446 17050 16432 22048
rect 16850 17120 21920 22095
rect 16850 17082 20076 17120
rect 11446 17022 15150 17050
rect 15124 16978 15150 17022
rect 15312 17022 16432 17050
rect 20050 17048 20076 17082
rect 20238 17082 21920 17120
rect 22414 17122 27401 22148
rect 22414 17094 27388 17122
rect 27917 17103 32903 22208
rect 38789 22128 43896 22566
rect 27917 17102 32784 17103
rect 20238 17048 20270 17082
rect 21581 17080 21920 17082
rect 25682 17086 26728 17094
rect 15312 16978 15344 17022
rect 15124 16902 15344 16978
rect 20050 16972 20270 17048
rect 25682 16990 26014 17086
rect 26278 16990 26728 17086
rect 25682 16938 26728 16990
rect 31314 16972 31572 17102
rect 33382 17060 38428 22128
rect 33382 17022 36870 17060
rect 31314 16926 31346 16972
rect 31320 16900 31346 16926
rect 31508 16926 31572 16972
rect 36844 16988 36870 17022
rect 37032 17022 38428 17060
rect 38789 17022 43928 22128
rect 37032 16988 37064 17022
rect 31508 16900 31540 16926
rect 36844 16912 37064 16988
rect 31320 16824 31540 16900
rect 11344 16566 16390 16584
rect 16868 16566 21914 16584
rect 22373 16566 27419 16584
rect 27857 16566 31014 16624
rect 5741 16534 31014 16566
rect 31938 16566 32903 16624
rect 38789 16584 43896 17022
rect 33382 16566 38428 16584
rect 38789 16566 43928 16584
rect 31938 16534 43928 16566
rect 5741 11472 43928 16534
rect 5741 11327 43896 11472
rect 6240 10758 7896 11327
rect 23602 11114 24522 11192
rect 23602 10920 23814 11114
rect 24168 10920 24522 11114
rect 23602 10888 24522 10920
rect 6240 9960 6468 10758
rect 7658 9960 7896 10758
rect 30570 10116 32058 10256
rect 6240 9746 7896 9960
rect 30246 9884 32058 10116
rect 6252 9744 7870 9746
rect 14402 8906 15928 9464
rect 14402 7974 14662 8906
rect 15370 7974 15928 8906
rect 30246 8768 30570 9884
rect 31732 8768 32058 9884
rect 30246 8198 32058 8768
rect 14402 5452 15928 7974
rect 30264 5480 31790 8198
rect 44804 7094 46990 34076
rect 51464 31844 53302 32112
rect 51464 31116 51706 31844
rect 53092 31116 53302 31844
rect 51464 30874 53302 31116
rect 51464 27844 53302 28112
rect 51464 27116 51706 27844
rect 53092 27116 53302 27844
rect 51464 26874 53302 27116
rect 51464 23844 53302 24112
rect 51464 23116 51706 23844
rect 53092 23116 53302 23844
rect 51464 22874 53302 23116
rect 51464 19844 53302 20112
rect 51464 19116 51706 19844
rect 53092 19116 53302 19844
rect 51464 18874 53302 19116
rect 51464 15844 53302 16112
rect 51464 15116 51706 15844
rect 53092 15116 53302 15844
rect 51464 14874 53302 15116
rect 51464 11844 53302 12112
rect 51464 11116 51706 11844
rect 53092 11116 53302 11844
rect 51464 10874 53302 11116
rect 51464 7844 53302 8112
rect 51464 7116 51706 7844
rect 53092 7116 53302 7844
rect 24120 5452 25896 5480
rect -6314 4882 -4476 5142
rect -6314 4154 -6072 4882
rect -4686 4154 -4476 4882
rect 280 4472 25896 5452
rect -6314 3912 -4476 4154
rect 374 3916 25896 4472
rect 374 3648 23860 3916
rect 24124 3676 25896 3916
rect 30246 4674 32058 5480
rect 44664 4674 47036 7094
rect 51464 6874 53302 7116
rect 30246 3716 47036 4674
rect 24124 3648 25848 3676
rect 374 3116 25848 3648
rect 30246 3474 31166 3716
rect 31396 3474 47036 3716
rect 30246 2814 47036 3474
rect 51464 3844 53302 4112
rect 51464 3116 51706 3844
rect 53092 3116 53302 3844
rect 51464 2874 53302 3116
rect 44664 2768 47036 2814
rect 27708 1260 28132 1332
rect -6314 882 -4476 1142
rect 27708 990 27780 1260
rect 28066 990 28132 1260
rect 27708 908 28132 990
rect -6314 154 -6072 882
rect -4686 154 -4476 882
rect -6314 -88 -4476 154
rect 51464 -156 53302 112
rect 51464 -884 51706 -156
rect 53092 -884 53302 -156
rect 51464 -1126 53302 -884
rect -3652 -2236 -1814 -1960
rect -3652 -2964 -3410 -2236
rect -2024 -2964 -1814 -2236
rect -3652 -3206 -1814 -2964
rect 348 -2060 536 -1964
rect 1076 -2060 2186 -1964
rect 348 -2236 2186 -2060
rect 348 -2964 590 -2236
rect 1976 -2964 2186 -2236
rect 348 -3206 2186 -2964
rect 4348 -2236 6186 -1964
rect 4348 -2964 4590 -2236
rect 5976 -2964 6186 -2236
rect 4348 -3206 6186 -2964
rect 8348 -2236 10186 -1964
rect 8348 -2964 8590 -2236
rect 9976 -2964 10186 -2236
rect 8348 -3206 10186 -2964
rect 12348 -2236 14186 -1964
rect 12348 -2964 12590 -2236
rect 13976 -2964 14186 -2236
rect 12348 -3206 14186 -2964
rect 16348 -2236 18186 -1964
rect 16348 -2964 16590 -2236
rect 17976 -2964 18186 -2236
rect 16348 -3206 18186 -2964
rect 20348 -2236 22186 -1964
rect 20348 -2964 20590 -2236
rect 21976 -2964 22186 -2236
rect 20348 -3206 22186 -2964
rect 24348 -2236 26186 -1964
rect 24348 -2964 24590 -2236
rect 25976 -2964 26186 -2236
rect 24348 -3206 26186 -2964
rect 28348 -2236 30186 -1964
rect 28348 -2964 28590 -2236
rect 29976 -2964 30186 -2236
rect 28348 -3206 30186 -2964
rect 32348 -2236 34186 -1964
rect 32348 -2964 32590 -2236
rect 33976 -2964 34186 -2236
rect 32348 -3206 34186 -2964
rect 36348 -2236 38186 -1964
rect 36348 -2964 36590 -2236
rect 37976 -2964 38186 -2236
rect 36348 -3206 38186 -2964
rect 40348 -2236 42186 -1964
rect 40348 -2964 40590 -2236
rect 41976 -2964 42186 -2236
rect 40348 -3206 42186 -2964
rect 44348 -2236 46186 -1964
rect 44348 -2964 44590 -2236
rect 45976 -2964 46186 -2236
rect 44348 -3206 46186 -2964
rect 48348 -2236 50186 -1964
rect 48348 -2964 48590 -2236
rect 49976 -2964 50186 -2236
rect 48348 -3206 50186 -2964
<< via3 >>
rect -4336 38318 -2950 39046
rect -336 38318 1050 39046
rect 3664 38318 5050 39046
rect 7664 38318 9050 39046
rect 11664 38318 13050 39046
rect 15664 38318 17050 39046
rect 19664 38318 21050 39046
rect 23664 38318 25050 39046
rect 27664 38318 29050 39046
rect 31664 38318 33050 39046
rect 35664 38318 37050 39046
rect 39664 38318 41050 39046
rect 43664 38318 45050 39046
rect 47664 38318 49050 39046
rect 51664 38318 53050 39046
rect -6072 36154 -4686 36882
rect 51706 35116 53092 35844
rect -6072 32154 -4686 32882
rect -6072 28154 -4686 28882
rect -6072 24154 -4686 24882
rect -6072 20154 -4686 20882
rect 3064 19246 3264 19480
rect -6072 16154 -4686 16882
rect -6072 12154 -4686 12882
rect -6072 8154 -4686 8882
rect 23814 10920 24168 11114
rect 6468 9960 7658 10758
rect 51706 31116 53092 31844
rect 51706 27116 53092 27844
rect 51706 23116 53092 23844
rect 51706 19116 53092 19844
rect 51706 15116 53092 15844
rect 51706 11116 53092 11844
rect 51706 7116 53092 7844
rect -6072 4154 -4686 4882
rect 51706 3116 53092 3844
rect 27780 990 28066 1260
rect -6072 154 -4686 882
rect 51706 -884 53092 -156
rect -3410 -2964 -2024 -2236
rect 590 -2964 1976 -2236
rect 4590 -2964 5976 -2236
rect 8590 -2964 9976 -2236
rect 12590 -2964 13976 -2236
rect 16590 -2964 17976 -2236
rect 20590 -2964 21976 -2236
rect 24590 -2964 25976 -2236
rect 28590 -2964 29976 -2236
rect 32590 -2964 33976 -2236
rect 36590 -2964 37976 -2236
rect 40590 -2964 41976 -2236
rect 44590 -2964 45976 -2236
rect 48590 -2964 49976 -2236
<< mimcap >>
rect 5986 31297 10786 33030
rect 5986 29675 6505 31297
rect 7769 29675 10786 31297
rect 5986 28204 10786 29675
rect 11566 31141 16366 33018
rect 11566 29679 14368 31141
rect 15763 29679 16366 31141
rect 11566 28198 16366 29679
rect 17066 31229 21866 33018
rect 17066 29767 20215 31229
rect 21610 29767 21866 31229
rect 17066 28198 21866 29767
rect 22566 31340 27366 33018
rect 22566 29878 25353 31340
rect 26748 29878 27366 31340
rect 22566 28198 27366 29878
rect 28066 31362 32866 33018
rect 28066 29900 31001 31362
rect 32396 29900 32866 31362
rect 28066 28198 32866 29900
rect 33566 31340 38366 33018
rect 33566 29878 36516 31340
rect 37911 29878 38366 31340
rect 33566 28198 38366 29878
rect 39066 31296 43866 33018
rect 39066 29834 39395 31296
rect 40790 29834 43866 31296
rect 39066 28198 43866 29834
rect 5986 25797 10786 27530
rect 5986 24175 6511 25797
rect 7769 24175 10786 25797
rect 5986 22698 10786 24175
rect 11566 25218 16366 27518
rect 11566 24140 12062 25218
rect 13168 24140 16366 25218
rect 11566 22698 16366 24140
rect 17066 26856 21866 27518
rect 17066 26760 17816 26856
rect 17066 25242 18938 26760
rect 17066 25110 17816 25242
rect 19002 25110 21866 26856
rect 17066 22698 21866 25110
rect 22566 24502 27366 27518
rect 22566 23288 23642 24502
rect 25588 23288 27366 24502
rect 22566 22698 27366 23288
rect 28066 27152 32866 27518
rect 28066 25406 28892 27152
rect 30078 26826 32866 27152
rect 28958 25406 32866 26826
rect 28066 22698 32866 25406
rect 33566 25554 38366 27518
rect 33566 24604 34112 25554
rect 35398 24604 38366 25554
rect 33566 22698 38366 24604
rect 39066 24829 43866 27518
rect 39066 23367 39572 24829
rect 40967 23367 43866 24829
rect 39066 22698 43866 23367
rect 5986 20297 10786 22018
rect 5986 18675 6511 20297
rect 7769 18675 10786 20297
rect 5986 17198 10786 18675
rect 11566 21582 16366 22018
rect 11566 21518 12178 21582
rect 11566 20064 13334 21518
rect 11566 20000 13300 20064
rect 13398 20000 16366 21582
rect 11566 19802 12178 20000
rect 13364 19802 16366 20000
rect 11566 17198 16366 19802
rect 17066 21310 21866 22018
rect 17066 19960 17882 21310
rect 18848 19960 21866 21310
rect 17066 17198 21866 19960
rect 22566 21178 27366 22018
rect 22566 19964 23618 21178
rect 23718 19964 25260 21050
rect 25564 19964 27366 21178
rect 22566 17198 27366 19964
rect 28066 21538 32866 22018
rect 28066 20240 29004 21538
rect 30224 20240 32866 21538
rect 28066 17198 32866 20240
rect 33566 21812 38366 22018
rect 33566 20066 34530 21812
rect 35716 21682 38366 21812
rect 34596 20164 38366 21682
rect 35716 20066 38366 20164
rect 33566 17198 38366 20066
rect 39066 20200 43866 22018
rect 39066 18738 39661 20200
rect 41056 18738 43866 20200
rect 39066 17198 43866 18738
rect 5986 14797 10786 16430
rect 5986 13175 6511 14797
rect 7769 13175 10786 14797
rect 5986 11604 10786 13175
rect 11486 14797 16286 16430
rect 11486 13175 12011 14797
rect 13269 13175 16286 14797
rect 11486 11604 16286 13175
rect 16986 14797 21786 16430
rect 16986 13175 17511 14797
rect 18769 13175 21786 14797
rect 16986 11604 21786 13175
rect 22486 14797 27286 16430
rect 22486 13175 23011 14797
rect 24269 13175 27286 14797
rect 22486 11604 27286 13175
rect 27986 14797 32786 16430
rect 27986 13175 28511 14797
rect 29769 13175 32786 14797
rect 27986 11604 32786 13175
rect 33486 14797 38286 16430
rect 33486 13175 34011 14797
rect 35269 13175 38286 14797
rect 33486 11604 38286 13175
rect 38986 14797 43786 16430
rect 38986 13175 39511 14797
rect 40769 13175 43786 14797
rect 38986 11604 43786 13175
<< mimcapcontact >>
rect 6505 29675 7769 31297
rect 14368 29679 15763 31141
rect 20215 29767 21610 31229
rect 25353 29878 26748 31340
rect 31001 29900 32396 31362
rect 36516 29878 37911 31340
rect 39395 29834 40790 31296
rect 6511 24175 7769 25797
rect 12062 24140 13168 25218
rect 17816 26760 19002 26856
rect 18938 25242 19002 26760
rect 17816 25110 19002 25242
rect 23642 23288 25588 24502
rect 28892 26826 30078 27152
rect 28892 25406 28958 26826
rect 34112 24604 35398 25554
rect 39572 23367 40967 24829
rect 6511 18675 7769 20297
rect 12178 21518 13398 21582
rect 13334 20064 13398 21518
rect 13300 20000 13398 20064
rect 12178 19802 13364 20000
rect 17882 19960 18848 21310
rect 23618 21050 25564 21178
rect 23618 19964 23718 21050
rect 25260 19964 25564 21050
rect 29004 20240 30224 21538
rect 34530 21682 35716 21812
rect 34530 20164 34596 21682
rect 34530 20066 35716 20164
rect 39661 18738 41056 20200
rect 6511 13175 7769 14797
rect 12011 13175 13269 14797
rect 17511 13175 18769 14797
rect 23011 13175 24269 14797
rect 28511 13175 29769 14797
rect 34011 13175 35269 14797
rect 39511 13175 40769 14797
<< metal4 >>
rect -4578 39046 -2740 39306
rect -4578 38318 -4336 39046
rect -2950 38318 -2740 39046
rect -4578 38076 -2740 38318
rect -578 39046 1260 39306
rect -578 38318 -336 39046
rect 1050 38318 1260 39046
rect -578 38076 1260 38318
rect 3422 39046 5260 39306
rect 3422 38318 3664 39046
rect 5050 38318 5260 39046
rect 3422 38076 5260 38318
rect 7422 39046 9260 39306
rect 7422 38318 7664 39046
rect 9050 38318 9260 39046
rect 7422 38076 9260 38318
rect 11422 39046 13260 39306
rect 11422 38318 11664 39046
rect 13050 38318 13260 39046
rect 11422 38076 13260 38318
rect 15422 39046 17260 39306
rect 15422 38318 15664 39046
rect 17050 38318 17260 39046
rect 15422 38076 17260 38318
rect 19422 39046 21260 39306
rect 19422 38318 19664 39046
rect 21050 38318 21260 39046
rect 19422 38076 21260 38318
rect 23422 39046 25260 39306
rect 23422 38318 23664 39046
rect 25050 38318 25260 39046
rect 23422 38076 25260 38318
rect 27422 39046 29260 39306
rect 27422 38318 27664 39046
rect 29050 38318 29260 39046
rect 27422 38076 29260 38318
rect 31422 39046 33260 39306
rect 31422 38318 31664 39046
rect 33050 38318 33260 39046
rect 31422 38076 33260 38318
rect 35422 39046 37260 39306
rect 35422 38318 35664 39046
rect 37050 38318 37260 39046
rect 35422 38076 37260 38318
rect 39422 39046 41260 39306
rect 39422 38318 39664 39046
rect 41050 38318 41260 39046
rect 39422 38076 41260 38318
rect 43422 39046 45260 39306
rect 43422 38318 43664 39046
rect 45050 38318 45260 39046
rect 43422 38076 45260 38318
rect 47422 39046 49260 39306
rect 47422 38318 47664 39046
rect 49050 38318 49260 39046
rect 47422 38076 49260 38318
rect 51422 39046 53260 39306
rect 51422 38318 51664 39046
rect 53050 38318 53260 39046
rect 51422 38076 53260 38318
rect -6314 36882 -4476 37142
rect -6314 36154 -6072 36882
rect -4686 36154 -4476 36882
rect 43222 36512 50344 36536
rect -6314 35912 -4476 36154
rect 33632 36416 50344 36512
rect 33632 35678 33836 36416
rect 35314 35678 50344 36416
rect 33632 35512 50344 35678
rect 33632 35468 43862 35512
rect 46664 35420 50344 35512
rect 51464 35844 53302 36112
rect 2710 34856 4018 34902
rect 2646 34635 19258 34856
rect 2646 33997 18009 34635
rect 18778 33997 19258 34635
rect 2646 33546 19258 33997
rect -6314 32882 -4476 33142
rect -6314 32154 -6072 32882
rect -4686 32154 -4476 32882
rect -6314 31912 -4476 32154
rect -6314 28882 -4476 29142
rect -6314 28154 -6072 28882
rect -4686 28154 -4476 28882
rect -6314 27912 -4476 28154
rect -6314 24882 -4476 25142
rect -6314 24154 -6072 24882
rect -4686 24154 -4476 24882
rect -6314 23912 -4476 24154
rect -6314 20882 -4476 21142
rect -6314 20154 -6072 20882
rect -4686 20154 -4476 20882
rect -6314 19912 -4476 20154
rect 2710 19480 4018 33546
rect 2710 19246 3064 19480
rect 3264 19246 4018 19480
rect -6314 16882 -4476 17142
rect -6314 16154 -6072 16882
rect -4686 16154 -4476 16882
rect -6314 15912 -4476 16154
rect -6314 12882 -4476 13142
rect -6314 12154 -6072 12882
rect -4686 12154 -4476 12882
rect -6314 11912 -4476 12154
rect -6314 8882 -4476 9142
rect -6314 8154 -6072 8882
rect -4686 8154 -4476 8882
rect -6314 7912 -4476 8154
rect 2710 7984 4018 19246
rect 6306 31662 7962 31695
rect 6306 31629 41045 31662
rect 6306 31362 41111 31629
rect 6306 31340 31001 31362
rect 6306 31297 25353 31340
rect 6306 29675 6505 31297
rect 7769 31229 25353 31297
rect 7769 31141 20215 31229
rect 7769 29679 14368 31141
rect 15763 29767 20215 31141
rect 21610 29878 25353 31229
rect 26748 29900 31001 31340
rect 32396 31340 41111 31362
rect 32396 29900 36516 31340
rect 26748 29878 36516 29900
rect 37911 31296 41111 31340
rect 37911 29878 39395 31296
rect 21610 29834 39395 29878
rect 40790 29834 41111 31296
rect 21610 29767 41111 29834
rect 15763 29679 41111 29767
rect 7769 29675 41111 29679
rect 6306 29410 41111 29675
rect 6306 25797 7962 29410
rect 6306 24175 6511 25797
rect 7769 24175 7962 25797
rect 6306 20297 7962 24175
rect 11754 26840 13604 27302
rect 17690 27026 19173 27287
rect 11754 25734 12138 26840
rect 13140 25734 13604 26840
rect 11754 25218 13604 25734
rect 11754 24140 12062 25218
rect 13168 24140 13604 25218
rect 17602 26856 19173 27026
rect 17602 26760 17816 26856
rect 17602 25242 17750 26760
rect 17602 25110 17816 25242
rect 19002 25110 19173 26856
rect 17602 24728 19173 25110
rect 28738 27152 30221 27229
rect 28738 25406 28892 27152
rect 30078 26826 30221 27152
rect 28738 25308 28958 25406
rect 30146 25308 30221 26826
rect 17602 24467 19085 24728
rect 23352 24502 25994 24768
rect 28738 24670 30221 25308
rect 33778 27020 35654 27534
rect 33778 26222 34344 27020
rect 35088 26222 35654 27020
rect 33778 25554 35654 26222
rect 11754 23910 13604 24140
rect 23352 23288 23642 24502
rect 25588 23288 25994 24502
rect 33778 24604 34112 25554
rect 35398 24604 35654 25554
rect 33778 23986 35654 24604
rect 39290 24829 41111 29410
rect 23352 22496 25994 23288
rect 39290 23367 39572 24829
rect 40967 23367 41111 24829
rect 23352 22112 25840 22496
rect 6306 18675 6511 20297
rect 7769 18675 7962 20297
rect 11618 21582 13992 22012
rect 23352 21824 25994 22112
rect 11618 21518 12178 21582
rect 11618 20000 12146 21518
rect 13398 20000 13992 21582
rect 11618 19802 12178 20000
rect 13364 19802 13992 20000
rect 17626 21310 19408 21792
rect 23352 21646 25818 21824
rect 17626 19960 17882 21310
rect 18848 19960 19408 21310
rect 11991 19233 13474 19802
rect 17626 19730 19408 19960
rect 17576 19630 19408 19730
rect 23300 21178 25818 21646
rect 23300 19964 23618 21178
rect 23300 19724 23718 19964
rect 25564 19964 25818 21178
rect 25260 19724 25818 19964
rect 6306 15137 7962 18675
rect 17576 18714 19358 19630
rect 23300 19326 25818 19724
rect 28646 21538 30632 21818
rect 28646 20240 29004 21538
rect 30224 20240 30632 21538
rect 17576 17822 18034 18714
rect 18696 17822 19358 18714
rect 17576 17568 19358 17822
rect 28646 18944 30632 20240
rect 34134 21812 36508 21846
rect 34134 20066 34530 21812
rect 35716 21682 36508 21812
rect 35784 20164 36508 21682
rect 35716 20066 36508 20164
rect 34134 19636 36508 20066
rect 39290 20200 41111 23367
rect 34408 19175 35891 19636
rect 28646 18052 28978 18944
rect 29640 18052 30632 18944
rect 28646 17772 30632 18052
rect 39290 18738 39661 20200
rect 41056 18738 41111 20200
rect 39290 15137 41111 18738
rect 6240 14797 41276 15137
rect 6240 13175 6511 14797
rect 7769 13175 12011 14797
rect 13269 13175 17511 14797
rect 18769 13175 23011 14797
rect 24269 13175 28511 14797
rect 29769 13175 34011 14797
rect 35269 13175 39511 14797
rect 40769 13175 41276 14797
rect 6240 12786 41276 13175
rect 6240 10758 7896 12786
rect 39290 12686 41111 12786
rect 23602 11156 24522 11192
rect 23602 10920 23814 11156
rect 24168 10920 24522 11156
rect 23602 10888 24522 10920
rect 6240 9960 6468 10758
rect 7658 9960 7896 10758
rect 6240 9746 7896 9960
rect 17640 9884 19222 10116
rect 17640 8768 17920 9884
rect 19082 8768 19222 9884
rect 17640 8396 19222 8768
rect 2416 6316 4120 7984
rect 10586 6762 13696 7042
rect 10586 6316 12480 6762
rect 2416 5826 12480 6316
rect 13508 5826 13696 6762
rect 2416 5594 13696 5826
rect -6314 4882 -4476 5142
rect -6314 4154 -6072 4882
rect -4686 4154 -4476 4882
rect 2416 4484 4120 5594
rect -6314 3912 -4476 4154
rect 17640 3512 19128 8396
rect 17454 2164 19128 3512
rect 47966 2164 50292 35420
rect 51464 35116 51706 35844
rect 53092 35116 53302 35844
rect 51464 34874 53302 35116
rect 51464 31844 53302 32112
rect 51464 31116 51706 31844
rect 53092 31116 53302 31844
rect 51464 30874 53302 31116
rect 51464 27844 53302 28112
rect 51464 27116 51706 27844
rect 53092 27116 53302 27844
rect 51464 26874 53302 27116
rect 51464 23844 53302 24112
rect 51464 23116 51706 23844
rect 53092 23116 53302 23844
rect 51464 22874 53302 23116
rect 51464 19844 53302 20112
rect 51464 19116 51706 19844
rect 53092 19116 53302 19844
rect 51464 18874 53302 19116
rect 51464 15844 53302 16112
rect 51464 15116 51706 15844
rect 53092 15116 53302 15844
rect 51464 14874 53302 15116
rect 51464 11844 53302 12112
rect 51464 11116 51706 11844
rect 53092 11116 53302 11844
rect 51464 10874 53302 11116
rect 51464 7844 53302 8112
rect 51464 7116 51706 7844
rect 53092 7116 53302 7844
rect 51464 6874 53302 7116
rect 51464 3844 53302 4112
rect 51464 3116 51706 3844
rect 53092 3116 53302 3844
rect 51464 2874 53302 3116
rect 17454 1260 50292 2164
rect -6314 882 -4476 1142
rect -6314 154 -6072 882
rect -4686 154 -4476 882
rect 17454 990 27780 1260
rect 28066 990 50292 1260
rect 17454 488 50292 990
rect 47966 350 50292 488
rect -6314 -88 -4476 154
rect 51464 -156 53302 112
rect 51464 -884 51706 -156
rect 53092 -884 53302 -156
rect 51464 -1126 53302 -884
rect -3652 -2236 -1814 -1960
rect -3652 -2964 -3410 -2236
rect -2024 -2964 -1814 -2236
rect -3652 -3206 -1814 -2964
rect 348 -2060 536 -1964
rect 1076 -2060 2186 -1964
rect 348 -2236 2186 -2060
rect 348 -2964 590 -2236
rect 1976 -2964 2186 -2236
rect 348 -3206 2186 -2964
rect 4348 -2236 6186 -1964
rect 4348 -2964 4590 -2236
rect 5976 -2964 6186 -2236
rect 4348 -3206 6186 -2964
rect 8348 -2236 10186 -1964
rect 8348 -2964 8590 -2236
rect 9976 -2964 10186 -2236
rect 8348 -3206 10186 -2964
rect 12348 -2236 14186 -1964
rect 12348 -2964 12590 -2236
rect 13976 -2964 14186 -2236
rect 12348 -3206 14186 -2964
rect 16348 -2236 18186 -1964
rect 16348 -2964 16590 -2236
rect 17976 -2964 18186 -2236
rect 16348 -3206 18186 -2964
rect 20348 -2236 22186 -1964
rect 20348 -2964 20590 -2236
rect 21976 -2964 22186 -2236
rect 20348 -3206 22186 -2964
rect 24348 -2236 26186 -1964
rect 24348 -2964 24590 -2236
rect 25976 -2964 26186 -2236
rect 24348 -3206 26186 -2964
rect 28348 -2236 30186 -1964
rect 28348 -2964 28590 -2236
rect 29976 -2964 30186 -2236
rect 28348 -3206 30186 -2964
rect 32348 -2236 34186 -1964
rect 32348 -2964 32590 -2236
rect 33976 -2964 34186 -2236
rect 32348 -3206 34186 -2964
rect 36348 -2236 38186 -1964
rect 36348 -2964 36590 -2236
rect 37976 -2964 38186 -2236
rect 36348 -3206 38186 -2964
rect 40348 -2236 42186 -1964
rect 40348 -2964 40590 -2236
rect 41976 -2964 42186 -2236
rect 40348 -3206 42186 -2964
rect 44348 -2236 46186 -1964
rect 44348 -2964 44590 -2236
rect 45976 -2964 46186 -2236
rect 44348 -3206 46186 -2964
rect 48348 -2236 50186 -1964
rect 48348 -2964 48590 -2236
rect 49976 -2964 50186 -2236
rect 48348 -3206 50186 -2964
<< via4 >>
rect 33836 35678 35314 36416
rect 18009 33997 18778 34635
rect 12138 25734 13140 26840
rect 17750 25242 18938 26760
rect 28958 25308 30146 26826
rect 34344 26222 35088 27020
rect 12146 20064 13334 21518
rect 12146 20000 13300 20064
rect 23718 19724 25260 21050
rect 18034 17822 18696 18714
rect 34596 20164 35784 21682
rect 28978 18052 29640 18944
rect 23814 11114 24168 11156
rect 23814 10920 24168 11114
rect 17920 8768 19082 9884
rect 12480 5826 13508 6762
<< metal5 >>
rect 12016 36416 35496 36672
rect 12016 35678 33836 36416
rect 35314 35706 35496 36416
rect 35314 35678 35524 35706
rect 12016 35298 35524 35678
rect 12050 27918 13352 35298
rect 17682 34702 29934 34880
rect 17682 34635 30114 34702
rect 17682 33997 18009 34635
rect 18778 33997 30114 34635
rect 17682 33822 30114 33997
rect 17766 33800 19130 33822
rect 11908 26840 13474 27918
rect 17766 27287 18958 33800
rect 17690 27114 19173 27287
rect 28922 27229 30114 33822
rect 34222 29770 35524 35298
rect 33778 29436 35524 29770
rect 11908 25734 12138 26840
rect 13140 25734 13474 26840
rect 11908 25400 13474 25734
rect 17532 26760 19344 27114
rect 17532 25242 17750 26760
rect 18938 25242 19344 26760
rect 17532 25140 19344 25242
rect 28738 26826 30221 27229
rect 28738 25308 28958 26826
rect 30146 25308 30221 26826
rect 33778 27020 35474 29436
rect 33778 26222 34344 27020
rect 35088 26222 35474 27020
rect 33778 26042 35474 26222
rect 17690 24728 19173 25140
rect 28738 24670 30221 25308
rect 11991 21762 13474 21792
rect 11830 21518 13642 21762
rect 11830 20000 12146 21518
rect 13334 20064 13642 21518
rect 34374 21682 36186 21920
rect 13300 20000 13642 20064
rect 11830 19788 13642 20000
rect 23326 21050 25362 21304
rect 11991 19233 13474 19788
rect 23326 19724 23718 21050
rect 25260 19724 25362 21050
rect 34374 20164 34596 21682
rect 35784 20164 36186 21682
rect 34374 19946 36186 20164
rect 12040 9202 13460 19233
rect 23326 19112 25362 19724
rect 34408 19494 35891 19946
rect 34396 19175 35891 19494
rect 17812 18714 19026 18846
rect 23326 18738 24906 19112
rect 17812 17822 18034 18714
rect 18696 17822 19026 18714
rect 23314 18112 24906 18738
rect 28778 18944 30038 19126
rect 17812 10260 19026 17822
rect 23376 11262 24816 18112
rect 28778 18072 28978 18944
rect 28808 18052 28978 18072
rect 29640 18072 30038 18944
rect 29640 18052 30022 18072
rect 23364 11156 24826 11262
rect 23364 10920 23814 11156
rect 24168 10920 24826 11156
rect 23364 10818 24826 10920
rect 28808 10260 30022 18052
rect 17744 9884 30068 10260
rect 12040 8268 13474 9202
rect 17744 8768 17920 9884
rect 19082 8768 30068 9884
rect 17744 8382 30068 8768
rect 34396 8538 35816 19175
rect 12072 7066 13474 8268
rect 34370 8314 35816 8538
rect 34370 7066 35772 8314
rect 12072 6762 35888 7066
rect 12072 5826 12480 6762
rect 13508 5826 35888 6762
rect 12072 5800 35888 5826
rect 12118 5754 35888 5800
rect 34370 5732 35772 5754
<< res0p35 >>
rect -1616 27376 -1542 32106
rect -1298 27376 -1224 32106
rect -980 27376 -906 32106
rect -662 27376 -588 32106
rect -1564 20098 -1490 24828
rect -1208 20080 -1134 24810
rect -890 20080 -816 24810
rect -492 20062 -418 24792
rect -1572 13598 -1498 18328
rect -1234 13618 -1160 18348
rect -916 13618 -842 18348
rect -546 13616 -472 18346
rect -1550 6846 -1476 11576
rect -1232 6846 -1158 11576
rect -914 6846 -840 11576
rect -596 6846 -522 11576
<< labels >>
flabel metal1 -842 25434 -842 25434 0 FreeSans 1600 0 0 0 vbias1
flabel metal1 -1178 25364 -1178 25364 0 FreeSans 1600 0 0 0 vbias2
flabel psubdiff -686 -2644 -686 -2644 0 FreeSans 1600 0 0 0 gnd
flabel metal3 46068 9984 46068 9984 0 FreeSans 1600 0 0 0 Bot_2
flabel metal4 49000 9040 49000 9040 0 FreeSans 1600 0 0 0 Top_2
flabel metal3 856 17074 856 17074 0 FreeSans 1600 0 0 0 Bot_1
flabel metal4 3404 17130 3404 17130 0 FreeSans 1600 0 0 0 Top_1
flabel metal1 -168 12900 -168 12900 0 FreeSans 1600 0 0 0 vinp2
flabel metal1 -1922 12880 -1922 12880 0 FreeSans 1600 0 0 0 vinp1
<< end >>
