magic
tech sky130A
magscale 1 2
timestamp 1634727530
<< nwell >>
rect -34584 18420 376 18716
rect -34584 17392 384 18420
rect -34584 520 376 17392
rect -34702 388 376 520
rect -34722 258 376 388
rect -34722 254 314 258
rect -34722 -262 272 254
rect -34722 -922 -506 -262
rect 54 -346 248 -262
rect -34586 -924 -506 -922
<< psubdiff >>
rect -62 -694 542 -678
rect -62 -746 -30 -694
rect 28 -746 370 -694
rect 428 -746 542 -694
rect -62 -760 542 -746
<< nsubdiff >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
<< psubdiffcont >>
rect -30 -746 28 -694
rect 370 -746 428 -694
<< nsubdiffcont >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
<< locali >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -32416 426 -31428 17046
rect -30764 426 -29776 17116
rect -29158 426 -28170 17046
rect -27458 426 -26470 17116
rect -25830 426 -24842 17092
rect -24154 426 -23166 17116
rect -22502 426 -21514 17070
rect -20872 426 -19884 17092
rect -19220 426 -18232 17070
rect -17520 426 -16532 17092
rect -15962 460 -14974 17092
rect -15962 426 -14964 460
rect -14214 426 -13226 17116
rect -12562 426 -11574 17116
rect -10932 426 -9944 17116
rect -9254 426 -8266 17116
rect -7556 426 -6568 17092
rect -5926 426 -4938 17140
rect -4250 426 -3262 17116
rect -2598 426 -1610 17140
rect -968 428 20 17116
rect -968 426 -4 428
rect -32422 388 -4 426
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -748 346 -4 388
rect -748 312 -72 346
rect -36 340 -4 346
rect -36 312 -2 340
rect -748 274 -2 312
rect 132 198 198 254
rect 380 134 448 158
rect -34586 -54 -734 116
rect 380 98 394 134
rect 432 98 448 134
rect 380 82 448 98
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect 130 -290 198 -276
rect 130 -334 138 -290
rect 184 -334 198 -290
rect 130 -342 198 -334
rect -34586 -828 -734 -520
rect -62 -694 542 -678
rect -62 -746 -30 -694
rect 28 -746 370 -694
rect 428 -746 542 -694
rect -62 -760 542 -746
<< viali >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -72 312 -36 346
rect 394 98 432 134
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 138 -334 184 -290
rect -30 -746 28 -694
rect 370 -746 428 -694
<< metal1 >>
rect 860 350192 1240 350420
rect -34456 18152 -32822 18174
rect -34456 18134 -328 18152
rect -34456 17946 372 18134
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 372 17946
rect -34456 17406 372 17480
rect -34456 17378 -32822 17406
rect -358 17400 372 17406
rect -34456 17376 -33498 17378
rect -358 17376 376 17400
rect -34456 15946 -33510 17376
rect 176 16710 376 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -32980 634 376 16710
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -90 372 -4 388
rect -92 346 130 372
rect -92 312 -72 346
rect -36 312 130 346
rect -92 280 130 312
rect -90 272 -12 280
rect -68 270 -18 272
rect -34586 -54 -734 116
rect 54 54 130 280
rect 380 134 610 156
rect 380 98 394 134
rect 432 98 610 134
rect 380 88 610 98
rect 230 58 266 60
rect 342 58 362 60
rect 230 56 362 58
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect 56 -26 138 54
rect 230 50 392 56
rect 226 48 392 50
rect 56 -90 72 -26
rect 128 -90 138 -26
rect 56 -142 138 -90
rect 190 -138 392 48
rect 438 -12 520 58
rect 438 -76 454 -12
rect 510 -76 520 -12
rect 438 -138 520 -76
rect 224 -140 392 -138
rect 288 -180 328 -140
rect 286 -226 330 -180
rect 126 -290 196 -280
rect 126 -334 138 -290
rect 184 -334 196 -290
rect 286 -296 934 -226
rect 288 -298 934 -296
rect 126 -444 196 -334
rect -34586 -828 -734 -520
rect -62 -694 542 -678
rect -62 -746 -30 -694
rect 28 -746 370 -694
rect 428 -746 542 -694
rect -62 -760 542 -746
<< via1 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 72 -90 128 -26
rect 454 -76 510 -12
rect -30 -746 28 -694
rect 370 -746 428 -694
<< metal2 >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect 54 -12 520 60
rect 54 -26 454 -12
rect 54 -90 72 -26
rect 128 -76 454 -26
rect 510 -76 520 -12
rect 128 -90 520 -76
rect 54 -142 520 -90
rect 56 -144 138 -142
rect -34586 -828 -734 -520
rect -62 -690 542 -678
rect -62 -746 -30 -690
rect 28 -746 370 -690
rect 428 -746 542 -690
rect -62 -760 542 -746
<< via2 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect -30 -694 28 -690
rect -30 -746 28 -694
rect 370 -694 428 -690
rect 370 -746 428 -694
<< metal3 >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
rect -62 -682 542 -678
rect -62 -746 -30 -682
rect 34 -746 370 -682
rect 434 -746 542 -682
rect -62 -760 542 -746
<< via3 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect -30 -690 34 -682
rect -30 -746 28 -690
rect 28 -746 34 -690
rect 370 -690 434 -682
rect 370 -746 428 -690
rect 428 -746 434 -690
<< metal4 >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
rect -62 -682 542 -678
rect -62 -746 -30 -682
rect 34 -746 370 -682
rect 434 -746 542 -682
rect -62 -760 542 -746
<< via4 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
<< metal5 >>
rect -34456 18152 -32822 18174
rect -34456 17946 -328 18152
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -328 17946
rect -34456 17406 -328 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 384 -33510 1480
rect -34586 116 -33510 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
use sky130_fd_pr__pfet_01v8_NZGT56  sky130_fd_pr__pfet_01v8_NZGT56_0
timestamp 1634714564
transform 1 0 163 0 1 -46
box -109 -300 109 300
use sky130_fd_pr__nfet_01v8_A8TGU8  sky130_fd_pr__nfet_01v8_A8TGU8_0
timestamp 1634714564
transform 1 0 413 0 1 -40
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_lvt_9PNB2P  sky130_fd_pr__pfet_01v8_lvt_9PNB2P_0
timestamp 1634714564
transform 1 0 -16337 0 1 3894
box -16645 -3254 16645 3254
use sky130_fd_pr__pfet_01v8_lvt_9PNB2P  sky130_fd_pr__pfet_01v8_lvt_9PNB2P_1
timestamp 1634714564
transform 1 0 -16335 0 1 10446
box -16645 -3254 16645 3254
use sky130_fd_pr__pfet_01v8_9PNB23  sky130_fd_pr__pfet_01v8_9PNB23_0
timestamp 1634714564
transform 1 0 -16341 0 1 15400
box -16645 -1618 16645 1618
use sky130_fd_pr__res_xhigh_po_0p35_Q5JWWA  sky130_fd_pr__res_xhigh_po_0p35_Q5JWWA_0
timestamp 1634716072
transform 1 0 896 0 1 175057
box -201 -175598 201 175598
<< labels >>
flabel metal1 56 314 56 314 0 FreeSans 320 0 0 0 net1
flabel metal1 1154 350306 1154 350306 0 FreeSans 320 0 0 0 GND!
flabel metal4 182 -728 182 -728 0 FreeSans 320 0 0 0 GND!
flabel metal1 228 17518 228 17518 0 FreeSans 320 0 0 0 VDD!
flabel metal1 536 116 536 116 0 FreeSans 320 0 0 0 clkb_in
flabel metal1 158 -422 158 -422 0 FreeSans 320 0 0 0 clk_in
flabel metal1 558 -270 558 -270 0 FreeSans 320 0 0 0 net2
<< end >>
