magic
tech sky130A
magscale 1 2
timestamp 1634911627
<< nwell >>
rect -804 1892 1298 1894
rect -804 514 6150 1892
rect -128 470 6150 514
rect -128 400 5162 470
rect 5940 468 6150 470
rect -128 390 94 400
rect 384 398 5162 400
rect 394 396 4120 398
rect 4776 396 5162 398
rect 394 392 1366 396
rect 2014 394 3454 396
rect 394 390 1062 392
rect 2990 390 3454 394
rect 932 -778 2152 -738
rect 930 -1284 2152 -778
rect 932 -1286 2152 -1284
rect 932 -1288 2120 -1286
rect 932 -1646 2090 -1288
rect 932 -2640 2088 -1646
rect 932 -3000 2084 -2640
<< nmos >>
rect 174 80 204 228
rect 270 80 300 228
rect 786 88 816 236
rect 882 88 912 236
rect 1364 84 1394 232
rect 1460 84 1490 232
rect 1938 92 1968 240
rect 2034 92 2064 240
rect 2516 92 2546 240
rect 2612 92 2642 240
rect 3094 92 3124 240
rect 3190 92 3220 240
rect 3676 96 3706 244
rect 3772 96 3802 244
rect 4252 92 4282 240
rect 4348 92 4378 240
rect 4822 88 4852 236
rect 4918 88 4948 236
rect 2232 -2258 2262 -1610
rect 2328 -2258 2358 -1610
rect 2424 -2258 2454 -1610
rect 2520 -2258 2550 -1610
rect 2616 -2258 2646 -1610
rect 2712 -2258 2742 -1610
rect 2808 -2258 2838 -1610
rect 2904 -2258 2934 -1610
rect 3000 -2258 3030 -1610
<< pmos >>
rect 170 490 200 826
rect 374 528 404 864
rect 782 498 812 834
rect 986 536 1016 872
rect 1360 494 1390 830
rect 1564 532 1594 868
rect 1934 502 1964 838
rect 2138 540 2168 876
rect 2512 502 2542 838
rect 2716 540 2746 876
rect 3090 502 3120 838
rect 3294 540 3324 876
rect 3672 506 3702 842
rect 3876 544 3906 880
rect 4248 502 4278 838
rect 4452 540 4482 876
rect 4818 498 4848 834
rect 5022 536 5052 872
rect 1564 -1564 1594 -1228
rect 1764 -1526 1794 -1190
rect 1966 -1566 1996 -1230
rect 1564 -2070 1594 -1734
rect 1764 -2032 1794 -1696
rect 1964 -2070 1994 -1734
rect 1564 -2578 1594 -2242
rect 1764 -2540 1794 -2204
rect 1964 -2578 1994 -2242
<< ndiff >>
rect 112 216 174 228
rect 112 92 124 216
rect 158 92 174 216
rect 112 80 174 92
rect 204 216 270 228
rect 204 92 220 216
rect 254 92 270 216
rect 204 80 270 92
rect 300 216 362 228
rect 300 92 316 216
rect 350 92 362 216
rect 300 80 362 92
rect 724 224 786 236
rect 724 100 736 224
rect 770 100 786 224
rect 724 88 786 100
rect 816 224 882 236
rect 816 100 832 224
rect 866 100 882 224
rect 816 88 882 100
rect 912 224 974 236
rect 912 100 928 224
rect 962 100 974 224
rect 912 88 974 100
rect 1302 220 1364 232
rect 1302 96 1314 220
rect 1348 96 1364 220
rect 1302 84 1364 96
rect 1394 220 1460 232
rect 1394 96 1410 220
rect 1444 96 1460 220
rect 1394 84 1460 96
rect 1490 220 1552 232
rect 1490 96 1506 220
rect 1540 96 1552 220
rect 1490 84 1552 96
rect 1876 228 1938 240
rect 1876 104 1888 228
rect 1922 104 1938 228
rect 1876 92 1938 104
rect 1968 228 2034 240
rect 1968 104 1984 228
rect 2018 104 2034 228
rect 1968 92 2034 104
rect 2064 228 2126 240
rect 2064 104 2080 228
rect 2114 104 2126 228
rect 2064 92 2126 104
rect 2454 228 2516 240
rect 2454 104 2466 228
rect 2500 104 2516 228
rect 2454 92 2516 104
rect 2546 228 2612 240
rect 2546 104 2562 228
rect 2596 104 2612 228
rect 2546 92 2612 104
rect 2642 228 2704 240
rect 2642 104 2658 228
rect 2692 104 2704 228
rect 2642 92 2704 104
rect 3032 228 3094 240
rect 3032 104 3044 228
rect 3078 104 3094 228
rect 3032 92 3094 104
rect 3124 228 3190 240
rect 3124 104 3140 228
rect 3174 104 3190 228
rect 3124 92 3190 104
rect 3220 228 3282 240
rect 3220 104 3236 228
rect 3270 104 3282 228
rect 3220 92 3282 104
rect 3614 232 3676 244
rect 3614 108 3626 232
rect 3660 108 3676 232
rect 3614 96 3676 108
rect 3706 232 3772 244
rect 3706 108 3722 232
rect 3756 108 3772 232
rect 3706 96 3772 108
rect 3802 232 3864 244
rect 3802 108 3818 232
rect 3852 108 3864 232
rect 3802 96 3864 108
rect 4190 228 4252 240
rect 4190 104 4202 228
rect 4236 104 4252 228
rect 4190 92 4252 104
rect 4282 228 4348 240
rect 4282 104 4298 228
rect 4332 104 4348 228
rect 4282 92 4348 104
rect 4378 228 4440 240
rect 4378 104 4394 228
rect 4428 104 4440 228
rect 4378 92 4440 104
rect 4760 224 4822 236
rect 4760 100 4772 224
rect 4806 100 4822 224
rect 4760 88 4822 100
rect 4852 224 4918 236
rect 4852 100 4868 224
rect 4902 100 4918 224
rect 4852 88 4918 100
rect 4948 224 5010 236
rect 4948 100 4964 224
rect 4998 100 5010 224
rect 4948 88 5010 100
rect 2170 -1622 2232 -1610
rect 2170 -2246 2182 -1622
rect 2216 -2246 2232 -1622
rect 2170 -2258 2232 -2246
rect 2262 -1622 2328 -1610
rect 2262 -2246 2278 -1622
rect 2312 -2246 2328 -1622
rect 2262 -2258 2328 -2246
rect 2358 -1622 2424 -1610
rect 2358 -2246 2374 -1622
rect 2408 -2246 2424 -1622
rect 2358 -2258 2424 -2246
rect 2454 -1622 2520 -1610
rect 2454 -2246 2470 -1622
rect 2504 -2246 2520 -1622
rect 2454 -2258 2520 -2246
rect 2550 -1622 2616 -1610
rect 2550 -2246 2566 -1622
rect 2600 -2246 2616 -1622
rect 2550 -2258 2616 -2246
rect 2646 -1622 2712 -1610
rect 2646 -2246 2662 -1622
rect 2696 -2246 2712 -1622
rect 2646 -2258 2712 -2246
rect 2742 -1622 2808 -1610
rect 2742 -2246 2758 -1622
rect 2792 -2246 2808 -1622
rect 2742 -2258 2808 -2246
rect 2838 -1622 2904 -1610
rect 2838 -2246 2854 -1622
rect 2888 -2246 2904 -1622
rect 2838 -2258 2904 -2246
rect 2934 -1622 3000 -1610
rect 2934 -2246 2950 -1622
rect 2984 -2246 3000 -1622
rect 2934 -2258 3000 -2246
rect 3030 -1622 3092 -1610
rect 3030 -2246 3046 -1622
rect 3080 -2246 3092 -1622
rect 3030 -2258 3092 -2246
<< pdiff >>
rect 316 852 374 864
rect 112 814 170 826
rect 112 502 124 814
rect 158 502 170 814
rect 112 490 170 502
rect 200 814 258 826
rect 200 502 212 814
rect 246 502 258 814
rect 316 540 328 852
rect 362 540 374 852
rect 316 528 374 540
rect 404 852 462 864
rect 404 540 416 852
rect 450 540 462 852
rect 928 860 986 872
rect 404 528 462 540
rect 724 822 782 834
rect 200 490 258 502
rect 724 510 736 822
rect 770 510 782 822
rect 724 498 782 510
rect 812 822 870 834
rect 812 510 824 822
rect 858 510 870 822
rect 928 548 940 860
rect 974 548 986 860
rect 928 536 986 548
rect 1016 860 1074 872
rect 1016 548 1028 860
rect 1062 548 1074 860
rect 1506 856 1564 868
rect 1016 536 1074 548
rect 1302 818 1360 830
rect 812 498 870 510
rect 1302 506 1314 818
rect 1348 506 1360 818
rect 1302 494 1360 506
rect 1390 818 1448 830
rect 1390 506 1402 818
rect 1436 506 1448 818
rect 1506 544 1518 856
rect 1552 544 1564 856
rect 1506 532 1564 544
rect 1594 856 1652 868
rect 1594 544 1606 856
rect 1640 544 1652 856
rect 2080 864 2138 876
rect 1594 532 1652 544
rect 1876 826 1934 838
rect 1390 494 1448 506
rect 1876 514 1888 826
rect 1922 514 1934 826
rect 1876 502 1934 514
rect 1964 826 2022 838
rect 1964 514 1976 826
rect 2010 514 2022 826
rect 2080 552 2092 864
rect 2126 552 2138 864
rect 2080 540 2138 552
rect 2168 864 2226 876
rect 2168 552 2180 864
rect 2214 552 2226 864
rect 2658 864 2716 876
rect 2168 540 2226 552
rect 2454 826 2512 838
rect 1964 502 2022 514
rect 2454 514 2466 826
rect 2500 514 2512 826
rect 2454 502 2512 514
rect 2542 826 2600 838
rect 2542 514 2554 826
rect 2588 514 2600 826
rect 2658 552 2670 864
rect 2704 552 2716 864
rect 2658 540 2716 552
rect 2746 864 2804 876
rect 2746 552 2758 864
rect 2792 552 2804 864
rect 3236 864 3294 876
rect 2746 540 2804 552
rect 3032 826 3090 838
rect 2542 502 2600 514
rect 3032 514 3044 826
rect 3078 514 3090 826
rect 3032 502 3090 514
rect 3120 826 3178 838
rect 3120 514 3132 826
rect 3166 514 3178 826
rect 3236 552 3248 864
rect 3282 552 3294 864
rect 3236 540 3294 552
rect 3324 864 3382 876
rect 3324 552 3336 864
rect 3370 552 3382 864
rect 3818 868 3876 880
rect 3324 540 3382 552
rect 3614 830 3672 842
rect 3120 502 3178 514
rect 3614 518 3626 830
rect 3660 518 3672 830
rect 3614 506 3672 518
rect 3702 830 3760 842
rect 3702 518 3714 830
rect 3748 518 3760 830
rect 3818 556 3830 868
rect 3864 556 3876 868
rect 3818 544 3876 556
rect 3906 868 3964 880
rect 3906 556 3918 868
rect 3952 556 3964 868
rect 4394 864 4452 876
rect 3906 544 3964 556
rect 4190 826 4248 838
rect 3702 506 3760 518
rect 4190 514 4202 826
rect 4236 514 4248 826
rect 4190 502 4248 514
rect 4278 826 4336 838
rect 4278 514 4290 826
rect 4324 514 4336 826
rect 4394 552 4406 864
rect 4440 552 4452 864
rect 4394 540 4452 552
rect 4482 864 4540 876
rect 4482 552 4494 864
rect 4528 552 4540 864
rect 4964 860 5022 872
rect 4482 540 4540 552
rect 4760 822 4818 834
rect 4278 502 4336 514
rect 4760 510 4772 822
rect 4806 510 4818 822
rect 4760 498 4818 510
rect 4848 822 4906 834
rect 4848 510 4860 822
rect 4894 510 4906 822
rect 4964 548 4976 860
rect 5010 548 5022 860
rect 4964 536 5022 548
rect 5052 860 5110 872
rect 5052 548 5064 860
rect 5098 548 5110 860
rect 5052 536 5110 548
rect 4848 498 4906 510
rect 1706 -1202 1764 -1190
rect 1506 -1240 1564 -1228
rect 1506 -1552 1518 -1240
rect 1552 -1552 1564 -1240
rect 1506 -1564 1564 -1552
rect 1594 -1240 1652 -1228
rect 1594 -1552 1606 -1240
rect 1640 -1552 1652 -1240
rect 1706 -1514 1718 -1202
rect 1752 -1514 1764 -1202
rect 1706 -1526 1764 -1514
rect 1794 -1202 1852 -1190
rect 1794 -1514 1806 -1202
rect 1840 -1514 1852 -1202
rect 1794 -1526 1852 -1514
rect 1908 -1242 1966 -1230
rect 1594 -1564 1652 -1552
rect 1908 -1554 1920 -1242
rect 1954 -1554 1966 -1242
rect 1908 -1566 1966 -1554
rect 1996 -1242 2054 -1230
rect 1996 -1554 2008 -1242
rect 2042 -1554 2054 -1242
rect 1996 -1566 2054 -1554
rect 1706 -1708 1764 -1696
rect 1506 -1746 1564 -1734
rect 1506 -2058 1518 -1746
rect 1552 -2058 1564 -1746
rect 1506 -2070 1564 -2058
rect 1594 -1746 1652 -1734
rect 1594 -2058 1606 -1746
rect 1640 -2058 1652 -1746
rect 1706 -2020 1718 -1708
rect 1752 -2020 1764 -1708
rect 1706 -2032 1764 -2020
rect 1794 -1708 1852 -1696
rect 1794 -2020 1806 -1708
rect 1840 -2020 1852 -1708
rect 1794 -2032 1852 -2020
rect 1906 -1746 1964 -1734
rect 1594 -2070 1652 -2058
rect 1906 -2058 1918 -1746
rect 1952 -2058 1964 -1746
rect 1906 -2070 1964 -2058
rect 1994 -1746 2052 -1734
rect 1994 -2058 2006 -1746
rect 2040 -2058 2052 -1746
rect 1994 -2070 2052 -2058
rect 1706 -2216 1764 -2204
rect 1506 -2254 1564 -2242
rect 1506 -2566 1518 -2254
rect 1552 -2566 1564 -2254
rect 1506 -2578 1564 -2566
rect 1594 -2254 1652 -2242
rect 1594 -2566 1606 -2254
rect 1640 -2566 1652 -2254
rect 1706 -2528 1718 -2216
rect 1752 -2528 1764 -2216
rect 1706 -2540 1764 -2528
rect 1794 -2216 1852 -2204
rect 1794 -2528 1806 -2216
rect 1840 -2528 1852 -2216
rect 1794 -2540 1852 -2528
rect 1906 -2254 1964 -2242
rect 1594 -2578 1652 -2566
rect 1906 -2566 1918 -2254
rect 1952 -2566 1964 -2254
rect 1906 -2578 1964 -2566
rect 1994 -2254 2052 -2242
rect 1994 -2566 2006 -2254
rect 2040 -2566 2052 -2254
rect 1994 -2578 2052 -2566
<< ndiffc >>
rect 124 92 158 216
rect 220 92 254 216
rect 316 92 350 216
rect 736 100 770 224
rect 832 100 866 224
rect 928 100 962 224
rect 1314 96 1348 220
rect 1410 96 1444 220
rect 1506 96 1540 220
rect 1888 104 1922 228
rect 1984 104 2018 228
rect 2080 104 2114 228
rect 2466 104 2500 228
rect 2562 104 2596 228
rect 2658 104 2692 228
rect 3044 104 3078 228
rect 3140 104 3174 228
rect 3236 104 3270 228
rect 3626 108 3660 232
rect 3722 108 3756 232
rect 3818 108 3852 232
rect 4202 104 4236 228
rect 4298 104 4332 228
rect 4394 104 4428 228
rect 4772 100 4806 224
rect 4868 100 4902 224
rect 4964 100 4998 224
rect 2182 -2246 2216 -1622
rect 2278 -2246 2312 -1622
rect 2374 -2246 2408 -1622
rect 2470 -2246 2504 -1622
rect 2566 -2246 2600 -1622
rect 2662 -2246 2696 -1622
rect 2758 -2246 2792 -1622
rect 2854 -2246 2888 -1622
rect 2950 -2246 2984 -1622
rect 3046 -2246 3080 -1622
<< pdiffc >>
rect 124 502 158 814
rect 212 502 246 814
rect 328 540 362 852
rect 416 540 450 852
rect 736 510 770 822
rect 824 510 858 822
rect 940 548 974 860
rect 1028 548 1062 860
rect 1314 506 1348 818
rect 1402 506 1436 818
rect 1518 544 1552 856
rect 1606 544 1640 856
rect 1888 514 1922 826
rect 1976 514 2010 826
rect 2092 552 2126 864
rect 2180 552 2214 864
rect 2466 514 2500 826
rect 2554 514 2588 826
rect 2670 552 2704 864
rect 2758 552 2792 864
rect 3044 514 3078 826
rect 3132 514 3166 826
rect 3248 552 3282 864
rect 3336 552 3370 864
rect 3626 518 3660 830
rect 3714 518 3748 830
rect 3830 556 3864 868
rect 3918 556 3952 868
rect 4202 514 4236 826
rect 4290 514 4324 826
rect 4406 552 4440 864
rect 4494 552 4528 864
rect 4772 510 4806 822
rect 4860 510 4894 822
rect 4976 548 5010 860
rect 5064 548 5098 860
rect 1518 -1552 1552 -1240
rect 1606 -1552 1640 -1240
rect 1718 -1514 1752 -1202
rect 1806 -1514 1840 -1202
rect 1920 -1554 1954 -1242
rect 2008 -1554 2042 -1242
rect 1518 -2058 1552 -1746
rect 1606 -2058 1640 -1746
rect 1718 -2020 1752 -1708
rect 1806 -2020 1840 -1708
rect 1918 -2058 1952 -1746
rect 2006 -2058 2040 -1746
rect 1518 -2566 1552 -2254
rect 1606 -2566 1640 -2254
rect 1718 -2528 1752 -2216
rect 1806 -2528 1840 -2216
rect 1918 -2566 1952 -2254
rect 2006 -2566 2040 -2254
<< psubdiff >>
rect -658 372 -344 416
rect -658 202 -586 372
rect -410 202 -344 372
rect 5198 360 5512 404
rect -658 152 -344 202
rect -658 -96 -346 152
rect 5198 190 5358 360
rect 5442 190 5512 360
rect 5198 152 5512 190
rect 5194 150 5512 152
rect 5602 226 6214 294
rect 5194 -96 5514 150
rect -658 -114 5514 -96
rect -658 -140 5512 -114
rect -658 -310 -594 -140
rect -418 -310 -134 -140
rect 42 -310 466 -140
rect 642 -310 1066 -140
rect 1242 -310 1666 -140
rect 1842 -310 2266 -140
rect 2442 -310 2866 -140
rect 3042 -310 3466 -140
rect 3642 -310 4066 -140
rect 4242 -310 4666 -140
rect 4842 -310 5266 -140
rect 5442 -310 5512 -140
rect 5602 -234 5662 226
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
rect -658 -314 5512 -310
rect -658 -360 1710 -314
rect 2174 -360 5512 -314
rect 2180 -966 3402 -914
rect 2180 -968 2568 -966
rect 2180 -970 2344 -968
rect 2268 -1118 2344 -970
rect 2494 -1116 2568 -968
rect 2718 -1116 2784 -966
rect 2934 -968 3184 -966
rect 2934 -1116 2976 -968
rect 2494 -1118 2976 -1116
rect 3126 -1116 3184 -968
rect 3334 -1116 3402 -966
rect 3126 -1118 3402 -1116
rect 2268 -1120 3402 -1118
rect 2180 -1162 3402 -1120
rect 2222 -1164 2252 -1162
rect 3148 -1190 3398 -1162
rect 3148 -1340 3194 -1190
rect 3344 -1340 3398 -1190
rect 3148 -1382 3398 -1340
rect 3148 -1532 3200 -1382
rect 3350 -1532 3398 -1382
rect 3148 -1576 3398 -1532
rect 3148 -1686 3204 -1576
rect 3150 -1726 3204 -1686
rect 3354 -1726 3398 -1576
rect 3150 -1762 3398 -1726
rect 3150 -1912 3206 -1762
rect 3356 -1912 3398 -1762
rect 3150 -1948 3398 -1912
rect 3150 -2068 3212 -1948
rect 3148 -2098 3212 -2068
rect 3362 -2098 3398 -1948
rect 3148 -2156 3398 -2098
rect 3148 -2306 3208 -2156
rect 3358 -2304 3398 -2156
rect 3358 -2306 3400 -2304
rect 3148 -2362 3400 -2306
rect 3148 -2392 3398 -2362
rect 3148 -2426 3202 -2392
rect 3106 -2430 3202 -2426
rect 3046 -2432 3202 -2430
rect 2118 -2468 3202 -2432
rect 2118 -2616 2150 -2468
rect 2300 -2470 3202 -2468
rect 2300 -2616 2362 -2470
rect 2118 -2620 2362 -2616
rect 2512 -2476 3202 -2470
rect 2512 -2620 2570 -2476
rect 2118 -2626 2570 -2620
rect 2720 -2478 3202 -2476
rect 2720 -2480 2990 -2478
rect 2720 -2626 2778 -2480
rect 2118 -2630 2778 -2626
rect 2928 -2628 2990 -2480
rect 3140 -2542 3202 -2478
rect 3352 -2436 3398 -2392
rect 3352 -2542 3400 -2436
rect 3140 -2628 3400 -2542
rect 2928 -2630 3400 -2628
rect 2118 -2650 3400 -2630
rect 2118 -2660 3398 -2650
rect 2146 -2664 3398 -2660
rect 3044 -2672 3398 -2664
<< nsubdiff >>
rect 2436 1718 2636 1720
rect 2436 1716 3702 1718
rect 3962 1716 5946 1718
rect 640 1714 5946 1716
rect -650 1594 5946 1714
rect -650 1570 5480 1594
rect -650 1324 226 1570
rect 474 1324 1226 1570
rect 1474 1324 2226 1570
rect 2474 1324 3226 1570
rect 3474 1324 4226 1570
rect 4474 1346 5480 1570
rect 5722 1346 5946 1594
rect 4474 1324 5946 1346
rect -650 1158 5946 1324
rect -650 1156 4746 1158
rect 5166 1156 5946 1158
rect -650 1152 112 1156
rect 636 1154 1124 1156
rect 1650 1154 3480 1156
rect 5170 1078 5946 1156
rect 5170 924 5952 1078
rect 5170 680 5450 924
rect 5698 680 5952 924
rect 5170 520 5952 680
rect 1132 -830 1400 -828
rect 2060 -830 2110 -824
rect 1132 -850 2110 -830
rect 1132 -852 1660 -850
rect 1132 -1046 1164 -852
rect 1130 -1050 1164 -1046
rect 1364 -1050 1420 -852
rect 1130 -1052 1420 -1050
rect 1620 -1050 1660 -852
rect 1860 -852 2110 -850
rect 1860 -1050 1894 -852
rect 1620 -1052 1894 -1050
rect 2068 -1052 2110 -852
rect 1130 -1074 2110 -1052
rect 1130 -1076 1648 -1074
rect 2060 -1076 2110 -1074
rect 1130 -1094 1386 -1076
rect 1132 -1104 1386 -1094
rect 1134 -1124 1386 -1104
rect 1134 -1136 1164 -1124
rect 1140 -1324 1164 -1136
rect 1364 -1146 1386 -1124
rect 1364 -1324 1384 -1146
rect 1140 -1358 1384 -1324
rect 1140 -1558 1164 -1358
rect 1364 -1558 1384 -1358
rect 1140 -1598 1384 -1558
rect 1140 -1798 1164 -1598
rect 1364 -1798 1384 -1598
rect 1140 -1836 1384 -1798
rect 1140 -2028 1162 -1836
rect 1362 -2028 1384 -1836
rect 1140 -2068 1384 -2028
rect 1140 -2268 1164 -2068
rect 1364 -2268 1384 -2068
rect 1140 -2304 1384 -2268
rect 1140 -2484 1162 -2304
rect 1130 -2504 1162 -2484
rect 1362 -2438 1384 -2304
rect 1362 -2504 1386 -2438
rect 1130 -2688 1386 -2504
rect 2004 -2688 2042 -2686
rect 1130 -2716 2048 -2688
rect 1130 -2728 1280 -2716
rect 1140 -2916 1280 -2728
rect 1480 -2718 2048 -2716
rect 1480 -2916 1586 -2718
rect 1140 -2918 1586 -2916
rect 1786 -2918 1866 -2718
rect 2028 -2918 2048 -2718
rect 1140 -2940 2048 -2918
rect 2000 -2942 2048 -2940
<< psubdiffcont >>
rect -586 202 -410 372
rect 5358 190 5442 360
rect -594 -310 -418 -140
rect -134 -310 42 -140
rect 466 -310 642 -140
rect 1066 -310 1242 -140
rect 1666 -310 1842 -140
rect 2266 -310 2442 -140
rect 2866 -310 3042 -140
rect 3466 -310 3642 -140
rect 4066 -310 4242 -140
rect 4666 -310 4842 -140
rect 5266 -310 5442 -140
rect 5662 -234 6142 226
rect 2180 -1120 2268 -970
rect 2344 -1118 2494 -968
rect 2568 -1116 2718 -966
rect 2784 -1116 2934 -966
rect 2976 -1118 3126 -968
rect 3184 -1116 3334 -966
rect 3194 -1340 3344 -1190
rect 3200 -1532 3350 -1382
rect 3204 -1726 3354 -1576
rect 3206 -1912 3356 -1762
rect 3212 -2098 3362 -1948
rect 3208 -2306 3358 -2156
rect 2150 -2616 2300 -2468
rect 2362 -2620 2512 -2470
rect 2570 -2626 2720 -2476
rect 2778 -2630 2928 -2480
rect 2990 -2628 3140 -2478
rect 3202 -2542 3352 -2392
<< nsubdiffcont >>
rect 226 1324 474 1570
rect 1226 1324 1474 1570
rect 2226 1324 2474 1570
rect 3226 1324 3474 1570
rect 4226 1324 4474 1570
rect 5480 1346 5722 1594
rect 5450 680 5698 924
rect 1164 -1050 1364 -852
rect 1420 -1052 1620 -852
rect 1660 -1050 1860 -850
rect 1894 -1052 2068 -852
rect 1164 -1324 1364 -1124
rect 1164 -1558 1364 -1358
rect 1164 -1798 1364 -1598
rect 1162 -2028 1362 -1836
rect 1164 -2268 1364 -2068
rect 1162 -2504 1362 -2304
rect 1280 -2916 1480 -2716
rect 1586 -2918 1786 -2718
rect 1866 -2918 2028 -2718
<< poly >>
rect 152 907 218 923
rect 152 873 168 907
rect 202 873 218 907
rect 764 915 830 931
rect 152 857 218 873
rect 374 864 404 890
rect 764 881 780 915
rect 814 881 830 915
rect 1342 911 1408 927
rect 764 865 830 881
rect 986 872 1016 898
rect 1342 877 1358 911
rect 1392 877 1408 911
rect 1916 919 1982 935
rect 170 826 200 857
rect 782 834 812 865
rect 374 497 404 528
rect 1342 861 1408 877
rect 1564 868 1594 894
rect 1916 885 1932 919
rect 1966 885 1982 919
rect 2494 919 2560 935
rect 1916 869 1982 885
rect 2138 876 2168 902
rect 2494 885 2510 919
rect 2544 885 2560 919
rect 3072 919 3138 935
rect 1360 830 1390 861
rect 986 505 1016 536
rect 170 464 200 490
rect 356 481 422 497
rect 356 447 372 481
rect 406 447 422 481
rect 782 472 812 498
rect 968 489 1034 505
rect 1934 838 1964 869
rect 1564 501 1594 532
rect 2494 869 2560 885
rect 2716 876 2746 902
rect 3072 885 3088 919
rect 3122 885 3138 919
rect 3654 923 3720 939
rect 2512 838 2542 869
rect 2138 509 2168 540
rect 356 431 422 447
rect 968 455 984 489
rect 1018 455 1034 489
rect 1360 468 1390 494
rect 1546 485 1612 501
rect 968 439 1034 455
rect 1546 451 1562 485
rect 1596 451 1612 485
rect 1934 476 1964 502
rect 2120 493 2186 509
rect 3072 869 3138 885
rect 3294 876 3324 902
rect 3654 889 3670 923
rect 3704 889 3720 923
rect 4230 919 4296 935
rect 3090 838 3120 869
rect 2716 509 2746 540
rect 1546 435 1612 451
rect 2120 459 2136 493
rect 2170 459 2186 493
rect 2512 476 2542 502
rect 2698 493 2764 509
rect 3654 873 3720 889
rect 3876 880 3906 906
rect 4230 885 4246 919
rect 4280 885 4296 919
rect 4800 915 4866 931
rect 3672 842 3702 873
rect 3294 509 3324 540
rect 2120 443 2186 459
rect 2698 459 2714 493
rect 2748 459 2764 493
rect 3090 476 3120 502
rect 3276 493 3342 509
rect 4230 869 4296 885
rect 4452 876 4482 902
rect 4800 881 4816 915
rect 4850 881 4866 915
rect 4248 838 4278 869
rect 3876 513 3906 544
rect 2698 443 2764 459
rect 3276 459 3292 493
rect 3326 459 3342 493
rect 3672 480 3702 506
rect 3858 497 3924 513
rect 4800 865 4866 881
rect 5022 872 5052 898
rect 4818 834 4848 865
rect 4452 509 4482 540
rect 3276 443 3342 459
rect 3858 463 3874 497
rect 3908 463 3924 497
rect 4248 476 4278 502
rect 4434 493 4500 509
rect 5022 505 5052 536
rect 3858 447 3924 463
rect 4434 459 4450 493
rect 4484 459 4500 493
rect 4818 472 4848 498
rect 5004 489 5070 505
rect 4434 443 4500 459
rect 5004 455 5020 489
rect 5054 455 5070 489
rect 5004 439 5070 455
rect 252 300 318 316
rect 252 266 268 300
rect 302 266 318 300
rect 174 228 204 254
rect 252 250 318 266
rect 864 308 930 324
rect 864 274 880 308
rect 914 274 930 308
rect 270 228 300 250
rect 786 236 816 262
rect 864 258 930 274
rect 1442 304 1508 320
rect 1442 270 1458 304
rect 1492 270 1508 304
rect 882 236 912 258
rect 1364 232 1394 258
rect 1442 254 1508 270
rect 2016 312 2082 328
rect 2016 278 2032 312
rect 2066 278 2082 312
rect 1460 232 1490 254
rect 1938 240 1968 266
rect 2016 262 2082 278
rect 2594 312 2660 328
rect 2594 278 2610 312
rect 2644 278 2660 312
rect 2034 240 2064 262
rect 2516 240 2546 266
rect 2594 262 2660 278
rect 3172 312 3238 328
rect 3172 278 3188 312
rect 3222 278 3238 312
rect 2612 240 2642 262
rect 3094 240 3124 266
rect 3172 262 3238 278
rect 3754 316 3820 332
rect 3754 282 3770 316
rect 3804 282 3820 316
rect 3190 240 3220 262
rect 3676 244 3706 270
rect 3754 266 3820 282
rect 4330 312 4396 328
rect 4330 278 4346 312
rect 4380 278 4396 312
rect 3772 244 3802 266
rect 174 58 204 80
rect 156 42 222 58
rect 270 54 300 80
rect 786 66 816 88
rect 156 8 172 42
rect 206 8 222 42
rect 156 -8 222 8
rect 768 50 834 66
rect 882 62 912 88
rect 4252 240 4282 266
rect 4330 262 4396 278
rect 4900 308 4966 324
rect 4900 274 4916 308
rect 4950 274 4966 308
rect 4348 240 4378 262
rect 1364 62 1394 84
rect 768 16 784 50
rect 818 16 834 50
rect 768 0 834 16
rect 1346 46 1412 62
rect 1460 58 1490 84
rect 1938 70 1968 92
rect 1346 12 1362 46
rect 1396 12 1412 46
rect 1346 -4 1412 12
rect 1920 54 1986 70
rect 2034 66 2064 92
rect 2516 70 2546 92
rect 1920 20 1936 54
rect 1970 20 1986 54
rect 1920 4 1986 20
rect 2498 54 2564 70
rect 2612 66 2642 92
rect 3094 70 3124 92
rect 2498 20 2514 54
rect 2548 20 2564 54
rect 2498 4 2564 20
rect 3076 54 3142 70
rect 3190 66 3220 92
rect 3676 74 3706 96
rect 3076 20 3092 54
rect 3126 20 3142 54
rect 3076 4 3142 20
rect 3658 58 3724 74
rect 3772 70 3802 96
rect 4822 236 4852 262
rect 4900 258 4966 274
rect 4918 236 4948 258
rect 4252 70 4282 92
rect 3658 24 3674 58
rect 3708 24 3724 58
rect 3658 8 3724 24
rect 4234 54 4300 70
rect 4348 66 4378 92
rect 4822 66 4852 88
rect 4234 20 4250 54
rect 4284 20 4300 54
rect 4234 4 4300 20
rect 4804 50 4870 66
rect 4918 62 4948 88
rect 4804 16 4820 50
rect 4854 16 4870 50
rect 4804 0 4870 16
rect 1546 -1147 1612 -1131
rect 1546 -1181 1562 -1147
rect 1596 -1181 1612 -1147
rect 1948 -1149 2014 -1133
rect 1546 -1197 1612 -1181
rect 1764 -1190 1794 -1164
rect 1948 -1183 1964 -1149
rect 1998 -1183 2014 -1149
rect 1564 -1228 1594 -1197
rect 1948 -1199 2014 -1183
rect 1966 -1230 1996 -1199
rect 1764 -1557 1794 -1526
rect 1564 -1590 1594 -1564
rect 1746 -1573 1812 -1557
rect 2310 -1538 2376 -1522
rect 1746 -1607 1762 -1573
rect 1796 -1607 1812 -1573
rect 1966 -1592 1996 -1566
rect 2310 -1572 2326 -1538
rect 2360 -1572 2376 -1538
rect 1746 -1623 1812 -1607
rect 2232 -1610 2262 -1584
rect 2310 -1588 2376 -1572
rect 2502 -1538 2568 -1522
rect 2502 -1572 2518 -1538
rect 2552 -1572 2568 -1538
rect 2328 -1610 2358 -1588
rect 2424 -1610 2454 -1584
rect 2502 -1588 2568 -1572
rect 2694 -1538 2760 -1522
rect 2694 -1572 2710 -1538
rect 2744 -1572 2760 -1538
rect 2520 -1610 2550 -1588
rect 2616 -1610 2646 -1584
rect 2694 -1588 2760 -1572
rect 2886 -1538 2952 -1522
rect 2886 -1572 2902 -1538
rect 2936 -1572 2952 -1538
rect 2712 -1610 2742 -1588
rect 2808 -1610 2838 -1584
rect 2886 -1588 2952 -1572
rect 2904 -1610 2934 -1588
rect 3000 -1610 3030 -1584
rect 1546 -1653 1612 -1637
rect 1546 -1687 1562 -1653
rect 1596 -1687 1612 -1653
rect 1946 -1653 2012 -1637
rect 1546 -1703 1612 -1687
rect 1764 -1696 1794 -1670
rect 1946 -1687 1962 -1653
rect 1996 -1687 2012 -1653
rect 1564 -1734 1594 -1703
rect 1946 -1703 2012 -1687
rect 1964 -1734 1994 -1703
rect 1764 -2063 1794 -2032
rect 1564 -2096 1594 -2070
rect 1746 -2079 1812 -2063
rect 1746 -2113 1762 -2079
rect 1796 -2113 1812 -2079
rect 1964 -2096 1994 -2070
rect 1746 -2129 1812 -2113
rect 1546 -2161 1612 -2145
rect 1546 -2195 1562 -2161
rect 1596 -2195 1612 -2161
rect 1946 -2161 2012 -2145
rect 1546 -2211 1612 -2195
rect 1764 -2204 1794 -2178
rect 1946 -2195 1962 -2161
rect 1996 -2195 2012 -2161
rect 1564 -2242 1594 -2211
rect 1946 -2211 2012 -2195
rect 1964 -2242 1994 -2211
rect 1764 -2571 1794 -2540
rect 1564 -2604 1594 -2578
rect 1746 -2587 1812 -2571
rect 2232 -2280 2262 -2258
rect 2214 -2296 2280 -2280
rect 2328 -2284 2358 -2258
rect 2424 -2280 2454 -2258
rect 2214 -2330 2230 -2296
rect 2264 -2330 2280 -2296
rect 2214 -2346 2280 -2330
rect 2406 -2296 2472 -2280
rect 2520 -2284 2550 -2258
rect 2616 -2280 2646 -2258
rect 2406 -2330 2422 -2296
rect 2456 -2330 2472 -2296
rect 2406 -2346 2472 -2330
rect 2598 -2296 2664 -2280
rect 2712 -2284 2742 -2258
rect 2808 -2280 2838 -2258
rect 2598 -2330 2614 -2296
rect 2648 -2330 2664 -2296
rect 2598 -2346 2664 -2330
rect 2790 -2296 2856 -2280
rect 2904 -2284 2934 -2258
rect 3000 -2280 3030 -2258
rect 2790 -2330 2806 -2296
rect 2840 -2330 2856 -2296
rect 2790 -2346 2856 -2330
rect 2982 -2296 3048 -2280
rect 2982 -2330 2998 -2296
rect 3032 -2330 3048 -2296
rect 2982 -2346 3048 -2330
rect 1746 -2621 1762 -2587
rect 1796 -2621 1812 -2587
rect 1964 -2604 1994 -2578
rect 1746 -2637 1812 -2621
<< polycont >>
rect 168 873 202 907
rect 780 881 814 915
rect 1358 877 1392 911
rect 1932 885 1966 919
rect 2510 885 2544 919
rect 372 447 406 481
rect 3088 885 3122 919
rect 984 455 1018 489
rect 1562 451 1596 485
rect 3670 889 3704 923
rect 2136 459 2170 493
rect 4246 885 4280 919
rect 2714 459 2748 493
rect 4816 881 4850 915
rect 3292 459 3326 493
rect 3874 463 3908 497
rect 4450 459 4484 493
rect 5020 455 5054 489
rect 268 266 302 300
rect 880 274 914 308
rect 1458 270 1492 304
rect 2032 278 2066 312
rect 2610 278 2644 312
rect 3188 278 3222 312
rect 3770 282 3804 316
rect 4346 278 4380 312
rect 172 8 206 42
rect 4916 274 4950 308
rect 784 16 818 50
rect 1362 12 1396 46
rect 1936 20 1970 54
rect 2514 20 2548 54
rect 3092 20 3126 54
rect 3674 24 3708 58
rect 4250 20 4284 54
rect 4820 16 4854 50
rect 1562 -1181 1596 -1147
rect 1964 -1183 1998 -1149
rect 1762 -1607 1796 -1573
rect 2326 -1572 2360 -1538
rect 2518 -1572 2552 -1538
rect 2710 -1572 2744 -1538
rect 2902 -1572 2936 -1538
rect 1562 -1687 1596 -1653
rect 1962 -1687 1996 -1653
rect 1762 -2113 1796 -2079
rect 1562 -2195 1596 -2161
rect 1962 -2195 1996 -2161
rect 2230 -2330 2264 -2296
rect 2422 -2330 2456 -2296
rect 2614 -2330 2648 -2296
rect 2806 -2330 2840 -2296
rect 2998 -2330 3032 -2296
rect 1762 -2621 1796 -2587
<< locali >>
rect -650 1658 -170 1696
rect -650 1600 -624 1658
rect -892 1590 -624 1600
rect -908 1316 -624 1590
rect -908 -638 -712 1316
rect -650 1266 -624 1316
rect -224 1600 -170 1658
rect -224 1592 192 1600
rect 5676 1596 5722 1598
rect 5484 1594 5736 1596
rect 4838 1592 5480 1594
rect -224 1570 5480 1592
rect -224 1324 226 1570
rect 474 1324 1226 1570
rect 1474 1324 2226 1570
rect 2474 1324 3226 1570
rect 3474 1324 4226 1570
rect 4474 1346 5480 1570
rect 5722 1346 5742 1594
rect 4474 1324 5742 1346
rect -224 1320 5742 1324
rect -224 1316 -146 1320
rect 4838 1316 5742 1320
rect -224 1266 -170 1316
rect 5224 1314 5742 1316
rect -650 1236 -170 1266
rect -556 1224 -240 1236
rect 5444 1078 5742 1314
rect 5438 1070 5742 1078
rect 5438 924 5734 1070
rect 3520 923 3720 924
rect 1782 919 1982 920
rect 630 915 830 916
rect 18 907 218 908
rect 18 874 168 907
rect -600 376 -506 378
rect -602 372 -394 376
rect -602 202 -586 372
rect -410 202 -394 372
rect 18 320 54 874
rect 152 873 168 874
rect 202 873 218 907
rect 630 882 780 915
rect 328 852 362 868
rect 124 814 158 830
rect 124 486 158 502
rect 212 814 246 830
rect 328 524 362 540
rect 416 854 450 868
rect 416 524 450 540
rect 212 486 246 502
rect 384 481 418 482
rect 356 447 372 481
rect 406 447 422 481
rect -22 302 54 320
rect 384 390 420 447
rect 630 390 666 882
rect 764 881 780 882
rect 814 881 830 915
rect 1208 911 1408 912
rect 1208 878 1358 911
rect 940 860 974 876
rect 736 822 770 838
rect 736 494 770 510
rect 824 822 858 838
rect 940 532 974 548
rect 1028 862 1062 876
rect 1028 532 1062 548
rect 824 494 858 510
rect 996 489 1030 490
rect 968 455 984 489
rect 1018 455 1034 489
rect 384 338 666 390
rect -22 300 314 302
rect -602 -140 -394 202
rect -84 284 268 300
rect -84 210 -72 284
rect 18 268 268 284
rect 18 266 50 268
rect 252 266 268 268
rect 302 266 318 300
rect 18 210 34 266
rect -84 196 34 210
rect 124 216 158 232
rect 220 216 254 232
rect 204 124 220 170
rect 124 76 158 92
rect 316 216 350 232
rect 254 124 270 170
rect 220 76 254 92
rect 316 76 350 92
rect 156 8 172 42
rect 206 8 222 42
rect 166 -12 222 8
rect 384 -12 420 338
rect 630 310 666 338
rect 996 370 1032 455
rect 1208 370 1244 878
rect 1342 877 1358 878
rect 1392 877 1408 911
rect 1782 886 1932 919
rect 1518 856 1552 872
rect 1406 834 1448 836
rect 1314 818 1348 834
rect 1314 490 1348 506
rect 1402 818 1448 834
rect 1436 528 1448 818
rect 1518 528 1552 544
rect 1606 858 1640 872
rect 1606 528 1640 544
rect 1402 490 1436 506
rect 1574 485 1608 486
rect 1546 451 1562 485
rect 1596 451 1612 485
rect 996 336 1244 370
rect 630 308 926 310
rect 630 276 880 308
rect 864 274 880 276
rect 914 274 930 308
rect 736 224 770 240
rect 724 100 736 152
rect 832 224 866 240
rect 770 100 786 152
rect 820 100 832 152
rect 928 224 962 240
rect 866 100 878 152
rect 724 94 786 100
rect 736 84 770 94
rect 832 84 866 100
rect 928 84 962 100
rect 768 16 784 50
rect 818 16 834 50
rect 166 -46 420 -12
rect 778 -4 834 16
rect 996 -4 1032 336
rect 1208 306 1244 336
rect 1574 378 1610 451
rect 1782 378 1818 886
rect 1916 885 1932 886
rect 1966 885 1982 919
rect 2360 919 2560 920
rect 2360 886 2510 919
rect 2092 864 2126 880
rect 1980 842 2022 844
rect 1888 826 1922 842
rect 1888 498 1922 514
rect 1976 826 2022 842
rect 2010 528 2022 826
rect 2092 536 2126 552
rect 2180 866 2214 880
rect 2180 536 2214 552
rect 1976 498 2010 514
rect 2148 493 2182 494
rect 2120 459 2136 493
rect 2170 459 2186 493
rect 1574 342 1818 378
rect 1208 304 1504 306
rect 1208 272 1458 304
rect 1442 270 1458 272
rect 1492 270 1508 304
rect 1314 220 1348 236
rect 1410 220 1444 236
rect 1394 120 1410 158
rect 1314 80 1348 96
rect 1506 220 1540 236
rect 1444 120 1458 158
rect 1410 80 1444 96
rect 1506 80 1540 96
rect 1346 12 1362 46
rect 1396 12 1412 46
rect 778 -38 1032 -4
rect 1356 -8 1412 12
rect 1574 -8 1610 342
rect 1782 314 1818 342
rect 2148 384 2184 459
rect 2360 384 2396 886
rect 2494 885 2510 886
rect 2544 885 2560 919
rect 2938 919 3138 920
rect 2938 886 3088 919
rect 2670 864 2704 880
rect 2466 826 2500 842
rect 2466 498 2500 514
rect 2554 826 2588 842
rect 2670 536 2704 552
rect 2758 866 2792 880
rect 2758 536 2792 552
rect 2554 498 2588 514
rect 2726 493 2760 494
rect 2698 459 2714 493
rect 2748 459 2764 493
rect 2148 348 2396 384
rect 1782 312 2078 314
rect 1782 280 2032 312
rect 2016 278 2032 280
rect 2066 278 2082 312
rect 1888 228 1922 244
rect 1984 228 2018 244
rect 1968 126 1984 192
rect 1888 88 1922 104
rect 2080 228 2114 244
rect 2018 136 2036 192
rect 2018 126 2032 136
rect 1984 88 2018 104
rect 2080 88 2114 104
rect 1920 20 1936 54
rect 1970 20 1986 54
rect 1356 -42 1610 -8
rect 1930 0 1986 20
rect 2148 0 2184 348
rect 2360 314 2396 348
rect 2726 388 2762 459
rect 2938 388 2974 886
rect 3072 885 3088 886
rect 3122 885 3138 919
rect 3520 890 3670 923
rect 3248 864 3282 880
rect 3044 826 3078 842
rect 3044 498 3078 514
rect 3132 826 3166 842
rect 3248 536 3282 552
rect 3336 866 3370 880
rect 3336 536 3370 552
rect 3132 498 3166 514
rect 3304 493 3338 494
rect 3276 459 3292 493
rect 3326 459 3342 493
rect 2726 352 2974 388
rect 2360 312 2656 314
rect 2360 280 2610 312
rect 2594 278 2610 280
rect 2644 278 2660 312
rect 2466 228 2500 244
rect 2562 228 2596 244
rect 2548 128 2562 182
rect 2466 88 2500 104
rect 2658 228 2692 244
rect 2596 146 2614 182
rect 2596 128 2612 146
rect 2562 88 2596 104
rect 2658 88 2692 104
rect 2498 20 2514 54
rect 2548 20 2564 54
rect 1930 -34 2184 0
rect 2508 0 2564 20
rect 2726 0 2762 352
rect 2938 314 2974 352
rect 3304 394 3340 459
rect 3520 394 3556 890
rect 3654 889 3670 890
rect 3704 889 3720 923
rect 4096 919 4296 920
rect 4096 886 4246 919
rect 3830 868 3864 884
rect 3626 830 3660 846
rect 3626 502 3660 518
rect 3714 830 3748 846
rect 3830 540 3864 556
rect 3918 870 3952 884
rect 3918 540 3952 556
rect 3714 502 3748 518
rect 3886 497 3920 498
rect 3858 463 3874 497
rect 3908 463 3924 497
rect 3304 358 3556 394
rect 2938 312 3234 314
rect 2938 280 3188 312
rect 3172 278 3188 280
rect 3222 278 3238 312
rect 3044 228 3078 244
rect 3140 228 3174 244
rect 3124 126 3140 182
rect 3044 88 3078 104
rect 3236 228 3270 244
rect 3174 140 3192 182
rect 3174 126 3188 140
rect 3140 88 3174 104
rect 3236 88 3270 104
rect 3076 20 3092 54
rect 3126 20 3142 54
rect 2508 -34 2762 0
rect 3086 0 3142 20
rect 3304 0 3340 358
rect 3520 318 3556 358
rect 3886 394 3922 463
rect 4096 394 4132 886
rect 4230 885 4246 886
rect 4280 885 4296 919
rect 4666 915 4866 916
rect 4666 882 4816 915
rect 4406 864 4440 880
rect 4202 826 4236 842
rect 4202 498 4236 514
rect 4290 826 4324 842
rect 4406 536 4440 552
rect 4494 866 4528 880
rect 4494 536 4528 552
rect 4290 498 4324 514
rect 4462 493 4496 494
rect 4434 459 4450 493
rect 4484 459 4500 493
rect 3886 358 4134 394
rect 4462 384 4498 459
rect 4666 384 4702 882
rect 4800 881 4816 882
rect 4850 881 4866 915
rect 4976 860 5010 876
rect 4772 822 4806 838
rect 4772 494 4806 510
rect 4860 822 4894 838
rect 4976 532 5010 548
rect 5064 862 5098 876
rect 5438 704 5450 924
rect 5434 680 5450 704
rect 5698 680 5734 924
rect 5434 670 5734 680
rect 5434 666 5714 670
rect 5064 532 5098 548
rect 4860 494 4894 510
rect 5032 489 5066 490
rect 5004 455 5020 489
rect 5054 455 5070 489
rect 3520 316 3816 318
rect 3520 284 3770 316
rect 3754 282 3770 284
rect 3804 282 3820 316
rect 3626 232 3660 248
rect 3722 232 3756 248
rect 3706 134 3722 188
rect 3626 92 3660 108
rect 3818 232 3852 248
rect 3756 146 3772 188
rect 3756 134 3770 146
rect 3722 92 3756 108
rect 3818 92 3852 108
rect 3658 24 3674 58
rect 3708 24 3724 58
rect 3086 -34 3340 0
rect 3668 4 3724 24
rect 3886 4 3922 358
rect 4096 314 4132 358
rect 4462 348 4702 384
rect 4096 312 4392 314
rect 4096 280 4346 312
rect 4330 278 4346 280
rect 4380 278 4396 312
rect 4202 228 4236 244
rect 4298 228 4332 244
rect 4282 126 4298 178
rect 4202 88 4236 104
rect 4394 228 4428 244
rect 4332 126 4346 178
rect 4298 88 4332 104
rect 4394 88 4428 104
rect 4234 20 4250 54
rect 4284 20 4300 54
rect 3668 -30 3922 4
rect 4244 0 4300 20
rect 4462 0 4498 348
rect 4666 310 4702 348
rect 4666 308 4962 310
rect 4666 276 4916 308
rect 4900 274 4916 276
rect 4950 274 4966 308
rect 4772 224 4806 240
rect 4544 94 4634 110
rect 4544 32 4558 94
rect 4620 50 4634 94
rect 4868 224 4902 240
rect 4854 128 4868 180
rect 4772 84 4806 100
rect 4964 224 4998 240
rect 4902 128 4918 180
rect 4868 84 4902 100
rect 4964 84 4998 100
rect 4620 32 4820 50
rect 4544 18 4820 32
rect 4244 -34 4498 0
rect 4560 16 4820 18
rect 4854 16 4872 50
rect 4560 -2 4872 16
rect 4814 -4 4872 -2
rect 5032 -4 5068 455
rect 5334 364 5402 366
rect 5334 360 5446 364
rect 5334 190 5358 360
rect 5442 234 5458 360
rect 5442 190 5460 234
rect 5334 152 5460 190
rect 4814 -38 5068 -4
rect 5264 126 5460 152
rect 5602 226 6214 294
rect 5602 126 5662 226
rect 5264 -62 5662 126
rect 3640 -140 4066 -136
rect 5264 -140 5458 -62
rect -602 -310 -594 -140
rect -418 -310 -134 -140
rect 42 -310 466 -140
rect 642 -310 1066 -140
rect 1242 -310 1666 -140
rect 1842 -310 2266 -140
rect 2442 -310 2866 -140
rect 3042 -310 3466 -140
rect 3642 -310 4066 -140
rect 4242 -310 4666 -140
rect 4842 -310 5266 -140
rect 5442 -310 5458 -140
rect 5602 -234 5662 -62
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
rect -602 -312 5268 -310
rect -602 -314 4858 -312
rect -602 -322 1710 -314
rect 2174 -322 3360 -314
rect -602 -324 178 -322
rect -602 -326 -192 -324
rect -908 -912 -718 -638
rect 1400 -844 2094 -840
rect 1148 -850 2094 -844
rect 1148 -852 1660 -850
rect 1148 -894 1164 -852
rect -908 -918 456 -912
rect 1118 -914 1164 -894
rect 930 -918 1164 -914
rect -908 -1004 1164 -918
rect -906 -1050 1164 -1004
rect 1364 -1050 1420 -852
rect -906 -1052 1420 -1050
rect 1620 -1050 1660 -852
rect 1860 -852 2094 -850
rect 1860 -1050 1894 -852
rect 1620 -1052 1894 -1050
rect 2068 -1052 2094 -852
rect 3164 -938 3360 -322
rect 2180 -948 3360 -938
rect 2180 -966 3370 -948
rect 2180 -968 2568 -966
rect 2180 -970 2344 -968
rect -906 -1064 2094 -1052
rect -906 -1066 2068 -1064
rect -906 -1068 1640 -1066
rect -906 -1070 1386 -1068
rect -906 -1104 1382 -1070
rect 1134 -1124 1382 -1104
rect 1134 -1136 1164 -1124
rect 1150 -1324 1164 -1136
rect 1364 -1136 1382 -1124
rect 2176 -1120 2180 -1036
rect 2268 -1118 2344 -970
rect 2494 -1116 2568 -968
rect 2718 -1116 2784 -966
rect 2934 -968 3184 -966
rect 2934 -1116 2976 -968
rect 2494 -1118 2976 -1116
rect 3126 -1116 3184 -968
rect 3334 -1116 3370 -966
rect 3126 -1118 3370 -1116
rect 2268 -1120 3370 -1118
rect 1364 -1270 1380 -1136
rect 1544 -1140 1602 -1132
rect 1544 -1147 1622 -1140
rect 1544 -1181 1562 -1147
rect 1596 -1181 1622 -1147
rect 2176 -1142 3370 -1120
rect 1544 -1182 1622 -1181
rect 1948 -1149 1998 -1148
rect 1544 -1190 1602 -1182
rect 1948 -1183 1964 -1149
rect 1998 -1183 2014 -1149
rect 1718 -1202 1752 -1186
rect 1518 -1240 1552 -1224
rect 1364 -1324 1518 -1270
rect 1150 -1338 1518 -1324
rect 1150 -1358 1380 -1338
rect 1150 -1558 1164 -1358
rect 1364 -1558 1380 -1358
rect 1150 -1598 1380 -1558
rect 1606 -1240 1640 -1224
rect 1552 -1338 1558 -1270
rect 1518 -1568 1552 -1552
rect 1718 -1530 1752 -1514
rect 1806 -1202 1840 -1186
rect 1948 -1190 1998 -1183
rect 1806 -1530 1840 -1514
rect 1920 -1242 1954 -1226
rect 1606 -1568 1640 -1552
rect 1920 -1570 1954 -1554
rect 2008 -1242 2042 -1226
rect 2176 -1478 2224 -1142
rect 2008 -1570 2042 -1554
rect 1150 -1798 1164 -1598
rect 1364 -1798 1380 -1598
rect 1746 -1607 1762 -1573
rect 1796 -1574 1812 -1573
rect 1796 -1607 1818 -1574
rect 1752 -1616 1818 -1607
rect 2178 -1622 2224 -1478
rect 3176 -1190 3370 -1142
rect 3176 -1340 3194 -1190
rect 3344 -1340 3370 -1190
rect 3176 -1382 3370 -1340
rect 2300 -1538 2388 -1528
rect 2300 -1572 2326 -1538
rect 2360 -1572 2388 -1538
rect 2488 -1538 2576 -1528
rect 2488 -1572 2518 -1538
rect 2552 -1572 2576 -1538
rect 2680 -1538 2768 -1526
rect 2680 -1572 2710 -1538
rect 2744 -1572 2768 -1538
rect 2870 -1538 2958 -1526
rect 2870 -1572 2902 -1538
rect 2936 -1572 2958 -1538
rect 3176 -1532 3200 -1382
rect 3350 -1532 3370 -1382
rect 3176 -1576 3370 -1532
rect 2178 -1638 2182 -1622
rect 1546 -1653 1612 -1652
rect 1950 -1653 2016 -1652
rect 1546 -1687 1562 -1653
rect 1596 -1687 1612 -1653
rect 1946 -1687 1962 -1653
rect 1996 -1687 2016 -1653
rect 1546 -1694 1612 -1687
rect 1718 -1708 1752 -1692
rect 1150 -1836 1380 -1798
rect 1150 -2028 1162 -1836
rect 1362 -2028 1380 -1836
rect 1150 -2068 1380 -2028
rect 1150 -2268 1164 -2068
rect 1364 -2268 1380 -2068
rect 1518 -1746 1552 -1730
rect 1518 -2074 1552 -2058
rect 1606 -1746 1640 -1730
rect 1718 -2036 1752 -2020
rect 1806 -1708 1840 -1692
rect 1950 -1694 2016 -1687
rect 2180 -1692 2182 -1638
rect 1806 -2036 1840 -2020
rect 1918 -1746 1952 -1730
rect 1606 -2074 1640 -2058
rect 1918 -2074 1952 -2058
rect 2006 -1746 2040 -1730
rect 2168 -1844 2182 -1692
rect 2172 -2052 2182 -1844
rect 2006 -2074 2040 -2058
rect 1748 -2079 1814 -2078
rect 1746 -2113 1762 -2079
rect 1796 -2113 1814 -2079
rect 1748 -2120 1814 -2113
rect 1946 -2161 2012 -2156
rect 1546 -2162 1562 -2161
rect 1454 -2195 1562 -2162
rect 1596 -2162 1612 -2161
rect 1596 -2195 1614 -2162
rect 1454 -2198 1614 -2195
rect 1946 -2195 1962 -2161
rect 1996 -2195 2012 -2161
rect 1946 -2198 2012 -2195
rect 1718 -2216 1752 -2200
rect 1150 -2304 1380 -2268
rect 1150 -2438 1162 -2304
rect 1144 -2504 1162 -2438
rect 1362 -2438 1380 -2304
rect 1518 -2254 1552 -2238
rect 1362 -2504 1386 -2438
rect 1144 -2694 1386 -2504
rect 1518 -2582 1552 -2566
rect 1606 -2254 1640 -2238
rect 1718 -2544 1752 -2528
rect 1806 -2216 1840 -2200
rect 1806 -2544 1840 -2528
rect 1918 -2254 1952 -2238
rect 1606 -2582 1640 -2566
rect 1918 -2582 1952 -2566
rect 2006 -2254 2040 -2238
rect 2216 -1692 2224 -1622
rect 2278 -1622 2312 -1606
rect 2216 -2052 2228 -1692
rect 2266 -1878 2278 -1702
rect 2272 -1988 2278 -1878
rect 2182 -2262 2216 -2246
rect 2374 -1622 2408 -1606
rect 2312 -1988 2320 -1796
rect 2364 -1878 2374 -1702
rect 2370 -1986 2374 -1878
rect 2278 -2262 2312 -2246
rect 2470 -1622 2504 -1606
rect 2408 -1986 2418 -1794
rect 2460 -2046 2470 -1690
rect 2374 -2262 2408 -2246
rect 2566 -1622 2600 -1606
rect 2504 -2046 2516 -1836
rect 2556 -1848 2566 -1684
rect 2554 -2058 2566 -1848
rect 2470 -2262 2504 -2246
rect 2662 -1622 2696 -1606
rect 2600 -2058 2610 -1848
rect 2650 -2052 2662 -1696
rect 2566 -2262 2600 -2246
rect 2758 -1622 2792 -1606
rect 2750 -1842 2758 -1694
rect 2696 -2052 2706 -1842
rect 2746 -2052 2758 -1842
rect 2662 -2262 2696 -2246
rect 2854 -1622 2888 -1606
rect 2792 -1842 2794 -1694
rect 2792 -2052 2802 -1842
rect 2848 -1846 2854 -1700
rect 2842 -2056 2854 -1846
rect 2758 -2262 2792 -2246
rect 2950 -1622 2984 -1606
rect 2888 -1846 2892 -1700
rect 2940 -1836 2950 -1716
rect 2888 -2056 2898 -1846
rect 2936 -2046 2950 -1836
rect 2854 -2262 2888 -2246
rect 3046 -1622 3080 -1606
rect 2984 -2046 2992 -1836
rect 2950 -2262 2984 -2246
rect 3176 -1726 3204 -1576
rect 3354 -1726 3370 -1576
rect 3176 -1762 3370 -1726
rect 3176 -1912 3206 -1762
rect 3356 -1912 3370 -1762
rect 3176 -1928 3370 -1912
rect 3174 -1948 3370 -1928
rect 3174 -2006 3212 -1948
rect 3046 -2262 3080 -2246
rect 3176 -2098 3212 -2006
rect 3362 -2098 3370 -1948
rect 3176 -2156 3370 -2098
rect 2214 -2298 2230 -2296
rect 2212 -2330 2230 -2298
rect 2264 -2298 2280 -2296
rect 2264 -2330 2298 -2298
rect 2212 -2344 2298 -2330
rect 2390 -2330 2422 -2296
rect 2456 -2330 2478 -2296
rect 2598 -2298 2614 -2296
rect 2390 -2342 2478 -2330
rect 2586 -2330 2614 -2298
rect 2648 -2298 2664 -2296
rect 2648 -2330 2674 -2298
rect 2586 -2344 2674 -2330
rect 2778 -2330 2806 -2296
rect 2840 -2330 2866 -2296
rect 2778 -2342 2866 -2330
rect 2966 -2330 2998 -2296
rect 3032 -2330 3054 -2296
rect 3176 -2306 3208 -2156
rect 3358 -2306 3370 -2156
rect 3176 -2316 3370 -2306
rect 2966 -2342 3054 -2330
rect 3174 -2392 3370 -2316
rect 3174 -2446 3202 -2392
rect 2006 -2582 2040 -2566
rect 2132 -2468 3202 -2446
rect 1746 -2587 1816 -2586
rect 1746 -2621 1762 -2587
rect 1796 -2621 1816 -2587
rect 1746 -2634 1816 -2621
rect 2132 -2616 2150 -2468
rect 2300 -2470 3202 -2468
rect 2300 -2616 2362 -2470
rect 2132 -2620 2362 -2616
rect 2512 -2476 3202 -2470
rect 2512 -2620 2570 -2476
rect 2132 -2626 2570 -2620
rect 2720 -2478 3202 -2476
rect 2720 -2480 2990 -2478
rect 2720 -2626 2778 -2480
rect 2132 -2630 2778 -2626
rect 2928 -2628 2990 -2480
rect 3140 -2542 3202 -2478
rect 3352 -2542 3370 -2392
rect 3140 -2628 3370 -2542
rect 2928 -2630 3370 -2628
rect 2132 -2650 3370 -2630
rect 2132 -2652 2206 -2650
rect 3302 -2652 3370 -2650
rect 1144 -2702 1566 -2694
rect 1144 -2716 2038 -2702
rect 1144 -2726 1280 -2716
rect 1150 -2916 1280 -2726
rect 1480 -2718 2038 -2716
rect 1480 -2916 1586 -2718
rect 1150 -2918 1586 -2916
rect 1786 -2918 1866 -2718
rect 2028 -2918 2038 -2718
rect 1150 -2932 2038 -2918
rect 1270 -2934 2038 -2932
<< viali >>
rect -624 1266 -224 1658
rect 124 502 158 814
rect 212 502 246 814
rect 328 540 362 852
rect 416 852 450 854
rect 416 540 450 852
rect 736 510 770 822
rect 824 510 858 822
rect 940 548 974 860
rect 1028 860 1062 862
rect 1028 548 1062 860
rect -72 210 18 284
rect 124 92 158 216
rect 316 92 350 216
rect 1314 506 1348 818
rect 1402 506 1436 818
rect 1518 544 1552 856
rect 1606 856 1640 858
rect 1606 544 1640 856
rect 736 100 770 224
rect 928 100 962 224
rect 1888 514 1922 826
rect 1976 514 2010 826
rect 2092 552 2126 864
rect 2180 864 2214 866
rect 2180 552 2214 864
rect 1314 96 1348 220
rect 1506 96 1540 220
rect 2466 514 2500 826
rect 2554 514 2588 826
rect 2670 552 2704 864
rect 2758 864 2792 866
rect 2758 552 2792 864
rect 1888 104 1922 228
rect 2080 104 2114 228
rect 3044 514 3078 826
rect 3132 514 3166 826
rect 3248 552 3282 864
rect 3336 864 3370 866
rect 3336 552 3370 864
rect 2466 104 2500 228
rect 2658 104 2692 228
rect 3626 518 3660 830
rect 3714 518 3748 830
rect 3830 556 3864 868
rect 3918 868 3952 870
rect 3918 556 3952 868
rect 3044 104 3078 228
rect 3236 104 3270 228
rect 4202 514 4236 826
rect 4290 514 4324 826
rect 4406 552 4440 864
rect 4494 864 4528 866
rect 4494 552 4528 864
rect 4772 510 4806 822
rect 4860 510 4894 822
rect 4976 548 5010 860
rect 5064 860 5098 862
rect 5064 548 5098 860
rect 3626 108 3660 232
rect 3818 108 3852 232
rect 4202 104 4236 228
rect 4394 104 4428 228
rect 4558 32 4620 94
rect 4772 100 4806 224
rect 4964 100 4998 224
rect 5662 -234 6142 226
rect 1518 -1552 1552 -1240
rect 1606 -1552 1640 -1240
rect 1718 -1514 1752 -1202
rect 1806 -1514 1840 -1202
rect 1920 -1554 1954 -1242
rect 2008 -1554 2042 -1242
rect 1518 -2058 1552 -1746
rect 1606 -2058 1640 -1746
rect 1718 -2020 1752 -1708
rect 1806 -2020 1840 -1708
rect 1918 -2058 1952 -1746
rect 2006 -2058 2040 -1746
rect 1518 -2566 1552 -2254
rect 1606 -2566 1640 -2254
rect 1718 -2528 1752 -2216
rect 1806 -2528 1840 -2216
rect 1918 -2566 1952 -2254
rect 2006 -2566 2040 -2254
rect 3046 -2246 3080 -1622
<< metal1 >>
rect -650 1658 -170 1696
rect -650 1266 -624 1658
rect -224 1266 -170 1658
rect -650 1236 -170 1266
rect -556 1224 -240 1236
rect 212 896 458 928
rect 824 904 1070 936
rect 212 826 246 896
rect 416 868 456 896
rect 316 852 372 864
rect 112 816 170 826
rect 112 498 114 816
rect 166 498 170 816
rect 112 492 170 498
rect 200 814 260 826
rect 200 502 212 814
rect 246 710 260 814
rect 246 502 258 710
rect 316 540 320 852
rect 316 528 372 540
rect 406 854 462 868
rect 406 540 416 854
rect 450 540 462 854
rect 824 834 858 904
rect 1028 876 1068 904
rect 1402 900 1648 932
rect 1976 908 2222 940
rect 2554 908 2800 940
rect 3132 908 3378 940
rect 3714 912 3960 944
rect 928 860 984 872
rect 406 526 462 540
rect 724 824 782 834
rect 124 488 158 492
rect 200 490 258 502
rect -84 284 34 300
rect -84 210 -72 284
rect 18 210 34 284
rect -84 196 34 210
rect 112 222 174 228
rect 112 80 174 88
rect 300 216 362 228
rect 300 92 316 216
rect 350 186 362 216
rect 416 202 452 526
rect 724 506 726 824
rect 778 506 782 824
rect 724 500 782 506
rect 812 822 872 834
rect 812 510 824 822
rect 858 718 872 822
rect 858 510 870 718
rect 928 548 932 860
rect 928 536 984 548
rect 1018 862 1074 876
rect 1018 548 1028 862
rect 1062 548 1074 862
rect 1402 830 1436 900
rect 1606 872 1646 900
rect 1506 856 1562 868
rect 1018 534 1074 548
rect 1302 820 1360 830
rect 736 496 770 500
rect 812 498 870 510
rect 724 230 786 236
rect 416 186 458 202
rect 350 148 458 186
rect 350 92 362 148
rect 418 134 458 148
rect 300 80 362 92
rect 724 88 786 96
rect 912 224 974 236
rect 912 100 928 224
rect 962 194 974 224
rect 1028 206 1064 534
rect 1302 502 1304 820
rect 1356 502 1360 820
rect 1302 496 1360 502
rect 1390 818 1450 830
rect 1390 506 1402 818
rect 1436 714 1450 818
rect 1436 506 1448 714
rect 1506 544 1510 856
rect 1506 532 1562 544
rect 1596 858 1652 872
rect 1596 544 1606 858
rect 1640 544 1652 858
rect 1976 838 2010 908
rect 2180 880 2220 908
rect 2080 864 2136 876
rect 1596 530 1652 544
rect 1876 828 1934 838
rect 1314 492 1348 496
rect 1390 494 1448 506
rect 1302 226 1364 234
rect 1504 232 1538 236
rect 1028 194 1076 206
rect 962 156 1076 194
rect 962 100 974 156
rect 1036 138 1076 156
rect 912 88 974 100
rect 1302 78 1364 92
rect 1490 220 1552 232
rect 1490 96 1506 220
rect 1540 190 1552 220
rect 1606 204 1642 530
rect 1876 510 1878 828
rect 1930 510 1934 828
rect 1876 504 1934 510
rect 1964 826 2024 838
rect 1964 514 1976 826
rect 2010 722 2024 826
rect 2010 514 2022 722
rect 2080 552 2084 864
rect 2080 540 2136 552
rect 2170 866 2226 880
rect 2170 552 2180 866
rect 2214 552 2226 866
rect 2554 838 2588 908
rect 2758 880 2798 908
rect 2658 864 2714 876
rect 2170 538 2226 552
rect 2454 828 2512 838
rect 1888 500 1922 504
rect 1964 502 2022 514
rect 2070 240 2114 244
rect 1876 234 1938 240
rect 1606 190 1654 204
rect 1540 152 1654 190
rect 1540 96 1552 152
rect 1614 136 1654 152
rect 1490 84 1552 96
rect 1876 92 1938 100
rect 2064 228 2126 240
rect 2064 104 2080 228
rect 2114 198 2126 228
rect 2180 210 2216 538
rect 2454 510 2456 828
rect 2508 510 2512 828
rect 2454 504 2512 510
rect 2542 826 2602 838
rect 2542 514 2554 826
rect 2588 722 2602 826
rect 2588 514 2600 722
rect 2658 552 2662 864
rect 2658 540 2714 552
rect 2748 866 2804 880
rect 2748 552 2758 866
rect 2792 552 2804 866
rect 3132 838 3166 908
rect 3336 880 3376 908
rect 3236 864 3292 876
rect 2748 538 2804 552
rect 3032 828 3090 838
rect 2466 500 2500 504
rect 2542 502 2600 514
rect 2650 240 2696 244
rect 2454 234 2516 240
rect 2180 198 2226 210
rect 2114 160 2226 198
rect 2114 104 2126 160
rect 2184 152 2226 160
rect 2186 142 2226 152
rect 2064 92 2126 104
rect 2454 92 2516 100
rect 2642 228 2704 240
rect 2642 104 2658 228
rect 2692 198 2704 228
rect 2758 198 2794 538
rect 3032 510 3034 828
rect 3086 510 3090 828
rect 3032 504 3090 510
rect 3120 826 3180 838
rect 3120 514 3132 826
rect 3166 722 3180 826
rect 3166 514 3178 722
rect 3236 552 3240 864
rect 3236 540 3292 552
rect 3326 866 3382 880
rect 3326 552 3336 866
rect 3370 552 3382 866
rect 3714 842 3748 912
rect 3918 884 3958 912
rect 4290 908 4536 940
rect 3818 868 3874 880
rect 3326 538 3382 552
rect 3614 832 3672 842
rect 3044 500 3078 504
rect 3120 502 3178 514
rect 3232 240 3264 244
rect 2692 160 2794 198
rect 3032 234 3094 240
rect 2692 158 2790 160
rect 2692 104 2704 158
rect 2642 92 2704 104
rect 3032 92 3094 100
rect 3220 228 3282 240
rect 3220 104 3236 228
rect 3270 198 3282 228
rect 3336 198 3372 538
rect 3614 514 3616 832
rect 3668 514 3672 832
rect 3614 508 3672 514
rect 3702 830 3762 842
rect 3702 518 3714 830
rect 3748 726 3762 830
rect 3748 518 3760 726
rect 3818 556 3822 868
rect 3818 544 3874 556
rect 3908 870 3964 884
rect 3908 556 3918 870
rect 3952 556 3964 870
rect 4290 838 4324 908
rect 4494 880 4534 908
rect 4860 904 5106 936
rect 4394 864 4450 876
rect 3908 542 3964 556
rect 4190 828 4248 838
rect 3626 504 3660 508
rect 3702 506 3760 518
rect 3812 244 3850 248
rect 3270 160 3372 198
rect 3614 238 3676 244
rect 3270 104 3282 160
rect 3220 92 3282 104
rect 3614 96 3676 104
rect 3802 232 3864 244
rect 3802 108 3818 232
rect 3852 202 3864 232
rect 3918 214 3954 542
rect 4190 510 4192 828
rect 4244 510 4248 828
rect 4190 504 4248 510
rect 4278 826 4338 838
rect 4278 514 4290 826
rect 4324 722 4338 826
rect 4324 514 4336 722
rect 4394 552 4398 864
rect 4394 540 4450 552
rect 4484 866 4540 880
rect 4484 552 4494 866
rect 4528 552 4540 866
rect 4860 834 4894 904
rect 5064 876 5104 904
rect 4964 860 5020 872
rect 4484 538 4540 552
rect 4760 824 4818 834
rect 4202 500 4236 504
rect 4278 502 4336 514
rect 4388 240 4426 244
rect 4190 234 4252 240
rect 3918 202 3960 214
rect 3852 164 3960 202
rect 3852 108 3864 164
rect 3926 156 3960 164
rect 3802 96 3864 108
rect 4190 92 4252 100
rect 4378 228 4440 240
rect 4378 104 4394 228
rect 4428 198 4440 228
rect 4494 214 4530 538
rect 4760 506 4762 824
rect 4814 506 4818 824
rect 4760 500 4818 506
rect 4848 822 4908 834
rect 4848 510 4860 822
rect 4894 718 4908 822
rect 4894 510 4906 718
rect 4964 548 4968 860
rect 4964 536 5020 548
rect 5054 862 5110 876
rect 5054 548 5064 862
rect 5098 548 5110 862
rect 5054 534 5110 548
rect 4772 496 4806 500
rect 4848 498 4906 510
rect 4760 230 4822 236
rect 4494 198 4534 214
rect 4428 160 4534 198
rect 4428 104 4440 160
rect 4500 156 4534 160
rect 4378 92 4440 104
rect 4544 94 4634 110
rect 4544 32 4558 94
rect 4620 32 4634 94
rect 4760 88 4822 96
rect 4948 224 5010 236
rect 4948 100 4964 224
rect 4998 194 5010 224
rect 5064 214 5100 534
rect 5602 226 6214 294
rect 5064 194 5108 214
rect 4998 156 5108 194
rect 4998 100 5010 156
rect 4948 88 5010 100
rect 5602 84 5662 226
rect 4544 18 4634 32
rect 5490 -6 5662 84
rect 5602 -234 5662 -6
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
rect 1592 -1074 1768 -1072
rect 1592 -1076 1910 -1074
rect 1592 -1120 2060 -1076
rect 1592 -1134 2058 -1120
rect 1506 -1240 1564 -1228
rect 1506 -1552 1508 -1240
rect 1562 -1552 1564 -1240
rect 1592 -1240 1654 -1134
rect 1734 -1136 2058 -1134
rect 1792 -1138 2058 -1136
rect 1792 -1190 1850 -1138
rect 1592 -1252 1606 -1240
rect 1506 -1564 1564 -1552
rect 1594 -1552 1606 -1252
rect 1640 -1252 1654 -1240
rect 1706 -1202 1764 -1190
rect 1640 -1552 1652 -1252
rect 1706 -1514 1708 -1202
rect 1762 -1514 1764 -1202
rect 1792 -1202 1852 -1190
rect 1792 -1256 1806 -1202
rect 1706 -1526 1764 -1514
rect 1794 -1514 1806 -1256
rect 1840 -1514 1852 -1202
rect 2000 -1228 2058 -1138
rect 1506 -1746 1564 -1734
rect 1506 -2058 1508 -1746
rect 1562 -2058 1564 -1746
rect 1506 -2070 1564 -2058
rect 1594 -1746 1652 -1552
rect 1594 -2058 1606 -1746
rect 1640 -2058 1652 -1746
rect 1706 -1708 1764 -1696
rect 1706 -2020 1708 -1708
rect 1762 -2020 1764 -1708
rect 1706 -2032 1764 -2020
rect 1794 -1708 1852 -1514
rect 1908 -1242 1966 -1230
rect 1908 -1554 1910 -1242
rect 1964 -1554 1966 -1242
rect 1908 -1566 1966 -1554
rect 1994 -1242 2058 -1228
rect 1994 -1554 2008 -1242
rect 2042 -1266 2058 -1242
rect 2042 -1554 2052 -1266
rect 1794 -2020 1806 -1708
rect 1840 -2020 1852 -1708
rect 1994 -1688 2052 -1554
rect 3030 -1622 3092 -1610
rect 3030 -1688 3046 -1622
rect 1994 -1728 3046 -1688
rect 1506 -2254 1564 -2242
rect 1506 -2566 1508 -2254
rect 1562 -2566 1564 -2254
rect 1506 -2578 1564 -2566
rect 1594 -2254 1652 -2058
rect 1594 -2566 1606 -2254
rect 1640 -2566 1652 -2254
rect 1706 -2216 1764 -2204
rect 1706 -2528 1708 -2216
rect 1762 -2528 1764 -2216
rect 1706 -2540 1764 -2528
rect 1794 -2216 1852 -2020
rect 1906 -1746 1964 -1734
rect 1906 -2058 1908 -1746
rect 1962 -2058 1964 -1746
rect 1906 -2070 1964 -2058
rect 1994 -1746 2052 -1728
rect 2082 -1730 2136 -1728
rect 1994 -2058 2006 -1746
rect 2040 -2058 2052 -1746
rect 1794 -2528 1806 -2216
rect 1840 -2528 1852 -2216
rect 1794 -2540 1852 -2528
rect 1906 -2254 1964 -2242
rect 1594 -2578 1652 -2566
rect 1906 -2566 1908 -2254
rect 1962 -2566 1964 -2254
rect 1906 -2578 1964 -2566
rect 1994 -2254 2052 -2058
rect 1994 -2566 2006 -2254
rect 2040 -2566 2052 -2254
rect 3030 -2246 3046 -1728
rect 3080 -2246 3092 -1622
rect 3030 -2258 3092 -2246
rect 1994 -2578 2052 -2566
<< via1 >>
rect -624 1266 -224 1658
rect 114 814 166 816
rect 114 502 124 814
rect 124 502 158 814
rect 158 502 166 814
rect 114 498 166 502
rect 320 540 328 852
rect 328 540 362 852
rect 362 540 372 852
rect -72 210 18 284
rect 112 216 174 222
rect 112 92 124 216
rect 124 92 158 216
rect 158 92 174 216
rect 112 88 174 92
rect 726 822 778 824
rect 726 510 736 822
rect 736 510 770 822
rect 770 510 778 822
rect 726 506 778 510
rect 932 548 940 860
rect 940 548 974 860
rect 974 548 984 860
rect 724 224 786 230
rect 724 100 736 224
rect 736 100 770 224
rect 770 100 786 224
rect 724 96 786 100
rect 1304 818 1356 820
rect 1304 506 1314 818
rect 1314 506 1348 818
rect 1348 506 1356 818
rect 1304 502 1356 506
rect 1510 544 1518 856
rect 1518 544 1552 856
rect 1552 544 1562 856
rect 1302 220 1364 226
rect 1302 96 1314 220
rect 1314 96 1348 220
rect 1348 96 1364 220
rect 1302 92 1364 96
rect 1878 826 1930 828
rect 1878 514 1888 826
rect 1888 514 1922 826
rect 1922 514 1930 826
rect 1878 510 1930 514
rect 2084 552 2092 864
rect 2092 552 2126 864
rect 2126 552 2136 864
rect 1876 228 1938 234
rect 1876 104 1888 228
rect 1888 104 1922 228
rect 1922 104 1938 228
rect 1876 100 1938 104
rect 2456 826 2508 828
rect 2456 514 2466 826
rect 2466 514 2500 826
rect 2500 514 2508 826
rect 2456 510 2508 514
rect 2662 552 2670 864
rect 2670 552 2704 864
rect 2704 552 2714 864
rect 2454 228 2516 234
rect 2454 104 2466 228
rect 2466 104 2500 228
rect 2500 104 2516 228
rect 2454 100 2516 104
rect 3034 826 3086 828
rect 3034 514 3044 826
rect 3044 514 3078 826
rect 3078 514 3086 826
rect 3034 510 3086 514
rect 3240 552 3248 864
rect 3248 552 3282 864
rect 3282 552 3292 864
rect 3032 228 3094 234
rect 3032 104 3044 228
rect 3044 104 3078 228
rect 3078 104 3094 228
rect 3032 100 3094 104
rect 3616 830 3668 832
rect 3616 518 3626 830
rect 3626 518 3660 830
rect 3660 518 3668 830
rect 3616 514 3668 518
rect 3822 556 3830 868
rect 3830 556 3864 868
rect 3864 556 3874 868
rect 3614 232 3676 238
rect 3614 108 3626 232
rect 3626 108 3660 232
rect 3660 108 3676 232
rect 3614 104 3676 108
rect 4192 826 4244 828
rect 4192 514 4202 826
rect 4202 514 4236 826
rect 4236 514 4244 826
rect 4192 510 4244 514
rect 4398 552 4406 864
rect 4406 552 4440 864
rect 4440 552 4450 864
rect 4190 228 4252 234
rect 4190 104 4202 228
rect 4202 104 4236 228
rect 4236 104 4252 228
rect 4190 100 4252 104
rect 4762 822 4814 824
rect 4762 510 4772 822
rect 4772 510 4806 822
rect 4806 510 4814 822
rect 4762 506 4814 510
rect 4968 548 4976 860
rect 4976 548 5010 860
rect 5010 548 5020 860
rect 4760 224 4822 230
rect 4558 32 4620 94
rect 4760 100 4772 224
rect 4772 100 4806 224
rect 4806 100 4822 224
rect 4760 96 4822 100
rect 5662 -234 6142 226
rect 1508 -1552 1518 -1240
rect 1518 -1552 1552 -1240
rect 1552 -1552 1562 -1240
rect 1708 -1514 1718 -1202
rect 1718 -1514 1752 -1202
rect 1752 -1514 1762 -1202
rect 1508 -2058 1518 -1746
rect 1518 -2058 1552 -1746
rect 1552 -2058 1562 -1746
rect 1708 -2020 1718 -1708
rect 1718 -2020 1752 -1708
rect 1752 -2020 1762 -1708
rect 1910 -1554 1920 -1242
rect 1920 -1554 1954 -1242
rect 1954 -1554 1964 -1242
rect 1508 -2566 1518 -2254
rect 1518 -2566 1552 -2254
rect 1552 -2566 1562 -2254
rect 1708 -2528 1718 -2216
rect 1718 -2528 1752 -2216
rect 1752 -2528 1762 -2216
rect 1908 -2058 1918 -1746
rect 1918 -2058 1952 -1746
rect 1952 -2058 1962 -1746
rect 1908 -2566 1918 -2254
rect 1918 -2566 1952 -2254
rect 1952 -2566 1962 -2254
<< metal2 >>
rect -650 1658 -170 1696
rect -650 1266 -624 1658
rect -224 1292 -170 1658
rect -224 1266 -162 1292
rect -650 1262 -162 1266
rect -650 1236 -288 1262
rect -556 1194 -288 1236
rect -554 1184 -288 1194
rect 40 1184 4934 1196
rect -554 1114 4934 1184
rect 112 826 170 1114
rect 316 852 374 864
rect 110 816 172 826
rect 110 498 114 816
rect 166 578 172 816
rect 316 578 320 852
rect 166 540 320 578
rect 372 540 374 852
rect 166 538 374 540
rect 166 498 172 538
rect 316 528 374 538
rect 722 824 784 1114
rect 110 490 172 498
rect 722 506 726 824
rect 778 586 784 824
rect 928 860 986 872
rect 928 586 932 860
rect 778 548 932 586
rect 984 548 986 860
rect 1302 830 1360 1114
rect 1506 856 1564 868
rect 778 546 986 548
rect 778 506 784 546
rect 928 536 986 546
rect 1300 820 1362 830
rect 722 496 784 506
rect 1300 502 1304 820
rect 1356 582 1362 820
rect 1506 582 1510 856
rect 1356 544 1510 582
rect 1562 544 1564 856
rect 1356 542 1564 544
rect 1356 502 1362 542
rect 1506 532 1564 542
rect 1870 828 1938 1114
rect 1300 494 1362 502
rect 1870 510 1878 828
rect 1930 590 1938 828
rect 2080 864 2138 876
rect 2080 590 2084 864
rect 1930 552 2084 590
rect 2136 552 2138 864
rect 1930 550 2138 552
rect 1930 510 1938 550
rect 2080 540 2138 550
rect 2450 828 2514 1114
rect 1870 498 1938 510
rect 2450 510 2456 828
rect 2508 590 2514 828
rect 2658 864 2716 876
rect 2658 590 2662 864
rect 2508 552 2662 590
rect 2714 552 2716 864
rect 2508 550 2716 552
rect 2508 510 2514 550
rect 2658 540 2716 550
rect 3026 838 3088 1114
rect 3236 864 3294 876
rect 3026 828 3092 838
rect 2450 502 2514 510
rect 3026 510 3034 828
rect 3086 590 3092 828
rect 3236 590 3240 864
rect 3086 552 3240 590
rect 3292 552 3294 864
rect 3086 550 3294 552
rect 3086 510 3092 550
rect 3236 540 3294 550
rect 3606 842 3668 1114
rect 3818 868 3876 880
rect 3606 832 3674 842
rect 3026 502 3092 510
rect 3606 514 3616 832
rect 3668 594 3674 832
rect 3818 594 3822 868
rect 3668 556 3822 594
rect 3874 556 3876 868
rect 3668 554 3876 556
rect 3668 514 3674 554
rect 3818 544 3876 554
rect 4188 838 4244 1114
rect 4394 864 4452 876
rect 4188 828 4250 838
rect 3606 506 3674 514
rect 4188 510 4192 828
rect 4244 590 4250 828
rect 4394 590 4398 864
rect 4244 552 4398 590
rect 4450 552 4452 864
rect 4244 550 4452 552
rect 4244 510 4250 550
rect 4394 540 4452 550
rect 4758 824 4820 1114
rect 3026 494 3088 502
rect 3606 500 3668 506
rect 4188 502 4250 510
rect 4758 506 4762 824
rect 4814 586 4820 824
rect 4964 860 5022 872
rect 4964 586 4968 860
rect 4814 548 4968 586
rect 5020 548 5022 860
rect 4814 546 5022 548
rect 4814 506 4820 546
rect 4964 536 5022 546
rect 4188 494 4244 502
rect 4758 496 4820 506
rect 112 488 170 490
rect -84 284 34 300
rect -84 210 -72 284
rect 18 210 34 284
rect 3614 244 3674 246
rect 3032 240 3092 242
rect 114 230 174 232
rect -84 196 34 210
rect 110 222 174 230
rect 110 88 112 222
rect 110 -30 174 88
rect 724 230 786 236
rect 1874 234 1938 240
rect 724 88 786 96
rect 1302 226 1364 234
rect 724 -30 784 88
rect 1302 78 1364 92
rect 1874 100 1876 234
rect 1874 92 1938 100
rect 2454 234 2516 240
rect 1874 90 1936 92
rect 1302 -30 1362 78
rect 1874 -30 1934 90
rect 2454 82 2516 100
rect 2456 -30 2516 82
rect 3032 234 3094 240
rect 3032 92 3094 100
rect 3614 238 3676 244
rect 3614 96 3676 104
rect 4190 234 4252 240
rect 4772 236 4820 238
rect 4760 230 4822 236
rect 3032 -30 3092 92
rect 3614 -30 3674 96
rect 4190 88 4252 100
rect 4192 -30 4252 88
rect 4544 94 4634 110
rect 4544 32 4558 94
rect 4620 32 4634 94
rect 4544 18 4634 32
rect 4760 88 4822 96
rect 5602 226 6214 294
rect 110 -32 4536 -30
rect 4760 -32 4820 88
rect 5602 84 5662 226
rect 5068 -10 5662 84
rect 5068 -32 5140 -10
rect 110 -82 5140 -32
rect 4534 -84 5140 -82
rect 5068 -86 5140 -84
rect 5602 -234 5662 -10
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
rect 1706 -1202 1766 -1190
rect 1504 -1240 1564 -1226
rect 1504 -1552 1508 -1240
rect 1562 -1272 1564 -1240
rect 1706 -1272 1708 -1202
rect 1562 -1326 1708 -1272
rect 1562 -1552 1564 -1326
rect 1504 -1746 1564 -1552
rect 1504 -2058 1508 -1746
rect 1562 -1952 1564 -1746
rect 1706 -1514 1708 -1326
rect 1762 -1272 1766 -1202
rect 1906 -1242 1966 -1230
rect 1906 -1272 1910 -1242
rect 1762 -1326 1910 -1272
rect 1762 -1514 1766 -1326
rect 1706 -1708 1766 -1514
rect 1706 -1952 1708 -1708
rect 1562 -2006 1708 -1952
rect 1562 -2058 1564 -2006
rect 1504 -2254 1564 -2058
rect 1504 -2396 1508 -2254
rect 1500 -2450 1508 -2396
rect 1504 -2566 1508 -2450
rect 1562 -2396 1564 -2254
rect 1706 -2020 1708 -2006
rect 1762 -1952 1766 -1708
rect 1906 -1554 1910 -1326
rect 1964 -1272 1966 -1242
rect 1964 -1326 1968 -1272
rect 1964 -1554 1966 -1326
rect 1906 -1746 1966 -1554
rect 1906 -1952 1908 -1746
rect 1762 -2006 1908 -1952
rect 1762 -2020 1766 -2006
rect 1706 -2216 1766 -2020
rect 1706 -2394 1708 -2216
rect 1704 -2396 1708 -2394
rect 1562 -2450 1708 -2396
rect 1562 -2566 1564 -2450
rect 1706 -2528 1708 -2450
rect 1762 -2394 1766 -2216
rect 1906 -2058 1908 -2006
rect 1962 -2058 1966 -1746
rect 1906 -2254 1966 -2058
rect 1906 -2394 1908 -2254
rect 1762 -2448 1908 -2394
rect 1762 -2528 1766 -2448
rect 1706 -2540 1766 -2528
rect 1504 -2582 1564 -2566
rect 1906 -2566 1908 -2448
rect 1962 -2566 1966 -2254
rect 1906 -2580 1966 -2566
<< via2 >>
rect -624 1266 -224 1658
rect -72 210 18 284
rect 4558 32 4620 94
rect 5662 -234 6142 226
<< metal3 >>
rect -656 1658 -166 1696
rect -656 1266 -624 1658
rect -224 1266 -166 1658
rect -656 1236 -166 1266
rect -84 284 34 302
rect -84 210 -72 284
rect 18 280 34 284
rect 18 220 4620 280
rect 18 210 34 220
rect -84 192 34 210
rect 4558 110 4620 220
rect 5602 226 6214 294
rect 4544 94 4634 110
rect 4544 32 4558 94
rect 4620 32 4634 94
rect 4544 18 4634 32
rect 5602 -234 5662 226
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
<< via3 >>
rect -624 1266 -224 1658
rect 5662 -234 6142 226
<< metal4 >>
rect -656 1658 -166 1696
rect -656 1266 -624 1658
rect -224 1266 -166 1658
rect -656 1236 -166 1266
rect 5602 226 6214 294
rect 5602 -234 5662 226
rect 6142 -234 6214 226
rect 5602 -304 6214 -234
<< metal5 >>
rect -656 1236 -166 1696
<< labels >>
flabel via3 5862 -40 5862 -40 0 FreeSans 1600 0 0 0 GND!
flabel viali -30 262 -30 262 0 FreeSans 400 0 0 0 n1
flabel locali 232 146 232 146 0 FreeSans 400 0 0 0 net9
flabel locali 844 152 844 152 0 FreeSans 400 0 0 0 net8
flabel locali 1428 148 1428 148 0 FreeSans 400 0 0 0 net7
flabel locali 524 354 524 354 0 FreeSans 400 0 0 0 n2
flabel locali 1102 352 1102 352 0 FreeSans 400 0 0 0 n3
flabel locali 1680 354 1680 354 0 FreeSans 400 0 0 0 n4
flabel locali 2278 366 2278 366 0 FreeSans 400 0 0 0 n5
flabel locali 2856 368 2856 368 0 FreeSans 400 0 0 0 n6
flabel locali 3424 376 3424 376 0 FreeSans 400 0 0 0 n7
flabel locali 4008 368 4008 368 0 FreeSans 400 0 0 0 n8
flabel locali 4592 362 4592 362 0 FreeSans 400 0 0 0 n9
flabel locali 2004 156 2004 156 0 FreeSans 400 0 0 0 net1
flabel locali 2578 160 2578 160 0 FreeSans 400 0 0 0 net2
flabel locali 3154 158 3154 158 0 FreeSans 400 0 0 0 net3
flabel locali 3736 154 3736 154 0 FreeSans 400 0 0 0 net4
flabel locali 4322 148 4322 148 0 FreeSans 400 0 0 0 net5
flabel locali 4882 154 4882 154 0 FreeSans 400 0 0 0 net6
flabel metal1 434 172 434 172 0 FreeSans 400 0 0 0 v1!
flabel metal1 1048 178 1048 178 0 FreeSans 400 0 0 0 v2!
flabel metal1 1632 174 1632 174 0 FreeSans 400 0 0 0 v3!
flabel metal1 2198 180 2198 180 0 FreeSans 400 0 0 0 v4!
flabel metal1 3938 178 3938 178 0 FreeSans 400 0 0 0 v7!
flabel metal1 4510 186 4510 186 0 FreeSans 400 0 0 0 v8!
flabel metal1 5082 190 5082 190 0 FreeSans 400 0 0 0 v9!
flabel metal1 3350 184 3350 184 0 FreeSans 400 0 0 0 v6!
flabel metal1 2784 180 2784 180 0 FreeSans 400 0 0 0 v5!
flabel locali -844 1410 -844 1410 0 FreeSans 1600 0 0 0 VDD
flabel metal1 2108 -1718 2108 -1718 0 FreeSans 400 0 0 0 vout
flabel locali 1468 -2178 1468 -2178 0 FreeSans 400 0 0 0 v1!
flabel locali 1980 -2184 1980 -2184 0 FreeSans 400 0 0 0 v3!
flabel locali 1782 -2102 1782 -2102 0 FreeSans 400 0 0 0 v4!
flabel locali 1590 -1674 1590 -1674 0 FreeSans 400 0 0 0 v5!
flabel locali 1976 -1670 1976 -1670 0 FreeSans 400 0 0 0 v6!
flabel locali 1784 -1598 1784 -1598 0 FreeSans 400 0 0 0 v7!
flabel locali 3014 -2308 3014 -2308 0 FreeSans 400 0 0 0 v1!
flabel locali 2914 -1554 2914 -1554 0 FreeSans 400 0 0 0 v2!
flabel locali 2728 -1552 2728 -1552 0 FreeSans 400 0 0 0 v4!
flabel locali 2528 -1558 2528 -1558 0 FreeSans 400 0 0 0 v6!
flabel locali 2342 -1554 2342 -1554 0 FreeSans 400 0 0 0 v8!
flabel locali 2824 -2318 2824 -2318 0 FreeSans 400 0 0 0 v3!
flabel locali 2438 -2316 2438 -2316 0 FreeSans 400 0 0 0 v7!
flabel locali 2242 -2318 2242 -2318 0 FreeSans 400 0 0 0 v9!
flabel locali 2626 -2314 2626 -2314 0 FreeSans 400 0 0 0 v5!
flabel locali 2292 -1852 2292 -1852 0 FreeSans 400 0 0 0 net17!
flabel locali 2388 -1920 2388 -1920 0 FreeSans 400 0 0 0 net16!
flabel locali 2482 -1860 2482 -1860 0 FreeSans 400 0 0 0 net15!
flabel locali 2564 -1938 2564 -1938 0 FreeSans 400 0 0 0 net14!
flabel locali 2656 -1874 2656 -1874 0 FreeSans 400 0 0 0 net13!
flabel locali 2762 -1950 2762 -1950 0 FreeSans 400 0 0 0 net12!
flabel locali 2852 -1882 2852 -1882 0 FreeSans 400 0 0 0 net11!
flabel locali 2954 -1934 2954 -1934 0 FreeSans 400 0 0 0 net10!
flabel locali 1956 -1180 1956 -1180 0 FreeSans 400 0 0 0 v9!
flabel locali 1550 -1170 1550 -1170 0 FreeSans 400 0 0 0 v8!
flabel locali 1792 -2624 1792 -2624 0 FreeSans 400 0 0 0 v2!
<< end >>
