magic
tech sky130A
magscale 1 2
timestamp 1634912583
<< nwell >>
rect -34584 520 35722 18716
rect -34702 388 35722 520
rect -34722 186 35722 388
rect -34722 -922 -506 186
rect -246 156 35714 186
rect -246 122 648 156
rect -124 -36 648 122
rect -38 -414 648 -36
rect 454 -416 648 -414
rect 984 -610 35714 156
rect 984 -918 35736 -610
rect -34586 -924 -506 -922
<< nmos >>
rect 42 -748 72 -548
rect 138 -748 168 -548
rect 234 -748 264 -548
rect 330 -748 360 -548
<< pmos >>
rect 90 -304 120 96
rect 186 -304 216 96
rect 282 -304 312 96
rect 378 -304 408 96
<< pmoslvt >>
rect -32754 15374 -31154 16774
rect -31096 15374 -29496 16774
rect -29438 15374 -27838 16774
rect -27780 15374 -26180 16774
rect -26122 15374 -24522 16774
rect -24464 15374 -22864 16774
rect -22806 15374 -21206 16774
rect -21148 15374 -19548 16774
rect -19490 15374 -17890 16774
rect -17832 15374 -16232 16774
rect -16174 15374 -14574 16774
rect -14516 15374 -12916 16774
rect -12858 15374 -11258 16774
rect -11200 15374 -9600 16774
rect -9542 15374 -7942 16774
rect -7884 15374 -6284 16774
rect -6226 15374 -4626 16774
rect -4568 15374 -2968 16774
rect -2910 15374 -1310 16774
rect -1252 15374 348 16774
rect 406 15374 2006 16774
rect 2064 15374 3664 16774
rect 3722 15374 5322 16774
rect 5380 15374 6980 16774
rect 7038 15374 8638 16774
rect 8696 15374 10296 16774
rect 10354 15374 11954 16774
rect 12012 15374 13612 16774
rect 13670 15374 15270 16774
rect 15328 15374 16928 16774
rect 16986 15374 18586 16774
rect 18644 15374 20244 16774
rect 20302 15374 21902 16774
rect 21960 15374 23560 16774
rect 23618 15374 25218 16774
rect 25276 15374 26876 16774
rect 26934 15374 28534 16774
rect 28592 15374 30192 16774
rect 30250 15374 31850 16774
rect 31908 15374 33508 16774
rect -32754 13738 -31154 15138
rect -31096 13738 -29496 15138
rect -29438 13738 -27838 15138
rect -27780 13738 -26180 15138
rect -26122 13738 -24522 15138
rect -24464 13738 -22864 15138
rect -22806 13738 -21206 15138
rect -21148 13738 -19548 15138
rect -19490 13738 -17890 15138
rect -17832 13738 -16232 15138
rect -16174 13738 -14574 15138
rect -14516 13738 -12916 15138
rect -12858 13738 -11258 15138
rect -11200 13738 -9600 15138
rect -9542 13738 -7942 15138
rect -7884 13738 -6284 15138
rect -6226 13738 -4626 15138
rect -4568 13738 -2968 15138
rect -2910 13738 -1310 15138
rect -1252 13738 348 15138
rect 406 13738 2006 15138
rect 2064 13738 3664 15138
rect 3722 13738 5322 15138
rect 5380 13738 6980 15138
rect 7038 13738 8638 15138
rect 8696 13738 10296 15138
rect 10354 13738 11954 15138
rect 12012 13738 13612 15138
rect 13670 13738 15270 15138
rect 15328 13738 16928 15138
rect 16986 13738 18586 15138
rect 18644 13738 20244 15138
rect 20302 13738 21902 15138
rect 21960 13738 23560 15138
rect 23618 13738 25218 15138
rect 25276 13738 26876 15138
rect 26934 13738 28534 15138
rect 28592 13738 30192 15138
rect 30250 13738 31850 15138
rect 31908 13738 33508 15138
rect -32752 11992 -31152 13392
rect -31094 11992 -29494 13392
rect -29436 11992 -27836 13392
rect -27778 11992 -26178 13392
rect -26120 11992 -24520 13392
rect -24462 11992 -22862 13392
rect -22804 11992 -21204 13392
rect -21146 11992 -19546 13392
rect -19488 11992 -17888 13392
rect -17830 11992 -16230 13392
rect -16172 11992 -14572 13392
rect -14514 11992 -12914 13392
rect -12856 11992 -11256 13392
rect -11198 11992 -9598 13392
rect -9540 11992 -7940 13392
rect -7882 11992 -6282 13392
rect -6224 11992 -4624 13392
rect -4566 11992 -2966 13392
rect -2908 11992 -1308 13392
rect -1250 11992 350 13392
rect 408 11992 2008 13392
rect 2066 11992 3666 13392
rect 3724 11992 5324 13392
rect 5382 11992 6982 13392
rect 7040 11992 8640 13392
rect 8698 11992 10298 13392
rect 10356 11992 11956 13392
rect 12014 11992 13614 13392
rect 13672 11992 15272 13392
rect 15330 11992 16930 13392
rect 16988 11992 18588 13392
rect 18646 11992 20246 13392
rect 20304 11992 21904 13392
rect 21962 11992 23562 13392
rect 23620 11992 25220 13392
rect 25278 11992 26878 13392
rect 26936 11992 28536 13392
rect 28594 11992 30194 13392
rect 30252 11992 31852 13392
rect 31910 11992 33510 13392
rect -32752 10356 -31152 11756
rect -31094 10356 -29494 11756
rect -29436 10356 -27836 11756
rect -27778 10356 -26178 11756
rect -26120 10356 -24520 11756
rect -24462 10356 -22862 11756
rect -22804 10356 -21204 11756
rect -21146 10356 -19546 11756
rect -19488 10356 -17888 11756
rect -17830 10356 -16230 11756
rect -16172 10356 -14572 11756
rect -14514 10356 -12914 11756
rect -12856 10356 -11256 11756
rect -11198 10356 -9598 11756
rect -9540 10356 -7940 11756
rect -7882 10356 -6282 11756
rect -6224 10356 -4624 11756
rect -4566 10356 -2966 11756
rect -2908 10356 -1308 11756
rect -1250 10356 350 11756
rect 408 10356 2008 11756
rect 2066 10356 3666 11756
rect 3724 10356 5324 11756
rect 5382 10356 6982 11756
rect 7040 10356 8640 11756
rect 8698 10356 10298 11756
rect 10356 10356 11956 11756
rect 12014 10356 13614 11756
rect 13672 10356 15272 11756
rect 15330 10356 16930 11756
rect 16988 10356 18588 11756
rect 18646 10356 20246 11756
rect 20304 10356 21904 11756
rect 21962 10356 23562 11756
rect 23620 10356 25220 11756
rect 25278 10356 26878 11756
rect 26936 10356 28536 11756
rect 28594 10356 30194 11756
rect 30252 10356 31852 11756
rect 31910 10356 33510 11756
rect -32752 8720 -31152 10120
rect -31094 8720 -29494 10120
rect -29436 8720 -27836 10120
rect -27778 8720 -26178 10120
rect -26120 8720 -24520 10120
rect -24462 8720 -22862 10120
rect -22804 8720 -21204 10120
rect -21146 8720 -19546 10120
rect -19488 8720 -17888 10120
rect -17830 8720 -16230 10120
rect -16172 8720 -14572 10120
rect -14514 8720 -12914 10120
rect -12856 8720 -11256 10120
rect -11198 8720 -9598 10120
rect -9540 8720 -7940 10120
rect -7882 8720 -6282 10120
rect -6224 8720 -4624 10120
rect -4566 8720 -2966 10120
rect -2908 8720 -1308 10120
rect -1250 8720 350 10120
rect 408 8720 2008 10120
rect 2066 8720 3666 10120
rect 3724 8720 5324 10120
rect 5382 8720 6982 10120
rect 7040 8720 8640 10120
rect 8698 8720 10298 10120
rect 10356 8720 11956 10120
rect 12014 8720 13614 10120
rect 13672 8720 15272 10120
rect 15330 8720 16930 10120
rect 16988 8720 18588 10120
rect 18646 8720 20246 10120
rect 20304 8720 21904 10120
rect 21962 8720 23562 10120
rect 23620 8720 25220 10120
rect 25278 8720 26878 10120
rect 26936 8720 28536 10120
rect 28594 8720 30194 10120
rect 30252 8720 31852 10120
rect 31910 8720 33510 10120
rect -32752 7084 -31152 8484
rect -31094 7084 -29494 8484
rect -29436 7084 -27836 8484
rect -27778 7084 -26178 8484
rect -26120 7084 -24520 8484
rect -24462 7084 -22862 8484
rect -22804 7084 -21204 8484
rect -21146 7084 -19546 8484
rect -19488 7084 -17888 8484
rect -17830 7084 -16230 8484
rect -16172 7084 -14572 8484
rect -14514 7084 -12914 8484
rect -12856 7084 -11256 8484
rect -11198 7084 -9598 8484
rect -9540 7084 -7940 8484
rect -7882 7084 -6282 8484
rect -6224 7084 -4624 8484
rect -4566 7084 -2966 8484
rect -2908 7084 -1308 8484
rect -1250 7084 350 8484
rect 408 7084 2008 8484
rect 2066 7084 3666 8484
rect 3724 7084 5324 8484
rect 5382 7084 6982 8484
rect 7040 7084 8640 8484
rect 8698 7084 10298 8484
rect 10356 7084 11956 8484
rect 12014 7084 13614 8484
rect 13672 7084 15272 8484
rect 15330 7084 16930 8484
rect 16988 7084 18588 8484
rect 18646 7084 20246 8484
rect 20304 7084 21904 8484
rect 21962 7084 23562 8484
rect 23620 7084 25220 8484
rect 25278 7084 26878 8484
rect 26936 7084 28536 8484
rect 28594 7084 30194 8484
rect 30252 7084 31852 8484
rect 31910 7084 33510 8484
rect -32752 5446 -31152 6846
rect -31094 5446 -29494 6846
rect -29436 5446 -27836 6846
rect -27778 5446 -26178 6846
rect -26120 5446 -24520 6846
rect -24462 5446 -22862 6846
rect -22804 5446 -21204 6846
rect -21146 5446 -19546 6846
rect -19488 5446 -17888 6846
rect -17830 5446 -16230 6846
rect -16172 5446 -14572 6846
rect -14514 5446 -12914 6846
rect -12856 5446 -11256 6846
rect -11198 5446 -9598 6846
rect -9540 5446 -7940 6846
rect -7882 5446 -6282 6846
rect -6224 5446 -4624 6846
rect -4566 5446 -2966 6846
rect -2908 5446 -1308 6846
rect -1250 5446 350 6846
rect 408 5446 2008 6846
rect 2066 5446 3666 6846
rect 3724 5446 5324 6846
rect 5382 5446 6982 6846
rect 7040 5446 8640 6846
rect 8698 5446 10298 6846
rect 10356 5446 11956 6846
rect 12014 5446 13614 6846
rect 13672 5446 15272 6846
rect 15330 5446 16930 6846
rect 16988 5446 18588 6846
rect 18646 5446 20246 6846
rect 20304 5446 21904 6846
rect 21962 5446 23562 6846
rect 23620 5446 25220 6846
rect 25278 5446 26878 6846
rect 26936 5446 28536 6846
rect 28594 5446 30194 6846
rect 30252 5446 31852 6846
rect 31910 5446 33510 6846
rect -32752 3810 -31152 5210
rect -31094 3810 -29494 5210
rect -29436 3810 -27836 5210
rect -27778 3810 -26178 5210
rect -26120 3810 -24520 5210
rect -24462 3810 -22862 5210
rect -22804 3810 -21204 5210
rect -21146 3810 -19546 5210
rect -19488 3810 -17888 5210
rect -17830 3810 -16230 5210
rect -16172 3810 -14572 5210
rect -14514 3810 -12914 5210
rect -12856 3810 -11256 5210
rect -11198 3810 -9598 5210
rect -9540 3810 -7940 5210
rect -7882 3810 -6282 5210
rect -6224 3810 -4624 5210
rect -4566 3810 -2966 5210
rect -2908 3810 -1308 5210
rect -1250 3810 350 5210
rect 408 3810 2008 5210
rect 2066 3810 3666 5210
rect 3724 3810 5324 5210
rect 5382 3810 6982 5210
rect 7040 3810 8640 5210
rect 8698 3810 10298 5210
rect 10356 3810 11956 5210
rect 12014 3810 13614 5210
rect 13672 3810 15272 5210
rect 15330 3810 16930 5210
rect 16988 3810 18588 5210
rect 18646 3810 20246 5210
rect 20304 3810 21904 5210
rect 21962 3810 23562 5210
rect 23620 3810 25220 5210
rect 25278 3810 26878 5210
rect 26936 3810 28536 5210
rect 28594 3810 30194 5210
rect 30252 3810 31852 5210
rect 31910 3810 33510 5210
rect -32752 2174 -31152 3574
rect -31094 2174 -29494 3574
rect -29436 2174 -27836 3574
rect -27778 2174 -26178 3574
rect -26120 2174 -24520 3574
rect -24462 2174 -22862 3574
rect -22804 2174 -21204 3574
rect -21146 2174 -19546 3574
rect -19488 2174 -17888 3574
rect -17830 2174 -16230 3574
rect -16172 2174 -14572 3574
rect -14514 2174 -12914 3574
rect -12856 2174 -11256 3574
rect -11198 2174 -9598 3574
rect -9540 2174 -7940 3574
rect -7882 2174 -6282 3574
rect -6224 2174 -4624 3574
rect -4566 2174 -2966 3574
rect -2908 2174 -1308 3574
rect -1250 2174 350 3574
rect 408 2174 2008 3574
rect 2066 2174 3666 3574
rect 3724 2174 5324 3574
rect 5382 2174 6982 3574
rect 7040 2174 8640 3574
rect 8698 2174 10298 3574
rect 10356 2174 11956 3574
rect 12014 2174 13614 3574
rect 13672 2174 15272 3574
rect 15330 2174 16930 3574
rect 16988 2174 18588 3574
rect 18646 2174 20246 3574
rect 20304 2174 21904 3574
rect 21962 2174 23562 3574
rect 23620 2174 25220 3574
rect 25278 2174 26878 3574
rect 26936 2174 28536 3574
rect 28594 2174 30194 3574
rect 30252 2174 31852 3574
rect 31910 2174 33510 3574
rect -32752 538 -31152 1938
rect -31094 538 -29494 1938
rect -29436 538 -27836 1938
rect -27778 538 -26178 1938
rect -26120 538 -24520 1938
rect -24462 538 -22862 1938
rect -22804 538 -21204 1938
rect -21146 538 -19546 1938
rect -19488 538 -17888 1938
rect -17830 538 -16230 1938
rect -16172 538 -14572 1938
rect -14514 538 -12914 1938
rect -12856 538 -11256 1938
rect -11198 538 -9598 1938
rect -9540 538 -7940 1938
rect -7882 538 -6282 1938
rect -6224 538 -4624 1938
rect -4566 538 -2966 1938
rect -2908 538 -1308 1938
rect -1250 538 350 1938
rect 408 538 2008 1938
rect 2066 538 3666 1938
rect 3724 538 5324 1938
rect 5382 538 6982 1938
rect 7040 538 8640 1938
rect 8698 538 10298 1938
rect 10356 538 11956 1938
rect 12014 538 13614 1938
rect 13672 538 15272 1938
rect 15330 538 16930 1938
rect 16988 538 18588 1938
rect 18646 538 20246 1938
rect 20304 538 21904 1938
rect 21962 538 23562 1938
rect 23620 538 25220 1938
rect 25278 538 26878 1938
rect 26936 538 28536 1938
rect 28594 538 30194 1938
rect 30252 538 31852 1938
rect 31910 538 33510 1938
<< ndiff >>
rect -16 -592 42 -548
rect -20 -604 42 -592
rect -20 -692 -8 -604
rect 26 -692 42 -604
rect -20 -704 42 -692
rect -16 -748 42 -704
rect 72 -604 138 -548
rect 72 -692 88 -604
rect 122 -692 138 -604
rect 72 -748 138 -692
rect 168 -604 234 -548
rect 168 -692 184 -604
rect 218 -692 234 -604
rect 168 -748 234 -692
rect 264 -604 330 -548
rect 264 -692 280 -604
rect 314 -692 330 -604
rect 264 -748 330 -692
rect 360 -592 418 -548
rect 360 -604 422 -592
rect 360 -692 376 -604
rect 410 -692 422 -604
rect 360 -704 422 -692
rect 360 -748 418 -704
<< pdiff >>
rect -32812 16418 -32754 16774
rect -32812 15730 -32800 16418
rect -32766 15730 -32754 16418
rect -32812 15374 -32754 15730
rect -31154 16418 -31096 16774
rect -31154 15730 -31142 16418
rect -31108 15730 -31096 16418
rect -31154 15374 -31096 15730
rect -29496 16418 -29438 16774
rect -29496 15730 -29484 16418
rect -29450 15730 -29438 16418
rect -29496 15374 -29438 15730
rect -27838 16418 -27780 16774
rect -27838 15730 -27826 16418
rect -27792 15730 -27780 16418
rect -27838 15374 -27780 15730
rect -26180 16418 -26122 16774
rect -26180 15730 -26168 16418
rect -26134 15730 -26122 16418
rect -26180 15374 -26122 15730
rect -24522 16418 -24464 16774
rect -24522 15730 -24510 16418
rect -24476 15730 -24464 16418
rect -24522 15374 -24464 15730
rect -22864 16418 -22806 16774
rect -22864 15730 -22852 16418
rect -22818 15730 -22806 16418
rect -22864 15374 -22806 15730
rect -21206 16418 -21148 16774
rect -21206 15730 -21194 16418
rect -21160 15730 -21148 16418
rect -21206 15374 -21148 15730
rect -19548 16418 -19490 16774
rect -19548 15730 -19536 16418
rect -19502 15730 -19490 16418
rect -19548 15374 -19490 15730
rect -17890 16418 -17832 16774
rect -17890 15730 -17878 16418
rect -17844 15730 -17832 16418
rect -17890 15374 -17832 15730
rect -16232 16418 -16174 16774
rect -16232 15730 -16220 16418
rect -16186 15730 -16174 16418
rect -16232 15374 -16174 15730
rect -14574 16418 -14516 16774
rect -14574 15730 -14562 16418
rect -14528 15730 -14516 16418
rect -14574 15374 -14516 15730
rect -12916 16418 -12858 16774
rect -12916 15730 -12904 16418
rect -12870 15730 -12858 16418
rect -12916 15374 -12858 15730
rect -11258 16418 -11200 16774
rect -11258 15730 -11246 16418
rect -11212 15730 -11200 16418
rect -11258 15374 -11200 15730
rect -9600 16418 -9542 16774
rect -9600 15730 -9588 16418
rect -9554 15730 -9542 16418
rect -9600 15374 -9542 15730
rect -7942 16418 -7884 16774
rect -7942 15730 -7930 16418
rect -7896 15730 -7884 16418
rect -7942 15374 -7884 15730
rect -6284 16418 -6226 16774
rect -6284 15730 -6272 16418
rect -6238 15730 -6226 16418
rect -6284 15374 -6226 15730
rect -4626 16418 -4568 16774
rect -4626 15730 -4614 16418
rect -4580 15730 -4568 16418
rect -4626 15374 -4568 15730
rect -2968 16418 -2910 16774
rect -2968 15730 -2956 16418
rect -2922 15730 -2910 16418
rect -2968 15374 -2910 15730
rect -1310 16418 -1252 16774
rect -1310 15730 -1298 16418
rect -1264 15730 -1252 16418
rect -1310 15374 -1252 15730
rect 348 16418 406 16774
rect 348 15730 360 16418
rect 394 15730 406 16418
rect 348 15374 406 15730
rect 2006 16418 2064 16774
rect 2006 15730 2018 16418
rect 2052 15730 2064 16418
rect 2006 15374 2064 15730
rect 3664 16418 3722 16774
rect 3664 15730 3676 16418
rect 3710 15730 3722 16418
rect 3664 15374 3722 15730
rect 5322 16418 5380 16774
rect 5322 15730 5334 16418
rect 5368 15730 5380 16418
rect 5322 15374 5380 15730
rect 6980 16418 7038 16774
rect 6980 15730 6992 16418
rect 7026 15730 7038 16418
rect 6980 15374 7038 15730
rect 8638 16418 8696 16774
rect 8638 15730 8650 16418
rect 8684 15730 8696 16418
rect 8638 15374 8696 15730
rect 10296 16418 10354 16774
rect 10296 15730 10308 16418
rect 10342 15730 10354 16418
rect 10296 15374 10354 15730
rect 11954 16418 12012 16774
rect 11954 15730 11966 16418
rect 12000 15730 12012 16418
rect 11954 15374 12012 15730
rect 13612 16418 13670 16774
rect 13612 15730 13624 16418
rect 13658 15730 13670 16418
rect 13612 15374 13670 15730
rect 15270 16418 15328 16774
rect 15270 15730 15282 16418
rect 15316 15730 15328 16418
rect 15270 15374 15328 15730
rect 16928 16418 16986 16774
rect 16928 15730 16940 16418
rect 16974 15730 16986 16418
rect 16928 15374 16986 15730
rect 18586 16418 18644 16774
rect 18586 15730 18598 16418
rect 18632 15730 18644 16418
rect 18586 15374 18644 15730
rect 20244 16418 20302 16774
rect 20244 15730 20256 16418
rect 20290 15730 20302 16418
rect 20244 15374 20302 15730
rect 21902 16418 21960 16774
rect 21902 15730 21914 16418
rect 21948 15730 21960 16418
rect 21902 15374 21960 15730
rect 23560 16418 23618 16774
rect 23560 15730 23572 16418
rect 23606 15730 23618 16418
rect 23560 15374 23618 15730
rect 25218 16418 25276 16774
rect 25218 15730 25230 16418
rect 25264 15730 25276 16418
rect 25218 15374 25276 15730
rect 26876 16418 26934 16774
rect 26876 15730 26888 16418
rect 26922 15730 26934 16418
rect 26876 15374 26934 15730
rect 28534 16418 28592 16774
rect 28534 15730 28546 16418
rect 28580 15730 28592 16418
rect 28534 15374 28592 15730
rect 30192 16418 30250 16774
rect 30192 15730 30204 16418
rect 30238 15730 30250 16418
rect 30192 15374 30250 15730
rect 31850 16418 31908 16774
rect 31850 15730 31862 16418
rect 31896 15730 31908 16418
rect 31850 15374 31908 15730
rect 33508 16418 33566 16774
rect 33508 15730 33520 16418
rect 33554 15730 33566 16418
rect 33508 15374 33566 15730
rect -32812 14782 -32754 15138
rect -32812 14094 -32800 14782
rect -32766 14094 -32754 14782
rect -32812 13738 -32754 14094
rect -31154 14782 -31096 15138
rect -31154 14094 -31142 14782
rect -31108 14094 -31096 14782
rect -31154 13738 -31096 14094
rect -29496 14782 -29438 15138
rect -29496 14094 -29484 14782
rect -29450 14094 -29438 14782
rect -29496 13738 -29438 14094
rect -27838 14782 -27780 15138
rect -27838 14094 -27826 14782
rect -27792 14094 -27780 14782
rect -27838 13738 -27780 14094
rect -26180 14782 -26122 15138
rect -26180 14094 -26168 14782
rect -26134 14094 -26122 14782
rect -26180 13738 -26122 14094
rect -24522 14782 -24464 15138
rect -24522 14094 -24510 14782
rect -24476 14094 -24464 14782
rect -24522 13738 -24464 14094
rect -22864 14782 -22806 15138
rect -22864 14094 -22852 14782
rect -22818 14094 -22806 14782
rect -22864 13738 -22806 14094
rect -21206 14782 -21148 15138
rect -21206 14094 -21194 14782
rect -21160 14094 -21148 14782
rect -21206 13738 -21148 14094
rect -19548 14782 -19490 15138
rect -19548 14094 -19536 14782
rect -19502 14094 -19490 14782
rect -19548 13738 -19490 14094
rect -17890 14782 -17832 15138
rect -17890 14094 -17878 14782
rect -17844 14094 -17832 14782
rect -17890 13738 -17832 14094
rect -16232 14782 -16174 15138
rect -16232 14094 -16220 14782
rect -16186 14094 -16174 14782
rect -16232 13738 -16174 14094
rect -14574 14782 -14516 15138
rect -14574 14094 -14562 14782
rect -14528 14094 -14516 14782
rect -14574 13738 -14516 14094
rect -12916 14782 -12858 15138
rect -12916 14094 -12904 14782
rect -12870 14094 -12858 14782
rect -12916 13738 -12858 14094
rect -11258 14782 -11200 15138
rect -11258 14094 -11246 14782
rect -11212 14094 -11200 14782
rect -11258 13738 -11200 14094
rect -9600 14782 -9542 15138
rect -9600 14094 -9588 14782
rect -9554 14094 -9542 14782
rect -9600 13738 -9542 14094
rect -7942 14782 -7884 15138
rect -7942 14094 -7930 14782
rect -7896 14094 -7884 14782
rect -7942 13738 -7884 14094
rect -6284 14782 -6226 15138
rect -6284 14094 -6272 14782
rect -6238 14094 -6226 14782
rect -6284 13738 -6226 14094
rect -4626 14782 -4568 15138
rect -4626 14094 -4614 14782
rect -4580 14094 -4568 14782
rect -4626 13738 -4568 14094
rect -2968 14782 -2910 15138
rect -2968 14094 -2956 14782
rect -2922 14094 -2910 14782
rect -2968 13738 -2910 14094
rect -1310 14782 -1252 15138
rect -1310 14094 -1298 14782
rect -1264 14094 -1252 14782
rect -1310 13738 -1252 14094
rect 348 14782 406 15138
rect 348 14094 360 14782
rect 394 14094 406 14782
rect 348 13738 406 14094
rect 2006 14782 2064 15138
rect 2006 14094 2018 14782
rect 2052 14094 2064 14782
rect 2006 13738 2064 14094
rect 3664 14782 3722 15138
rect 3664 14094 3676 14782
rect 3710 14094 3722 14782
rect 3664 13738 3722 14094
rect 5322 14782 5380 15138
rect 5322 14094 5334 14782
rect 5368 14094 5380 14782
rect 5322 13738 5380 14094
rect 6980 14782 7038 15138
rect 6980 14094 6992 14782
rect 7026 14094 7038 14782
rect 6980 13738 7038 14094
rect 8638 14782 8696 15138
rect 8638 14094 8650 14782
rect 8684 14094 8696 14782
rect 8638 13738 8696 14094
rect 10296 14782 10354 15138
rect 10296 14094 10308 14782
rect 10342 14094 10354 14782
rect 10296 13738 10354 14094
rect 11954 14782 12012 15138
rect 11954 14094 11966 14782
rect 12000 14094 12012 14782
rect 11954 13738 12012 14094
rect 13612 14782 13670 15138
rect 13612 14094 13624 14782
rect 13658 14094 13670 14782
rect 13612 13738 13670 14094
rect 15270 14782 15328 15138
rect 15270 14094 15282 14782
rect 15316 14094 15328 14782
rect 15270 13738 15328 14094
rect 16928 14782 16986 15138
rect 16928 14094 16940 14782
rect 16974 14094 16986 14782
rect 16928 13738 16986 14094
rect 18586 14782 18644 15138
rect 18586 14094 18598 14782
rect 18632 14094 18644 14782
rect 18586 13738 18644 14094
rect 20244 14782 20302 15138
rect 20244 14094 20256 14782
rect 20290 14094 20302 14782
rect 20244 13738 20302 14094
rect 21902 14782 21960 15138
rect 21902 14094 21914 14782
rect 21948 14094 21960 14782
rect 21902 13738 21960 14094
rect 23560 14782 23618 15138
rect 23560 14094 23572 14782
rect 23606 14094 23618 14782
rect 23560 13738 23618 14094
rect 25218 14782 25276 15138
rect 25218 14094 25230 14782
rect 25264 14094 25276 14782
rect 25218 13738 25276 14094
rect 26876 14782 26934 15138
rect 26876 14094 26888 14782
rect 26922 14094 26934 14782
rect 26876 13738 26934 14094
rect 28534 14782 28592 15138
rect 28534 14094 28546 14782
rect 28580 14094 28592 14782
rect 28534 13738 28592 14094
rect 30192 14782 30250 15138
rect 30192 14094 30204 14782
rect 30238 14094 30250 14782
rect 30192 13738 30250 14094
rect 31850 14782 31908 15138
rect 31850 14094 31862 14782
rect 31896 14094 31908 14782
rect 31850 13738 31908 14094
rect 33508 14782 33566 15138
rect 33508 14094 33520 14782
rect 33554 14094 33566 14782
rect 33508 13738 33566 14094
rect -32810 13036 -32752 13392
rect -32810 12348 -32798 13036
rect -32764 12348 -32752 13036
rect -32810 11992 -32752 12348
rect -31152 13036 -31094 13392
rect -31152 12348 -31140 13036
rect -31106 12348 -31094 13036
rect -31152 11992 -31094 12348
rect -29494 13036 -29436 13392
rect -29494 12348 -29482 13036
rect -29448 12348 -29436 13036
rect -29494 11992 -29436 12348
rect -27836 13036 -27778 13392
rect -27836 12348 -27824 13036
rect -27790 12348 -27778 13036
rect -27836 11992 -27778 12348
rect -26178 13036 -26120 13392
rect -26178 12348 -26166 13036
rect -26132 12348 -26120 13036
rect -26178 11992 -26120 12348
rect -24520 13036 -24462 13392
rect -24520 12348 -24508 13036
rect -24474 12348 -24462 13036
rect -24520 11992 -24462 12348
rect -22862 13036 -22804 13392
rect -22862 12348 -22850 13036
rect -22816 12348 -22804 13036
rect -22862 11992 -22804 12348
rect -21204 13036 -21146 13392
rect -21204 12348 -21192 13036
rect -21158 12348 -21146 13036
rect -21204 11992 -21146 12348
rect -19546 13036 -19488 13392
rect -19546 12348 -19534 13036
rect -19500 12348 -19488 13036
rect -19546 11992 -19488 12348
rect -17888 13036 -17830 13392
rect -17888 12348 -17876 13036
rect -17842 12348 -17830 13036
rect -17888 11992 -17830 12348
rect -16230 13036 -16172 13392
rect -16230 12348 -16218 13036
rect -16184 12348 -16172 13036
rect -16230 11992 -16172 12348
rect -14572 13036 -14514 13392
rect -14572 12348 -14560 13036
rect -14526 12348 -14514 13036
rect -14572 11992 -14514 12348
rect -12914 13036 -12856 13392
rect -12914 12348 -12902 13036
rect -12868 12348 -12856 13036
rect -12914 11992 -12856 12348
rect -11256 13036 -11198 13392
rect -11256 12348 -11244 13036
rect -11210 12348 -11198 13036
rect -11256 11992 -11198 12348
rect -9598 13036 -9540 13392
rect -9598 12348 -9586 13036
rect -9552 12348 -9540 13036
rect -9598 11992 -9540 12348
rect -7940 13036 -7882 13392
rect -7940 12348 -7928 13036
rect -7894 12348 -7882 13036
rect -7940 11992 -7882 12348
rect -6282 13036 -6224 13392
rect -6282 12348 -6270 13036
rect -6236 12348 -6224 13036
rect -6282 11992 -6224 12348
rect -4624 13036 -4566 13392
rect -4624 12348 -4612 13036
rect -4578 12348 -4566 13036
rect -4624 11992 -4566 12348
rect -2966 13036 -2908 13392
rect -2966 12348 -2954 13036
rect -2920 12348 -2908 13036
rect -2966 11992 -2908 12348
rect -1308 13036 -1250 13392
rect -1308 12348 -1296 13036
rect -1262 12348 -1250 13036
rect -1308 11992 -1250 12348
rect 350 13036 408 13392
rect 350 12348 362 13036
rect 396 12348 408 13036
rect 350 11992 408 12348
rect 2008 13036 2066 13392
rect 2008 12348 2020 13036
rect 2054 12348 2066 13036
rect 2008 11992 2066 12348
rect 3666 13036 3724 13392
rect 3666 12348 3678 13036
rect 3712 12348 3724 13036
rect 3666 11992 3724 12348
rect 5324 13036 5382 13392
rect 5324 12348 5336 13036
rect 5370 12348 5382 13036
rect 5324 11992 5382 12348
rect 6982 13036 7040 13392
rect 6982 12348 6994 13036
rect 7028 12348 7040 13036
rect 6982 11992 7040 12348
rect 8640 13036 8698 13392
rect 8640 12348 8652 13036
rect 8686 12348 8698 13036
rect 8640 11992 8698 12348
rect 10298 13036 10356 13392
rect 10298 12348 10310 13036
rect 10344 12348 10356 13036
rect 10298 11992 10356 12348
rect 11956 13036 12014 13392
rect 11956 12348 11968 13036
rect 12002 12348 12014 13036
rect 11956 11992 12014 12348
rect 13614 13036 13672 13392
rect 13614 12348 13626 13036
rect 13660 12348 13672 13036
rect 13614 11992 13672 12348
rect 15272 13036 15330 13392
rect 15272 12348 15284 13036
rect 15318 12348 15330 13036
rect 15272 11992 15330 12348
rect 16930 13036 16988 13392
rect 16930 12348 16942 13036
rect 16976 12348 16988 13036
rect 16930 11992 16988 12348
rect 18588 13036 18646 13392
rect 18588 12348 18600 13036
rect 18634 12348 18646 13036
rect 18588 11992 18646 12348
rect 20246 13036 20304 13392
rect 20246 12348 20258 13036
rect 20292 12348 20304 13036
rect 20246 11992 20304 12348
rect 21904 13036 21962 13392
rect 21904 12348 21916 13036
rect 21950 12348 21962 13036
rect 21904 11992 21962 12348
rect 23562 13036 23620 13392
rect 23562 12348 23574 13036
rect 23608 12348 23620 13036
rect 23562 11992 23620 12348
rect 25220 13036 25278 13392
rect 25220 12348 25232 13036
rect 25266 12348 25278 13036
rect 25220 11992 25278 12348
rect 26878 13036 26936 13392
rect 26878 12348 26890 13036
rect 26924 12348 26936 13036
rect 26878 11992 26936 12348
rect 28536 13036 28594 13392
rect 28536 12348 28548 13036
rect 28582 12348 28594 13036
rect 28536 11992 28594 12348
rect 30194 13036 30252 13392
rect 30194 12348 30206 13036
rect 30240 12348 30252 13036
rect 30194 11992 30252 12348
rect 31852 13036 31910 13392
rect 31852 12348 31864 13036
rect 31898 12348 31910 13036
rect 31852 11992 31910 12348
rect 33510 13036 33568 13392
rect 33510 12348 33522 13036
rect 33556 12348 33568 13036
rect 33510 11992 33568 12348
rect -32810 11400 -32752 11756
rect -32810 10712 -32798 11400
rect -32764 10712 -32752 11400
rect -32810 10356 -32752 10712
rect -31152 11400 -31094 11756
rect -31152 10712 -31140 11400
rect -31106 10712 -31094 11400
rect -31152 10356 -31094 10712
rect -29494 11400 -29436 11756
rect -29494 10712 -29482 11400
rect -29448 10712 -29436 11400
rect -29494 10356 -29436 10712
rect -27836 11400 -27778 11756
rect -27836 10712 -27824 11400
rect -27790 10712 -27778 11400
rect -27836 10356 -27778 10712
rect -26178 11400 -26120 11756
rect -26178 10712 -26166 11400
rect -26132 10712 -26120 11400
rect -26178 10356 -26120 10712
rect -24520 11400 -24462 11756
rect -24520 10712 -24508 11400
rect -24474 10712 -24462 11400
rect -24520 10356 -24462 10712
rect -22862 11400 -22804 11756
rect -22862 10712 -22850 11400
rect -22816 10712 -22804 11400
rect -22862 10356 -22804 10712
rect -21204 11400 -21146 11756
rect -21204 10712 -21192 11400
rect -21158 10712 -21146 11400
rect -21204 10356 -21146 10712
rect -19546 11400 -19488 11756
rect -19546 10712 -19534 11400
rect -19500 10712 -19488 11400
rect -19546 10356 -19488 10712
rect -17888 11400 -17830 11756
rect -17888 10712 -17876 11400
rect -17842 10712 -17830 11400
rect -17888 10356 -17830 10712
rect -16230 11400 -16172 11756
rect -16230 10712 -16218 11400
rect -16184 10712 -16172 11400
rect -16230 10356 -16172 10712
rect -14572 11400 -14514 11756
rect -14572 10712 -14560 11400
rect -14526 10712 -14514 11400
rect -14572 10356 -14514 10712
rect -12914 11400 -12856 11756
rect -12914 10712 -12902 11400
rect -12868 10712 -12856 11400
rect -12914 10356 -12856 10712
rect -11256 11400 -11198 11756
rect -11256 10712 -11244 11400
rect -11210 10712 -11198 11400
rect -11256 10356 -11198 10712
rect -9598 11400 -9540 11756
rect -9598 10712 -9586 11400
rect -9552 10712 -9540 11400
rect -9598 10356 -9540 10712
rect -7940 11400 -7882 11756
rect -7940 10712 -7928 11400
rect -7894 10712 -7882 11400
rect -7940 10356 -7882 10712
rect -6282 11400 -6224 11756
rect -6282 10712 -6270 11400
rect -6236 10712 -6224 11400
rect -6282 10356 -6224 10712
rect -4624 11400 -4566 11756
rect -4624 10712 -4612 11400
rect -4578 10712 -4566 11400
rect -4624 10356 -4566 10712
rect -2966 11400 -2908 11756
rect -2966 10712 -2954 11400
rect -2920 10712 -2908 11400
rect -2966 10356 -2908 10712
rect -1308 11400 -1250 11756
rect -1308 10712 -1296 11400
rect -1262 10712 -1250 11400
rect -1308 10356 -1250 10712
rect 350 11400 408 11756
rect 350 10712 362 11400
rect 396 10712 408 11400
rect 350 10356 408 10712
rect 2008 11400 2066 11756
rect 2008 10712 2020 11400
rect 2054 10712 2066 11400
rect 2008 10356 2066 10712
rect 3666 11400 3724 11756
rect 3666 10712 3678 11400
rect 3712 10712 3724 11400
rect 3666 10356 3724 10712
rect 5324 11400 5382 11756
rect 5324 10712 5336 11400
rect 5370 10712 5382 11400
rect 5324 10356 5382 10712
rect 6982 11400 7040 11756
rect 6982 10712 6994 11400
rect 7028 10712 7040 11400
rect 6982 10356 7040 10712
rect 8640 11400 8698 11756
rect 8640 10712 8652 11400
rect 8686 10712 8698 11400
rect 8640 10356 8698 10712
rect 10298 11400 10356 11756
rect 10298 10712 10310 11400
rect 10344 10712 10356 11400
rect 10298 10356 10356 10712
rect 11956 11400 12014 11756
rect 11956 10712 11968 11400
rect 12002 10712 12014 11400
rect 11956 10356 12014 10712
rect 13614 11400 13672 11756
rect 13614 10712 13626 11400
rect 13660 10712 13672 11400
rect 13614 10356 13672 10712
rect 15272 11400 15330 11756
rect 15272 10712 15284 11400
rect 15318 10712 15330 11400
rect 15272 10356 15330 10712
rect 16930 11400 16988 11756
rect 16930 10712 16942 11400
rect 16976 10712 16988 11400
rect 16930 10356 16988 10712
rect 18588 11400 18646 11756
rect 18588 10712 18600 11400
rect 18634 10712 18646 11400
rect 18588 10356 18646 10712
rect 20246 11400 20304 11756
rect 20246 10712 20258 11400
rect 20292 10712 20304 11400
rect 20246 10356 20304 10712
rect 21904 11400 21962 11756
rect 21904 10712 21916 11400
rect 21950 10712 21962 11400
rect 21904 10356 21962 10712
rect 23562 11400 23620 11756
rect 23562 10712 23574 11400
rect 23608 10712 23620 11400
rect 23562 10356 23620 10712
rect 25220 11400 25278 11756
rect 25220 10712 25232 11400
rect 25266 10712 25278 11400
rect 25220 10356 25278 10712
rect 26878 11400 26936 11756
rect 26878 10712 26890 11400
rect 26924 10712 26936 11400
rect 26878 10356 26936 10712
rect 28536 11400 28594 11756
rect 28536 10712 28548 11400
rect 28582 10712 28594 11400
rect 28536 10356 28594 10712
rect 30194 11400 30252 11756
rect 30194 10712 30206 11400
rect 30240 10712 30252 11400
rect 30194 10356 30252 10712
rect 31852 11400 31910 11756
rect 31852 10712 31864 11400
rect 31898 10712 31910 11400
rect 31852 10356 31910 10712
rect 33510 11400 33568 11756
rect 33510 10712 33522 11400
rect 33556 10712 33568 11400
rect 33510 10356 33568 10712
rect -32810 9764 -32752 10120
rect -32810 9076 -32798 9764
rect -32764 9076 -32752 9764
rect -32810 8720 -32752 9076
rect -31152 9764 -31094 10120
rect -31152 9076 -31140 9764
rect -31106 9076 -31094 9764
rect -31152 8720 -31094 9076
rect -29494 9764 -29436 10120
rect -29494 9076 -29482 9764
rect -29448 9076 -29436 9764
rect -29494 8720 -29436 9076
rect -27836 9764 -27778 10120
rect -27836 9076 -27824 9764
rect -27790 9076 -27778 9764
rect -27836 8720 -27778 9076
rect -26178 9764 -26120 10120
rect -26178 9076 -26166 9764
rect -26132 9076 -26120 9764
rect -26178 8720 -26120 9076
rect -24520 9764 -24462 10120
rect -24520 9076 -24508 9764
rect -24474 9076 -24462 9764
rect -24520 8720 -24462 9076
rect -22862 9764 -22804 10120
rect -22862 9076 -22850 9764
rect -22816 9076 -22804 9764
rect -22862 8720 -22804 9076
rect -21204 9764 -21146 10120
rect -21204 9076 -21192 9764
rect -21158 9076 -21146 9764
rect -21204 8720 -21146 9076
rect -19546 9764 -19488 10120
rect -19546 9076 -19534 9764
rect -19500 9076 -19488 9764
rect -19546 8720 -19488 9076
rect -17888 9764 -17830 10120
rect -17888 9076 -17876 9764
rect -17842 9076 -17830 9764
rect -17888 8720 -17830 9076
rect -16230 9764 -16172 10120
rect -16230 9076 -16218 9764
rect -16184 9076 -16172 9764
rect -16230 8720 -16172 9076
rect -14572 9764 -14514 10120
rect -14572 9076 -14560 9764
rect -14526 9076 -14514 9764
rect -14572 8720 -14514 9076
rect -12914 9764 -12856 10120
rect -12914 9076 -12902 9764
rect -12868 9076 -12856 9764
rect -12914 8720 -12856 9076
rect -11256 9764 -11198 10120
rect -11256 9076 -11244 9764
rect -11210 9076 -11198 9764
rect -11256 8720 -11198 9076
rect -9598 9764 -9540 10120
rect -9598 9076 -9586 9764
rect -9552 9076 -9540 9764
rect -9598 8720 -9540 9076
rect -7940 9764 -7882 10120
rect -7940 9076 -7928 9764
rect -7894 9076 -7882 9764
rect -7940 8720 -7882 9076
rect -6282 9764 -6224 10120
rect -6282 9076 -6270 9764
rect -6236 9076 -6224 9764
rect -6282 8720 -6224 9076
rect -4624 9764 -4566 10120
rect -4624 9076 -4612 9764
rect -4578 9076 -4566 9764
rect -4624 8720 -4566 9076
rect -2966 9764 -2908 10120
rect -2966 9076 -2954 9764
rect -2920 9076 -2908 9764
rect -2966 8720 -2908 9076
rect -1308 9764 -1250 10120
rect -1308 9076 -1296 9764
rect -1262 9076 -1250 9764
rect -1308 8720 -1250 9076
rect 350 9764 408 10120
rect 350 9076 362 9764
rect 396 9076 408 9764
rect 350 8720 408 9076
rect 2008 9764 2066 10120
rect 2008 9076 2020 9764
rect 2054 9076 2066 9764
rect 2008 8720 2066 9076
rect 3666 9764 3724 10120
rect 3666 9076 3678 9764
rect 3712 9076 3724 9764
rect 3666 8720 3724 9076
rect 5324 9764 5382 10120
rect 5324 9076 5336 9764
rect 5370 9076 5382 9764
rect 5324 8720 5382 9076
rect 6982 9764 7040 10120
rect 6982 9076 6994 9764
rect 7028 9076 7040 9764
rect 6982 8720 7040 9076
rect 8640 9764 8698 10120
rect 8640 9076 8652 9764
rect 8686 9076 8698 9764
rect 8640 8720 8698 9076
rect 10298 9764 10356 10120
rect 10298 9076 10310 9764
rect 10344 9076 10356 9764
rect 10298 8720 10356 9076
rect 11956 9764 12014 10120
rect 11956 9076 11968 9764
rect 12002 9076 12014 9764
rect 11956 8720 12014 9076
rect 13614 9764 13672 10120
rect 13614 9076 13626 9764
rect 13660 9076 13672 9764
rect 13614 8720 13672 9076
rect 15272 9764 15330 10120
rect 15272 9076 15284 9764
rect 15318 9076 15330 9764
rect 15272 8720 15330 9076
rect 16930 9764 16988 10120
rect 16930 9076 16942 9764
rect 16976 9076 16988 9764
rect 16930 8720 16988 9076
rect 18588 9764 18646 10120
rect 18588 9076 18600 9764
rect 18634 9076 18646 9764
rect 18588 8720 18646 9076
rect 20246 9764 20304 10120
rect 20246 9076 20258 9764
rect 20292 9076 20304 9764
rect 20246 8720 20304 9076
rect 21904 9764 21962 10120
rect 21904 9076 21916 9764
rect 21950 9076 21962 9764
rect 21904 8720 21962 9076
rect 23562 9764 23620 10120
rect 23562 9076 23574 9764
rect 23608 9076 23620 9764
rect 23562 8720 23620 9076
rect 25220 9764 25278 10120
rect 25220 9076 25232 9764
rect 25266 9076 25278 9764
rect 25220 8720 25278 9076
rect 26878 9764 26936 10120
rect 26878 9076 26890 9764
rect 26924 9076 26936 9764
rect 26878 8720 26936 9076
rect 28536 9764 28594 10120
rect 28536 9076 28548 9764
rect 28582 9076 28594 9764
rect 28536 8720 28594 9076
rect 30194 9764 30252 10120
rect 30194 9076 30206 9764
rect 30240 9076 30252 9764
rect 30194 8720 30252 9076
rect 31852 9764 31910 10120
rect 31852 9076 31864 9764
rect 31898 9076 31910 9764
rect 31852 8720 31910 9076
rect 33510 9764 33568 10120
rect 33510 9076 33522 9764
rect 33556 9076 33568 9764
rect 33510 8720 33568 9076
rect -32810 8128 -32752 8484
rect -32810 7440 -32798 8128
rect -32764 7440 -32752 8128
rect -32810 7084 -32752 7440
rect -31152 8128 -31094 8484
rect -31152 7440 -31140 8128
rect -31106 7440 -31094 8128
rect -31152 7084 -31094 7440
rect -29494 8128 -29436 8484
rect -29494 7440 -29482 8128
rect -29448 7440 -29436 8128
rect -29494 7084 -29436 7440
rect -27836 8128 -27778 8484
rect -27836 7440 -27824 8128
rect -27790 7440 -27778 8128
rect -27836 7084 -27778 7440
rect -26178 8128 -26120 8484
rect -26178 7440 -26166 8128
rect -26132 7440 -26120 8128
rect -26178 7084 -26120 7440
rect -24520 8128 -24462 8484
rect -24520 7440 -24508 8128
rect -24474 7440 -24462 8128
rect -24520 7084 -24462 7440
rect -22862 8128 -22804 8484
rect -22862 7440 -22850 8128
rect -22816 7440 -22804 8128
rect -22862 7084 -22804 7440
rect -21204 8128 -21146 8484
rect -21204 7440 -21192 8128
rect -21158 7440 -21146 8128
rect -21204 7084 -21146 7440
rect -19546 8128 -19488 8484
rect -19546 7440 -19534 8128
rect -19500 7440 -19488 8128
rect -19546 7084 -19488 7440
rect -17888 8128 -17830 8484
rect -17888 7440 -17876 8128
rect -17842 7440 -17830 8128
rect -17888 7084 -17830 7440
rect -16230 8128 -16172 8484
rect -16230 7440 -16218 8128
rect -16184 7440 -16172 8128
rect -16230 7084 -16172 7440
rect -14572 8128 -14514 8484
rect -14572 7440 -14560 8128
rect -14526 7440 -14514 8128
rect -14572 7084 -14514 7440
rect -12914 8128 -12856 8484
rect -12914 7440 -12902 8128
rect -12868 7440 -12856 8128
rect -12914 7084 -12856 7440
rect -11256 8128 -11198 8484
rect -11256 7440 -11244 8128
rect -11210 7440 -11198 8128
rect -11256 7084 -11198 7440
rect -9598 8128 -9540 8484
rect -9598 7440 -9586 8128
rect -9552 7440 -9540 8128
rect -9598 7084 -9540 7440
rect -7940 8128 -7882 8484
rect -7940 7440 -7928 8128
rect -7894 7440 -7882 8128
rect -7940 7084 -7882 7440
rect -6282 8128 -6224 8484
rect -6282 7440 -6270 8128
rect -6236 7440 -6224 8128
rect -6282 7084 -6224 7440
rect -4624 8128 -4566 8484
rect -4624 7440 -4612 8128
rect -4578 7440 -4566 8128
rect -4624 7084 -4566 7440
rect -2966 8128 -2908 8484
rect -2966 7440 -2954 8128
rect -2920 7440 -2908 8128
rect -2966 7084 -2908 7440
rect -1308 8128 -1250 8484
rect -1308 7440 -1296 8128
rect -1262 7440 -1250 8128
rect -1308 7084 -1250 7440
rect 350 8128 408 8484
rect 350 7440 362 8128
rect 396 7440 408 8128
rect 350 7084 408 7440
rect 2008 8128 2066 8484
rect 2008 7440 2020 8128
rect 2054 7440 2066 8128
rect 2008 7084 2066 7440
rect 3666 8128 3724 8484
rect 3666 7440 3678 8128
rect 3712 7440 3724 8128
rect 3666 7084 3724 7440
rect 5324 8128 5382 8484
rect 5324 7440 5336 8128
rect 5370 7440 5382 8128
rect 5324 7084 5382 7440
rect 6982 8128 7040 8484
rect 6982 7440 6994 8128
rect 7028 7440 7040 8128
rect 6982 7084 7040 7440
rect 8640 8128 8698 8484
rect 8640 7440 8652 8128
rect 8686 7440 8698 8128
rect 8640 7084 8698 7440
rect 10298 8128 10356 8484
rect 10298 7440 10310 8128
rect 10344 7440 10356 8128
rect 10298 7084 10356 7440
rect 11956 8128 12014 8484
rect 11956 7440 11968 8128
rect 12002 7440 12014 8128
rect 11956 7084 12014 7440
rect 13614 8128 13672 8484
rect 13614 7440 13626 8128
rect 13660 7440 13672 8128
rect 13614 7084 13672 7440
rect 15272 8128 15330 8484
rect 15272 7440 15284 8128
rect 15318 7440 15330 8128
rect 15272 7084 15330 7440
rect 16930 8128 16988 8484
rect 16930 7440 16942 8128
rect 16976 7440 16988 8128
rect 16930 7084 16988 7440
rect 18588 8128 18646 8484
rect 18588 7440 18600 8128
rect 18634 7440 18646 8128
rect 18588 7084 18646 7440
rect 20246 8128 20304 8484
rect 20246 7440 20258 8128
rect 20292 7440 20304 8128
rect 20246 7084 20304 7440
rect 21904 8128 21962 8484
rect 21904 7440 21916 8128
rect 21950 7440 21962 8128
rect 21904 7084 21962 7440
rect 23562 8128 23620 8484
rect 23562 7440 23574 8128
rect 23608 7440 23620 8128
rect 23562 7084 23620 7440
rect 25220 8128 25278 8484
rect 25220 7440 25232 8128
rect 25266 7440 25278 8128
rect 25220 7084 25278 7440
rect 26878 8128 26936 8484
rect 26878 7440 26890 8128
rect 26924 7440 26936 8128
rect 26878 7084 26936 7440
rect 28536 8128 28594 8484
rect 28536 7440 28548 8128
rect 28582 7440 28594 8128
rect 28536 7084 28594 7440
rect 30194 8128 30252 8484
rect 30194 7440 30206 8128
rect 30240 7440 30252 8128
rect 30194 7084 30252 7440
rect 31852 8128 31910 8484
rect 31852 7440 31864 8128
rect 31898 7440 31910 8128
rect 31852 7084 31910 7440
rect 33510 8128 33568 8484
rect 33510 7440 33522 8128
rect 33556 7440 33568 8128
rect 33510 7084 33568 7440
rect -32810 6490 -32752 6846
rect -32810 5802 -32798 6490
rect -32764 5802 -32752 6490
rect -32810 5446 -32752 5802
rect -31152 6490 -31094 6846
rect -31152 5802 -31140 6490
rect -31106 5802 -31094 6490
rect -31152 5446 -31094 5802
rect -29494 6490 -29436 6846
rect -29494 5802 -29482 6490
rect -29448 5802 -29436 6490
rect -29494 5446 -29436 5802
rect -27836 6490 -27778 6846
rect -27836 5802 -27824 6490
rect -27790 5802 -27778 6490
rect -27836 5446 -27778 5802
rect -26178 6490 -26120 6846
rect -26178 5802 -26166 6490
rect -26132 5802 -26120 6490
rect -26178 5446 -26120 5802
rect -24520 6490 -24462 6846
rect -24520 5802 -24508 6490
rect -24474 5802 -24462 6490
rect -24520 5446 -24462 5802
rect -22862 6490 -22804 6846
rect -22862 5802 -22850 6490
rect -22816 5802 -22804 6490
rect -22862 5446 -22804 5802
rect -21204 6490 -21146 6846
rect -21204 5802 -21192 6490
rect -21158 5802 -21146 6490
rect -21204 5446 -21146 5802
rect -19546 6490 -19488 6846
rect -19546 5802 -19534 6490
rect -19500 5802 -19488 6490
rect -19546 5446 -19488 5802
rect -17888 6490 -17830 6846
rect -17888 5802 -17876 6490
rect -17842 5802 -17830 6490
rect -17888 5446 -17830 5802
rect -16230 6490 -16172 6846
rect -16230 5802 -16218 6490
rect -16184 5802 -16172 6490
rect -16230 5446 -16172 5802
rect -14572 6490 -14514 6846
rect -14572 5802 -14560 6490
rect -14526 5802 -14514 6490
rect -14572 5446 -14514 5802
rect -12914 6490 -12856 6846
rect -12914 5802 -12902 6490
rect -12868 5802 -12856 6490
rect -12914 5446 -12856 5802
rect -11256 6490 -11198 6846
rect -11256 5802 -11244 6490
rect -11210 5802 -11198 6490
rect -11256 5446 -11198 5802
rect -9598 6490 -9540 6846
rect -9598 5802 -9586 6490
rect -9552 5802 -9540 6490
rect -9598 5446 -9540 5802
rect -7940 6490 -7882 6846
rect -7940 5802 -7928 6490
rect -7894 5802 -7882 6490
rect -7940 5446 -7882 5802
rect -6282 6490 -6224 6846
rect -6282 5802 -6270 6490
rect -6236 5802 -6224 6490
rect -6282 5446 -6224 5802
rect -4624 6490 -4566 6846
rect -4624 5802 -4612 6490
rect -4578 5802 -4566 6490
rect -4624 5446 -4566 5802
rect -2966 6490 -2908 6846
rect -2966 5802 -2954 6490
rect -2920 5802 -2908 6490
rect -2966 5446 -2908 5802
rect -1308 6490 -1250 6846
rect -1308 5802 -1296 6490
rect -1262 5802 -1250 6490
rect -1308 5446 -1250 5802
rect 350 6490 408 6846
rect 350 5802 362 6490
rect 396 5802 408 6490
rect 350 5446 408 5802
rect 2008 6490 2066 6846
rect 2008 5802 2020 6490
rect 2054 5802 2066 6490
rect 2008 5446 2066 5802
rect 3666 6490 3724 6846
rect 3666 5802 3678 6490
rect 3712 5802 3724 6490
rect 3666 5446 3724 5802
rect 5324 6490 5382 6846
rect 5324 5802 5336 6490
rect 5370 5802 5382 6490
rect 5324 5446 5382 5802
rect 6982 6490 7040 6846
rect 6982 5802 6994 6490
rect 7028 5802 7040 6490
rect 6982 5446 7040 5802
rect 8640 6490 8698 6846
rect 8640 5802 8652 6490
rect 8686 5802 8698 6490
rect 8640 5446 8698 5802
rect 10298 6490 10356 6846
rect 10298 5802 10310 6490
rect 10344 5802 10356 6490
rect 10298 5446 10356 5802
rect 11956 6490 12014 6846
rect 11956 5802 11968 6490
rect 12002 5802 12014 6490
rect 11956 5446 12014 5802
rect 13614 6490 13672 6846
rect 13614 5802 13626 6490
rect 13660 5802 13672 6490
rect 13614 5446 13672 5802
rect 15272 6490 15330 6846
rect 15272 5802 15284 6490
rect 15318 5802 15330 6490
rect 15272 5446 15330 5802
rect 16930 6490 16988 6846
rect 16930 5802 16942 6490
rect 16976 5802 16988 6490
rect 16930 5446 16988 5802
rect 18588 6490 18646 6846
rect 18588 5802 18600 6490
rect 18634 5802 18646 6490
rect 18588 5446 18646 5802
rect 20246 6490 20304 6846
rect 20246 5802 20258 6490
rect 20292 5802 20304 6490
rect 20246 5446 20304 5802
rect 21904 6490 21962 6846
rect 21904 5802 21916 6490
rect 21950 5802 21962 6490
rect 21904 5446 21962 5802
rect 23562 6490 23620 6846
rect 23562 5802 23574 6490
rect 23608 5802 23620 6490
rect 23562 5446 23620 5802
rect 25220 6490 25278 6846
rect 25220 5802 25232 6490
rect 25266 5802 25278 6490
rect 25220 5446 25278 5802
rect 26878 6490 26936 6846
rect 26878 5802 26890 6490
rect 26924 5802 26936 6490
rect 26878 5446 26936 5802
rect 28536 6490 28594 6846
rect 28536 5802 28548 6490
rect 28582 5802 28594 6490
rect 28536 5446 28594 5802
rect 30194 6490 30252 6846
rect 30194 5802 30206 6490
rect 30240 5802 30252 6490
rect 30194 5446 30252 5802
rect 31852 6490 31910 6846
rect 31852 5802 31864 6490
rect 31898 5802 31910 6490
rect 31852 5446 31910 5802
rect 33510 6490 33568 6846
rect 33510 5802 33522 6490
rect 33556 5802 33568 6490
rect 33510 5446 33568 5802
rect -32810 4854 -32752 5210
rect -32810 4166 -32798 4854
rect -32764 4166 -32752 4854
rect -32810 3810 -32752 4166
rect -31152 4854 -31094 5210
rect -31152 4166 -31140 4854
rect -31106 4166 -31094 4854
rect -31152 3810 -31094 4166
rect -29494 4854 -29436 5210
rect -29494 4166 -29482 4854
rect -29448 4166 -29436 4854
rect -29494 3810 -29436 4166
rect -27836 4854 -27778 5210
rect -27836 4166 -27824 4854
rect -27790 4166 -27778 4854
rect -27836 3810 -27778 4166
rect -26178 4854 -26120 5210
rect -26178 4166 -26166 4854
rect -26132 4166 -26120 4854
rect -26178 3810 -26120 4166
rect -24520 4854 -24462 5210
rect -24520 4166 -24508 4854
rect -24474 4166 -24462 4854
rect -24520 3810 -24462 4166
rect -22862 4854 -22804 5210
rect -22862 4166 -22850 4854
rect -22816 4166 -22804 4854
rect -22862 3810 -22804 4166
rect -21204 4854 -21146 5210
rect -21204 4166 -21192 4854
rect -21158 4166 -21146 4854
rect -21204 3810 -21146 4166
rect -19546 4854 -19488 5210
rect -19546 4166 -19534 4854
rect -19500 4166 -19488 4854
rect -19546 3810 -19488 4166
rect -17888 4854 -17830 5210
rect -17888 4166 -17876 4854
rect -17842 4166 -17830 4854
rect -17888 3810 -17830 4166
rect -16230 4854 -16172 5210
rect -16230 4166 -16218 4854
rect -16184 4166 -16172 4854
rect -16230 3810 -16172 4166
rect -14572 4854 -14514 5210
rect -14572 4166 -14560 4854
rect -14526 4166 -14514 4854
rect -14572 3810 -14514 4166
rect -12914 4854 -12856 5210
rect -12914 4166 -12902 4854
rect -12868 4166 -12856 4854
rect -12914 3810 -12856 4166
rect -11256 4854 -11198 5210
rect -11256 4166 -11244 4854
rect -11210 4166 -11198 4854
rect -11256 3810 -11198 4166
rect -9598 4854 -9540 5210
rect -9598 4166 -9586 4854
rect -9552 4166 -9540 4854
rect -9598 3810 -9540 4166
rect -7940 4854 -7882 5210
rect -7940 4166 -7928 4854
rect -7894 4166 -7882 4854
rect -7940 3810 -7882 4166
rect -6282 4854 -6224 5210
rect -6282 4166 -6270 4854
rect -6236 4166 -6224 4854
rect -6282 3810 -6224 4166
rect -4624 4854 -4566 5210
rect -4624 4166 -4612 4854
rect -4578 4166 -4566 4854
rect -4624 3810 -4566 4166
rect -2966 4854 -2908 5210
rect -2966 4166 -2954 4854
rect -2920 4166 -2908 4854
rect -2966 3810 -2908 4166
rect -1308 4854 -1250 5210
rect -1308 4166 -1296 4854
rect -1262 4166 -1250 4854
rect -1308 3810 -1250 4166
rect 350 4854 408 5210
rect 350 4166 362 4854
rect 396 4166 408 4854
rect 350 3810 408 4166
rect 2008 4854 2066 5210
rect 2008 4166 2020 4854
rect 2054 4166 2066 4854
rect 2008 3810 2066 4166
rect 3666 4854 3724 5210
rect 3666 4166 3678 4854
rect 3712 4166 3724 4854
rect 3666 3810 3724 4166
rect 5324 4854 5382 5210
rect 5324 4166 5336 4854
rect 5370 4166 5382 4854
rect 5324 3810 5382 4166
rect 6982 4854 7040 5210
rect 6982 4166 6994 4854
rect 7028 4166 7040 4854
rect 6982 3810 7040 4166
rect 8640 4854 8698 5210
rect 8640 4166 8652 4854
rect 8686 4166 8698 4854
rect 8640 3810 8698 4166
rect 10298 4854 10356 5210
rect 10298 4166 10310 4854
rect 10344 4166 10356 4854
rect 10298 3810 10356 4166
rect 11956 4854 12014 5210
rect 11956 4166 11968 4854
rect 12002 4166 12014 4854
rect 11956 3810 12014 4166
rect 13614 4854 13672 5210
rect 13614 4166 13626 4854
rect 13660 4166 13672 4854
rect 13614 3810 13672 4166
rect 15272 4854 15330 5210
rect 15272 4166 15284 4854
rect 15318 4166 15330 4854
rect 15272 3810 15330 4166
rect 16930 4854 16988 5210
rect 16930 4166 16942 4854
rect 16976 4166 16988 4854
rect 16930 3810 16988 4166
rect 18588 4854 18646 5210
rect 18588 4166 18600 4854
rect 18634 4166 18646 4854
rect 18588 3810 18646 4166
rect 20246 4854 20304 5210
rect 20246 4166 20258 4854
rect 20292 4166 20304 4854
rect 20246 3810 20304 4166
rect 21904 4854 21962 5210
rect 21904 4166 21916 4854
rect 21950 4166 21962 4854
rect 21904 3810 21962 4166
rect 23562 4854 23620 5210
rect 23562 4166 23574 4854
rect 23608 4166 23620 4854
rect 23562 3810 23620 4166
rect 25220 4854 25278 5210
rect 25220 4166 25232 4854
rect 25266 4166 25278 4854
rect 25220 3810 25278 4166
rect 26878 4854 26936 5210
rect 26878 4166 26890 4854
rect 26924 4166 26936 4854
rect 26878 3810 26936 4166
rect 28536 4854 28594 5210
rect 28536 4166 28548 4854
rect 28582 4166 28594 4854
rect 28536 3810 28594 4166
rect 30194 4854 30252 5210
rect 30194 4166 30206 4854
rect 30240 4166 30252 4854
rect 30194 3810 30252 4166
rect 31852 4854 31910 5210
rect 31852 4166 31864 4854
rect 31898 4166 31910 4854
rect 31852 3810 31910 4166
rect 33510 4854 33568 5210
rect 33510 4166 33522 4854
rect 33556 4166 33568 4854
rect 33510 3810 33568 4166
rect -32810 3218 -32752 3574
rect -32810 2530 -32798 3218
rect -32764 2530 -32752 3218
rect -32810 2174 -32752 2530
rect -31152 3218 -31094 3574
rect -31152 2530 -31140 3218
rect -31106 2530 -31094 3218
rect -31152 2174 -31094 2530
rect -29494 3218 -29436 3574
rect -29494 2530 -29482 3218
rect -29448 2530 -29436 3218
rect -29494 2174 -29436 2530
rect -27836 3218 -27778 3574
rect -27836 2530 -27824 3218
rect -27790 2530 -27778 3218
rect -27836 2174 -27778 2530
rect -26178 3218 -26120 3574
rect -26178 2530 -26166 3218
rect -26132 2530 -26120 3218
rect -26178 2174 -26120 2530
rect -24520 3218 -24462 3574
rect -24520 2530 -24508 3218
rect -24474 2530 -24462 3218
rect -24520 2174 -24462 2530
rect -22862 3218 -22804 3574
rect -22862 2530 -22850 3218
rect -22816 2530 -22804 3218
rect -22862 2174 -22804 2530
rect -21204 3218 -21146 3574
rect -21204 2530 -21192 3218
rect -21158 2530 -21146 3218
rect -21204 2174 -21146 2530
rect -19546 3218 -19488 3574
rect -19546 2530 -19534 3218
rect -19500 2530 -19488 3218
rect -19546 2174 -19488 2530
rect -17888 3218 -17830 3574
rect -17888 2530 -17876 3218
rect -17842 2530 -17830 3218
rect -17888 2174 -17830 2530
rect -16230 3218 -16172 3574
rect -16230 2530 -16218 3218
rect -16184 2530 -16172 3218
rect -16230 2174 -16172 2530
rect -14572 3218 -14514 3574
rect -14572 2530 -14560 3218
rect -14526 2530 -14514 3218
rect -14572 2174 -14514 2530
rect -12914 3218 -12856 3574
rect -12914 2530 -12902 3218
rect -12868 2530 -12856 3218
rect -12914 2174 -12856 2530
rect -11256 3218 -11198 3574
rect -11256 2530 -11244 3218
rect -11210 2530 -11198 3218
rect -11256 2174 -11198 2530
rect -9598 3218 -9540 3574
rect -9598 2530 -9586 3218
rect -9552 2530 -9540 3218
rect -9598 2174 -9540 2530
rect -7940 3218 -7882 3574
rect -7940 2530 -7928 3218
rect -7894 2530 -7882 3218
rect -7940 2174 -7882 2530
rect -6282 3218 -6224 3574
rect -6282 2530 -6270 3218
rect -6236 2530 -6224 3218
rect -6282 2174 -6224 2530
rect -4624 3218 -4566 3574
rect -4624 2530 -4612 3218
rect -4578 2530 -4566 3218
rect -4624 2174 -4566 2530
rect -2966 3218 -2908 3574
rect -2966 2530 -2954 3218
rect -2920 2530 -2908 3218
rect -2966 2174 -2908 2530
rect -1308 3218 -1250 3574
rect -1308 2530 -1296 3218
rect -1262 2530 -1250 3218
rect -1308 2174 -1250 2530
rect 350 3218 408 3574
rect 350 2530 362 3218
rect 396 2530 408 3218
rect 350 2174 408 2530
rect 2008 3218 2066 3574
rect 2008 2530 2020 3218
rect 2054 2530 2066 3218
rect 2008 2174 2066 2530
rect 3666 3218 3724 3574
rect 3666 2530 3678 3218
rect 3712 2530 3724 3218
rect 3666 2174 3724 2530
rect 5324 3218 5382 3574
rect 5324 2530 5336 3218
rect 5370 2530 5382 3218
rect 5324 2174 5382 2530
rect 6982 3218 7040 3574
rect 6982 2530 6994 3218
rect 7028 2530 7040 3218
rect 6982 2174 7040 2530
rect 8640 3218 8698 3574
rect 8640 2530 8652 3218
rect 8686 2530 8698 3218
rect 8640 2174 8698 2530
rect 10298 3218 10356 3574
rect 10298 2530 10310 3218
rect 10344 2530 10356 3218
rect 10298 2174 10356 2530
rect 11956 3218 12014 3574
rect 11956 2530 11968 3218
rect 12002 2530 12014 3218
rect 11956 2174 12014 2530
rect 13614 3218 13672 3574
rect 13614 2530 13626 3218
rect 13660 2530 13672 3218
rect 13614 2174 13672 2530
rect 15272 3218 15330 3574
rect 15272 2530 15284 3218
rect 15318 2530 15330 3218
rect 15272 2174 15330 2530
rect 16930 3218 16988 3574
rect 16930 2530 16942 3218
rect 16976 2530 16988 3218
rect 16930 2174 16988 2530
rect 18588 3218 18646 3574
rect 18588 2530 18600 3218
rect 18634 2530 18646 3218
rect 18588 2174 18646 2530
rect 20246 3218 20304 3574
rect 20246 2530 20258 3218
rect 20292 2530 20304 3218
rect 20246 2174 20304 2530
rect 21904 3218 21962 3574
rect 21904 2530 21916 3218
rect 21950 2530 21962 3218
rect 21904 2174 21962 2530
rect 23562 3218 23620 3574
rect 23562 2530 23574 3218
rect 23608 2530 23620 3218
rect 23562 2174 23620 2530
rect 25220 3218 25278 3574
rect 25220 2530 25232 3218
rect 25266 2530 25278 3218
rect 25220 2174 25278 2530
rect 26878 3218 26936 3574
rect 26878 2530 26890 3218
rect 26924 2530 26936 3218
rect 26878 2174 26936 2530
rect 28536 3218 28594 3574
rect 28536 2530 28548 3218
rect 28582 2530 28594 3218
rect 28536 2174 28594 2530
rect 30194 3218 30252 3574
rect 30194 2530 30206 3218
rect 30240 2530 30252 3218
rect 30194 2174 30252 2530
rect 31852 3218 31910 3574
rect 31852 2530 31864 3218
rect 31898 2530 31910 3218
rect 31852 2174 31910 2530
rect 33510 3218 33568 3574
rect 33510 2530 33522 3218
rect 33556 2530 33568 3218
rect 33510 2174 33568 2530
rect -32810 1582 -32752 1938
rect -32810 894 -32798 1582
rect -32764 894 -32752 1582
rect -32810 538 -32752 894
rect -31152 1582 -31094 1938
rect -31152 894 -31140 1582
rect -31106 894 -31094 1582
rect -31152 538 -31094 894
rect -29494 1582 -29436 1938
rect -29494 894 -29482 1582
rect -29448 894 -29436 1582
rect -29494 538 -29436 894
rect -27836 1582 -27778 1938
rect -27836 894 -27824 1582
rect -27790 894 -27778 1582
rect -27836 538 -27778 894
rect -26178 1582 -26120 1938
rect -26178 894 -26166 1582
rect -26132 894 -26120 1582
rect -26178 538 -26120 894
rect -24520 1582 -24462 1938
rect -24520 894 -24508 1582
rect -24474 894 -24462 1582
rect -24520 538 -24462 894
rect -22862 1582 -22804 1938
rect -22862 894 -22850 1582
rect -22816 894 -22804 1582
rect -22862 538 -22804 894
rect -21204 1582 -21146 1938
rect -21204 894 -21192 1582
rect -21158 894 -21146 1582
rect -21204 538 -21146 894
rect -19546 1582 -19488 1938
rect -19546 894 -19534 1582
rect -19500 894 -19488 1582
rect -19546 538 -19488 894
rect -17888 1582 -17830 1938
rect -17888 894 -17876 1582
rect -17842 894 -17830 1582
rect -17888 538 -17830 894
rect -16230 1582 -16172 1938
rect -16230 894 -16218 1582
rect -16184 894 -16172 1582
rect -16230 538 -16172 894
rect -14572 1582 -14514 1938
rect -14572 894 -14560 1582
rect -14526 894 -14514 1582
rect -14572 538 -14514 894
rect -12914 1582 -12856 1938
rect -12914 894 -12902 1582
rect -12868 894 -12856 1582
rect -12914 538 -12856 894
rect -11256 1582 -11198 1938
rect -11256 894 -11244 1582
rect -11210 894 -11198 1582
rect -11256 538 -11198 894
rect -9598 1582 -9540 1938
rect -9598 894 -9586 1582
rect -9552 894 -9540 1582
rect -9598 538 -9540 894
rect -7940 1582 -7882 1938
rect -7940 894 -7928 1582
rect -7894 894 -7882 1582
rect -7940 538 -7882 894
rect -6282 1582 -6224 1938
rect -6282 894 -6270 1582
rect -6236 894 -6224 1582
rect -6282 538 -6224 894
rect -4624 1582 -4566 1938
rect -4624 894 -4612 1582
rect -4578 894 -4566 1582
rect -4624 538 -4566 894
rect -2966 1582 -2908 1938
rect -2966 894 -2954 1582
rect -2920 894 -2908 1582
rect -2966 538 -2908 894
rect -1308 1582 -1250 1938
rect -1308 894 -1296 1582
rect -1262 894 -1250 1582
rect -1308 538 -1250 894
rect 350 1582 408 1938
rect 350 894 362 1582
rect 396 894 408 1582
rect 350 538 408 894
rect 2008 1582 2066 1938
rect 2008 894 2020 1582
rect 2054 894 2066 1582
rect 2008 538 2066 894
rect 3666 1582 3724 1938
rect 3666 894 3678 1582
rect 3712 894 3724 1582
rect 3666 538 3724 894
rect 5324 1582 5382 1938
rect 5324 894 5336 1582
rect 5370 894 5382 1582
rect 5324 538 5382 894
rect 6982 1582 7040 1938
rect 6982 894 6994 1582
rect 7028 894 7040 1582
rect 6982 538 7040 894
rect 8640 1582 8698 1938
rect 8640 894 8652 1582
rect 8686 894 8698 1582
rect 8640 538 8698 894
rect 10298 1582 10356 1938
rect 10298 894 10310 1582
rect 10344 894 10356 1582
rect 10298 538 10356 894
rect 11956 1582 12014 1938
rect 11956 894 11968 1582
rect 12002 894 12014 1582
rect 11956 538 12014 894
rect 13614 1582 13672 1938
rect 13614 894 13626 1582
rect 13660 894 13672 1582
rect 13614 538 13672 894
rect 15272 1582 15330 1938
rect 15272 894 15284 1582
rect 15318 894 15330 1582
rect 15272 538 15330 894
rect 16930 1582 16988 1938
rect 16930 894 16942 1582
rect 16976 894 16988 1582
rect 16930 538 16988 894
rect 18588 1582 18646 1938
rect 18588 894 18600 1582
rect 18634 894 18646 1582
rect 18588 538 18646 894
rect 20246 1582 20304 1938
rect 20246 894 20258 1582
rect 20292 894 20304 1582
rect 20246 538 20304 894
rect 21904 1582 21962 1938
rect 21904 894 21916 1582
rect 21950 894 21962 1582
rect 21904 538 21962 894
rect 23562 1582 23620 1938
rect 23562 894 23574 1582
rect 23608 894 23620 1582
rect 23562 538 23620 894
rect 25220 1582 25278 1938
rect 25220 894 25232 1582
rect 25266 894 25278 1582
rect 25220 538 25278 894
rect 26878 1582 26936 1938
rect 26878 894 26890 1582
rect 26924 894 26936 1582
rect 26878 538 26936 894
rect 28536 1582 28594 1938
rect 28536 894 28548 1582
rect 28582 894 28594 1582
rect 28536 538 28594 894
rect 30194 1582 30252 1938
rect 30194 894 30206 1582
rect 30240 894 30252 1582
rect 30194 538 30252 894
rect 31852 1582 31910 1938
rect 31852 894 31864 1582
rect 31898 894 31910 1582
rect 31852 538 31910 894
rect 33510 1582 33568 1938
rect 33510 894 33522 1582
rect 33556 894 33568 1582
rect 33510 538 33568 894
rect 32 2 90 96
rect 28 -10 90 2
rect 28 -198 40 -10
rect 74 -198 90 -10
rect 28 -210 90 -198
rect 32 -304 90 -210
rect 120 -10 186 96
rect 120 -198 136 -10
rect 170 -198 186 -10
rect 120 -304 186 -198
rect 216 -10 282 96
rect 216 -198 232 -10
rect 266 -198 282 -10
rect 216 -304 282 -198
rect 312 -10 378 96
rect 312 -198 328 -10
rect 362 -198 378 -10
rect 312 -304 378 -198
rect 408 2 466 96
rect 408 -10 470 2
rect 408 -198 424 -10
rect 458 -198 470 -10
rect 408 -210 470 -198
rect 408 -304 466 -210
<< ndiffc >>
rect -8 -692 26 -604
rect 88 -692 122 -604
rect 184 -692 218 -604
rect 280 -692 314 -604
rect 376 -692 410 -604
<< pdiffc >>
rect -32800 15730 -32766 16418
rect -31142 15730 -31108 16418
rect -29484 15730 -29450 16418
rect -27826 15730 -27792 16418
rect -26168 15730 -26134 16418
rect -24510 15730 -24476 16418
rect -22852 15730 -22818 16418
rect -21194 15730 -21160 16418
rect -19536 15730 -19502 16418
rect -17878 15730 -17844 16418
rect -16220 15730 -16186 16418
rect -14562 15730 -14528 16418
rect -12904 15730 -12870 16418
rect -11246 15730 -11212 16418
rect -9588 15730 -9554 16418
rect -7930 15730 -7896 16418
rect -6272 15730 -6238 16418
rect -4614 15730 -4580 16418
rect -2956 15730 -2922 16418
rect -1298 15730 -1264 16418
rect 360 15730 394 16418
rect 2018 15730 2052 16418
rect 3676 15730 3710 16418
rect 5334 15730 5368 16418
rect 6992 15730 7026 16418
rect 8650 15730 8684 16418
rect 10308 15730 10342 16418
rect 11966 15730 12000 16418
rect 13624 15730 13658 16418
rect 15282 15730 15316 16418
rect 16940 15730 16974 16418
rect 18598 15730 18632 16418
rect 20256 15730 20290 16418
rect 21914 15730 21948 16418
rect 23572 15730 23606 16418
rect 25230 15730 25264 16418
rect 26888 15730 26922 16418
rect 28546 15730 28580 16418
rect 30204 15730 30238 16418
rect 31862 15730 31896 16418
rect 33520 15730 33554 16418
rect -32800 14094 -32766 14782
rect -31142 14094 -31108 14782
rect -29484 14094 -29450 14782
rect -27826 14094 -27792 14782
rect -26168 14094 -26134 14782
rect -24510 14094 -24476 14782
rect -22852 14094 -22818 14782
rect -21194 14094 -21160 14782
rect -19536 14094 -19502 14782
rect -17878 14094 -17844 14782
rect -16220 14094 -16186 14782
rect -14562 14094 -14528 14782
rect -12904 14094 -12870 14782
rect -11246 14094 -11212 14782
rect -9588 14094 -9554 14782
rect -7930 14094 -7896 14782
rect -6272 14094 -6238 14782
rect -4614 14094 -4580 14782
rect -2956 14094 -2922 14782
rect -1298 14094 -1264 14782
rect 360 14094 394 14782
rect 2018 14094 2052 14782
rect 3676 14094 3710 14782
rect 5334 14094 5368 14782
rect 6992 14094 7026 14782
rect 8650 14094 8684 14782
rect 10308 14094 10342 14782
rect 11966 14094 12000 14782
rect 13624 14094 13658 14782
rect 15282 14094 15316 14782
rect 16940 14094 16974 14782
rect 18598 14094 18632 14782
rect 20256 14094 20290 14782
rect 21914 14094 21948 14782
rect 23572 14094 23606 14782
rect 25230 14094 25264 14782
rect 26888 14094 26922 14782
rect 28546 14094 28580 14782
rect 30204 14094 30238 14782
rect 31862 14094 31896 14782
rect 33520 14094 33554 14782
rect -32798 12348 -32764 13036
rect -31140 12348 -31106 13036
rect -29482 12348 -29448 13036
rect -27824 12348 -27790 13036
rect -26166 12348 -26132 13036
rect -24508 12348 -24474 13036
rect -22850 12348 -22816 13036
rect -21192 12348 -21158 13036
rect -19534 12348 -19500 13036
rect -17876 12348 -17842 13036
rect -16218 12348 -16184 13036
rect -14560 12348 -14526 13036
rect -12902 12348 -12868 13036
rect -11244 12348 -11210 13036
rect -9586 12348 -9552 13036
rect -7928 12348 -7894 13036
rect -6270 12348 -6236 13036
rect -4612 12348 -4578 13036
rect -2954 12348 -2920 13036
rect -1296 12348 -1262 13036
rect 362 12348 396 13036
rect 2020 12348 2054 13036
rect 3678 12348 3712 13036
rect 5336 12348 5370 13036
rect 6994 12348 7028 13036
rect 8652 12348 8686 13036
rect 10310 12348 10344 13036
rect 11968 12348 12002 13036
rect 13626 12348 13660 13036
rect 15284 12348 15318 13036
rect 16942 12348 16976 13036
rect 18600 12348 18634 13036
rect 20258 12348 20292 13036
rect 21916 12348 21950 13036
rect 23574 12348 23608 13036
rect 25232 12348 25266 13036
rect 26890 12348 26924 13036
rect 28548 12348 28582 13036
rect 30206 12348 30240 13036
rect 31864 12348 31898 13036
rect 33522 12348 33556 13036
rect -32798 10712 -32764 11400
rect -31140 10712 -31106 11400
rect -29482 10712 -29448 11400
rect -27824 10712 -27790 11400
rect -26166 10712 -26132 11400
rect -24508 10712 -24474 11400
rect -22850 10712 -22816 11400
rect -21192 10712 -21158 11400
rect -19534 10712 -19500 11400
rect -17876 10712 -17842 11400
rect -16218 10712 -16184 11400
rect -14560 10712 -14526 11400
rect -12902 10712 -12868 11400
rect -11244 10712 -11210 11400
rect -9586 10712 -9552 11400
rect -7928 10712 -7894 11400
rect -6270 10712 -6236 11400
rect -4612 10712 -4578 11400
rect -2954 10712 -2920 11400
rect -1296 10712 -1262 11400
rect 362 10712 396 11400
rect 2020 10712 2054 11400
rect 3678 10712 3712 11400
rect 5336 10712 5370 11400
rect 6994 10712 7028 11400
rect 8652 10712 8686 11400
rect 10310 10712 10344 11400
rect 11968 10712 12002 11400
rect 13626 10712 13660 11400
rect 15284 10712 15318 11400
rect 16942 10712 16976 11400
rect 18600 10712 18634 11400
rect 20258 10712 20292 11400
rect 21916 10712 21950 11400
rect 23574 10712 23608 11400
rect 25232 10712 25266 11400
rect 26890 10712 26924 11400
rect 28548 10712 28582 11400
rect 30206 10712 30240 11400
rect 31864 10712 31898 11400
rect 33522 10712 33556 11400
rect -32798 9076 -32764 9764
rect -31140 9076 -31106 9764
rect -29482 9076 -29448 9764
rect -27824 9076 -27790 9764
rect -26166 9076 -26132 9764
rect -24508 9076 -24474 9764
rect -22850 9076 -22816 9764
rect -21192 9076 -21158 9764
rect -19534 9076 -19500 9764
rect -17876 9076 -17842 9764
rect -16218 9076 -16184 9764
rect -14560 9076 -14526 9764
rect -12902 9076 -12868 9764
rect -11244 9076 -11210 9764
rect -9586 9076 -9552 9764
rect -7928 9076 -7894 9764
rect -6270 9076 -6236 9764
rect -4612 9076 -4578 9764
rect -2954 9076 -2920 9764
rect -1296 9076 -1262 9764
rect 362 9076 396 9764
rect 2020 9076 2054 9764
rect 3678 9076 3712 9764
rect 5336 9076 5370 9764
rect 6994 9076 7028 9764
rect 8652 9076 8686 9764
rect 10310 9076 10344 9764
rect 11968 9076 12002 9764
rect 13626 9076 13660 9764
rect 15284 9076 15318 9764
rect 16942 9076 16976 9764
rect 18600 9076 18634 9764
rect 20258 9076 20292 9764
rect 21916 9076 21950 9764
rect 23574 9076 23608 9764
rect 25232 9076 25266 9764
rect 26890 9076 26924 9764
rect 28548 9076 28582 9764
rect 30206 9076 30240 9764
rect 31864 9076 31898 9764
rect 33522 9076 33556 9764
rect -32798 7440 -32764 8128
rect -31140 7440 -31106 8128
rect -29482 7440 -29448 8128
rect -27824 7440 -27790 8128
rect -26166 7440 -26132 8128
rect -24508 7440 -24474 8128
rect -22850 7440 -22816 8128
rect -21192 7440 -21158 8128
rect -19534 7440 -19500 8128
rect -17876 7440 -17842 8128
rect -16218 7440 -16184 8128
rect -14560 7440 -14526 8128
rect -12902 7440 -12868 8128
rect -11244 7440 -11210 8128
rect -9586 7440 -9552 8128
rect -7928 7440 -7894 8128
rect -6270 7440 -6236 8128
rect -4612 7440 -4578 8128
rect -2954 7440 -2920 8128
rect -1296 7440 -1262 8128
rect 362 7440 396 8128
rect 2020 7440 2054 8128
rect 3678 7440 3712 8128
rect 5336 7440 5370 8128
rect 6994 7440 7028 8128
rect 8652 7440 8686 8128
rect 10310 7440 10344 8128
rect 11968 7440 12002 8128
rect 13626 7440 13660 8128
rect 15284 7440 15318 8128
rect 16942 7440 16976 8128
rect 18600 7440 18634 8128
rect 20258 7440 20292 8128
rect 21916 7440 21950 8128
rect 23574 7440 23608 8128
rect 25232 7440 25266 8128
rect 26890 7440 26924 8128
rect 28548 7440 28582 8128
rect 30206 7440 30240 8128
rect 31864 7440 31898 8128
rect 33522 7440 33556 8128
rect -32798 5802 -32764 6490
rect -31140 5802 -31106 6490
rect -29482 5802 -29448 6490
rect -27824 5802 -27790 6490
rect -26166 5802 -26132 6490
rect -24508 5802 -24474 6490
rect -22850 5802 -22816 6490
rect -21192 5802 -21158 6490
rect -19534 5802 -19500 6490
rect -17876 5802 -17842 6490
rect -16218 5802 -16184 6490
rect -14560 5802 -14526 6490
rect -12902 5802 -12868 6490
rect -11244 5802 -11210 6490
rect -9586 5802 -9552 6490
rect -7928 5802 -7894 6490
rect -6270 5802 -6236 6490
rect -4612 5802 -4578 6490
rect -2954 5802 -2920 6490
rect -1296 5802 -1262 6490
rect 362 5802 396 6490
rect 2020 5802 2054 6490
rect 3678 5802 3712 6490
rect 5336 5802 5370 6490
rect 6994 5802 7028 6490
rect 8652 5802 8686 6490
rect 10310 5802 10344 6490
rect 11968 5802 12002 6490
rect 13626 5802 13660 6490
rect 15284 5802 15318 6490
rect 16942 5802 16976 6490
rect 18600 5802 18634 6490
rect 20258 5802 20292 6490
rect 21916 5802 21950 6490
rect 23574 5802 23608 6490
rect 25232 5802 25266 6490
rect 26890 5802 26924 6490
rect 28548 5802 28582 6490
rect 30206 5802 30240 6490
rect 31864 5802 31898 6490
rect 33522 5802 33556 6490
rect -32798 4166 -32764 4854
rect -31140 4166 -31106 4854
rect -29482 4166 -29448 4854
rect -27824 4166 -27790 4854
rect -26166 4166 -26132 4854
rect -24508 4166 -24474 4854
rect -22850 4166 -22816 4854
rect -21192 4166 -21158 4854
rect -19534 4166 -19500 4854
rect -17876 4166 -17842 4854
rect -16218 4166 -16184 4854
rect -14560 4166 -14526 4854
rect -12902 4166 -12868 4854
rect -11244 4166 -11210 4854
rect -9586 4166 -9552 4854
rect -7928 4166 -7894 4854
rect -6270 4166 -6236 4854
rect -4612 4166 -4578 4854
rect -2954 4166 -2920 4854
rect -1296 4166 -1262 4854
rect 362 4166 396 4854
rect 2020 4166 2054 4854
rect 3678 4166 3712 4854
rect 5336 4166 5370 4854
rect 6994 4166 7028 4854
rect 8652 4166 8686 4854
rect 10310 4166 10344 4854
rect 11968 4166 12002 4854
rect 13626 4166 13660 4854
rect 15284 4166 15318 4854
rect 16942 4166 16976 4854
rect 18600 4166 18634 4854
rect 20258 4166 20292 4854
rect 21916 4166 21950 4854
rect 23574 4166 23608 4854
rect 25232 4166 25266 4854
rect 26890 4166 26924 4854
rect 28548 4166 28582 4854
rect 30206 4166 30240 4854
rect 31864 4166 31898 4854
rect 33522 4166 33556 4854
rect -32798 2530 -32764 3218
rect -31140 2530 -31106 3218
rect -29482 2530 -29448 3218
rect -27824 2530 -27790 3218
rect -26166 2530 -26132 3218
rect -24508 2530 -24474 3218
rect -22850 2530 -22816 3218
rect -21192 2530 -21158 3218
rect -19534 2530 -19500 3218
rect -17876 2530 -17842 3218
rect -16218 2530 -16184 3218
rect -14560 2530 -14526 3218
rect -12902 2530 -12868 3218
rect -11244 2530 -11210 3218
rect -9586 2530 -9552 3218
rect -7928 2530 -7894 3218
rect -6270 2530 -6236 3218
rect -4612 2530 -4578 3218
rect -2954 2530 -2920 3218
rect -1296 2530 -1262 3218
rect 362 2530 396 3218
rect 2020 2530 2054 3218
rect 3678 2530 3712 3218
rect 5336 2530 5370 3218
rect 6994 2530 7028 3218
rect 8652 2530 8686 3218
rect 10310 2530 10344 3218
rect 11968 2530 12002 3218
rect 13626 2530 13660 3218
rect 15284 2530 15318 3218
rect 16942 2530 16976 3218
rect 18600 2530 18634 3218
rect 20258 2530 20292 3218
rect 21916 2530 21950 3218
rect 23574 2530 23608 3218
rect 25232 2530 25266 3218
rect 26890 2530 26924 3218
rect 28548 2530 28582 3218
rect 30206 2530 30240 3218
rect 31864 2530 31898 3218
rect 33522 2530 33556 3218
rect -32798 894 -32764 1582
rect -31140 894 -31106 1582
rect -29482 894 -29448 1582
rect -27824 894 -27790 1582
rect -26166 894 -26132 1582
rect -24508 894 -24474 1582
rect -22850 894 -22816 1582
rect -21192 894 -21158 1582
rect -19534 894 -19500 1582
rect -17876 894 -17842 1582
rect -16218 894 -16184 1582
rect -14560 894 -14526 1582
rect -12902 894 -12868 1582
rect -11244 894 -11210 1582
rect -9586 894 -9552 1582
rect -7928 894 -7894 1582
rect -6270 894 -6236 1582
rect -4612 894 -4578 1582
rect -2954 894 -2920 1582
rect -1296 894 -1262 1582
rect 362 894 396 1582
rect 2020 894 2054 1582
rect 3678 894 3712 1582
rect 5336 894 5370 1582
rect 6994 894 7028 1582
rect 8652 894 8686 1582
rect 10310 894 10344 1582
rect 11968 894 12002 1582
rect 13626 894 13660 1582
rect 15284 894 15318 1582
rect 16942 894 16976 1582
rect 18600 894 18634 1582
rect 20258 894 20292 1582
rect 21916 894 21950 1582
rect 23574 894 23608 1582
rect 25232 894 25266 1582
rect 26890 894 26924 1582
rect 28548 894 28582 1582
rect 30206 894 30240 1582
rect 31864 894 31898 1582
rect 33522 894 33556 1582
rect 40 -198 74 -10
rect 136 -198 170 -10
rect 232 -198 266 -10
rect 328 -198 362 -10
rect 424 -198 458 -10
<< psubdiff >>
rect -86 -916 518 -900
rect -86 -968 -54 -916
rect 4 -968 346 -916
rect 404 -968 518 -916
rect -86 -982 518 -968
<< nsubdiff >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect 33976 13946 35004 15480
rect -34456 11946 -33510 13480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect 33976 11946 35004 13480
rect -34456 9946 -33510 11480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect 33976 3946 35004 5480
rect -34456 1946 -33510 3480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect 33976 1946 35004 3480
rect -34456 388 -33510 1480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect 33976 52 35004 1480
rect 1532 -54 35054 52
rect -34586 -828 -734 -520
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
<< psubdiffcont >>
rect -54 -968 4 -916
rect 346 -968 404 -916
<< nsubdiffcont >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect 34166 15480 34698 15946
rect -34234 13480 -33702 13946
rect 34166 13480 34698 13946
rect -34234 11480 -33702 11946
rect 34166 11480 34698 11946
rect -34234 9480 -33702 9946
rect 34166 9480 34698 9946
rect -34234 7480 -33702 7946
rect 34166 7480 34698 7946
rect -34234 5480 -33702 5946
rect 34166 5480 34698 5946
rect -34234 3480 -33702 3946
rect 34166 3480 34698 3946
rect -34234 1480 -33702 1946
rect 34166 1480 34698 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
<< poly >>
rect -32362 16855 -31546 16871
rect -32362 16838 -32346 16855
rect -32754 16821 -32346 16838
rect -31562 16838 -31546 16855
rect -30704 16855 -29888 16871
rect -30704 16838 -30688 16855
rect -31562 16821 -31154 16838
rect -32754 16774 -31154 16821
rect -31096 16821 -30688 16838
rect -29904 16838 -29888 16855
rect -29046 16855 -28230 16871
rect -29046 16838 -29030 16855
rect -29904 16821 -29496 16838
rect -31096 16774 -29496 16821
rect -29438 16821 -29030 16838
rect -28246 16838 -28230 16855
rect -27388 16855 -26572 16871
rect -27388 16838 -27372 16855
rect -28246 16821 -27838 16838
rect -29438 16774 -27838 16821
rect -27780 16821 -27372 16838
rect -26588 16838 -26572 16855
rect -25730 16855 -24914 16871
rect -25730 16838 -25714 16855
rect -26588 16821 -26180 16838
rect -27780 16774 -26180 16821
rect -26122 16821 -25714 16838
rect -24930 16838 -24914 16855
rect -24072 16855 -23256 16871
rect -24072 16838 -24056 16855
rect -24930 16821 -24522 16838
rect -26122 16774 -24522 16821
rect -24464 16821 -24056 16838
rect -23272 16838 -23256 16855
rect -22414 16855 -21598 16871
rect -22414 16838 -22398 16855
rect -23272 16821 -22864 16838
rect -24464 16774 -22864 16821
rect -22806 16821 -22398 16838
rect -21614 16838 -21598 16855
rect -20756 16855 -19940 16871
rect -20756 16838 -20740 16855
rect -21614 16821 -21206 16838
rect -22806 16774 -21206 16821
rect -21148 16821 -20740 16838
rect -19956 16838 -19940 16855
rect -19098 16855 -18282 16871
rect -19098 16838 -19082 16855
rect -19956 16821 -19548 16838
rect -21148 16774 -19548 16821
rect -19490 16821 -19082 16838
rect -18298 16838 -18282 16855
rect -17440 16855 -16624 16871
rect -17440 16838 -17424 16855
rect -18298 16821 -17890 16838
rect -19490 16774 -17890 16821
rect -17832 16821 -17424 16838
rect -16640 16838 -16624 16855
rect -15782 16855 -14966 16871
rect -15782 16838 -15766 16855
rect -16640 16821 -16232 16838
rect -17832 16774 -16232 16821
rect -16174 16821 -15766 16838
rect -14982 16838 -14966 16855
rect -14124 16855 -13308 16871
rect -14124 16838 -14108 16855
rect -14982 16821 -14574 16838
rect -16174 16774 -14574 16821
rect -14516 16821 -14108 16838
rect -13324 16838 -13308 16855
rect -12466 16855 -11650 16871
rect -12466 16838 -12450 16855
rect -13324 16821 -12916 16838
rect -14516 16774 -12916 16821
rect -12858 16821 -12450 16838
rect -11666 16838 -11650 16855
rect -10808 16855 -9992 16871
rect -10808 16838 -10792 16855
rect -11666 16821 -11258 16838
rect -12858 16774 -11258 16821
rect -11200 16821 -10792 16838
rect -10008 16838 -9992 16855
rect -9150 16855 -8334 16871
rect -9150 16838 -9134 16855
rect -10008 16821 -9600 16838
rect -11200 16774 -9600 16821
rect -9542 16821 -9134 16838
rect -8350 16838 -8334 16855
rect -7492 16855 -6676 16871
rect -7492 16838 -7476 16855
rect -8350 16821 -7942 16838
rect -9542 16774 -7942 16821
rect -7884 16821 -7476 16838
rect -6692 16838 -6676 16855
rect -5834 16855 -5018 16871
rect -5834 16838 -5818 16855
rect -6692 16821 -6284 16838
rect -7884 16774 -6284 16821
rect -6226 16821 -5818 16838
rect -5034 16838 -5018 16855
rect -4176 16855 -3360 16871
rect -4176 16838 -4160 16855
rect -5034 16821 -4626 16838
rect -6226 16774 -4626 16821
rect -4568 16821 -4160 16838
rect -3376 16838 -3360 16855
rect -2518 16855 -1702 16871
rect -2518 16838 -2502 16855
rect -3376 16821 -2968 16838
rect -4568 16774 -2968 16821
rect -2910 16821 -2502 16838
rect -1718 16838 -1702 16855
rect -860 16855 -44 16871
rect -860 16838 -844 16855
rect -1718 16821 -1310 16838
rect -2910 16774 -1310 16821
rect -1252 16821 -844 16838
rect -60 16838 -44 16855
rect 798 16855 1614 16871
rect 798 16838 814 16855
rect -60 16821 348 16838
rect -1252 16774 348 16821
rect 406 16821 814 16838
rect 1598 16838 1614 16855
rect 2456 16855 3272 16871
rect 2456 16838 2472 16855
rect 1598 16821 2006 16838
rect 406 16774 2006 16821
rect 2064 16821 2472 16838
rect 3256 16838 3272 16855
rect 4114 16855 4930 16871
rect 4114 16838 4130 16855
rect 3256 16821 3664 16838
rect 2064 16774 3664 16821
rect 3722 16821 4130 16838
rect 4914 16838 4930 16855
rect 5772 16855 6588 16871
rect 5772 16838 5788 16855
rect 4914 16821 5322 16838
rect 3722 16774 5322 16821
rect 5380 16821 5788 16838
rect 6572 16838 6588 16855
rect 7430 16855 8246 16871
rect 7430 16838 7446 16855
rect 6572 16821 6980 16838
rect 5380 16774 6980 16821
rect 7038 16821 7446 16838
rect 8230 16838 8246 16855
rect 9088 16855 9904 16871
rect 9088 16838 9104 16855
rect 8230 16821 8638 16838
rect 7038 16774 8638 16821
rect 8696 16821 9104 16838
rect 9888 16838 9904 16855
rect 10746 16855 11562 16871
rect 10746 16838 10762 16855
rect 9888 16821 10296 16838
rect 8696 16774 10296 16821
rect 10354 16821 10762 16838
rect 11546 16838 11562 16855
rect 12404 16855 13220 16871
rect 12404 16838 12420 16855
rect 11546 16821 11954 16838
rect 10354 16774 11954 16821
rect 12012 16821 12420 16838
rect 13204 16838 13220 16855
rect 14062 16855 14878 16871
rect 14062 16838 14078 16855
rect 13204 16821 13612 16838
rect 12012 16774 13612 16821
rect 13670 16821 14078 16838
rect 14862 16838 14878 16855
rect 15720 16855 16536 16871
rect 15720 16838 15736 16855
rect 14862 16821 15270 16838
rect 13670 16774 15270 16821
rect 15328 16821 15736 16838
rect 16520 16838 16536 16855
rect 17378 16855 18194 16871
rect 17378 16838 17394 16855
rect 16520 16821 16928 16838
rect 15328 16774 16928 16821
rect 16986 16821 17394 16838
rect 18178 16838 18194 16855
rect 19036 16855 19852 16871
rect 19036 16838 19052 16855
rect 18178 16821 18586 16838
rect 16986 16774 18586 16821
rect 18644 16821 19052 16838
rect 19836 16838 19852 16855
rect 20694 16855 21510 16871
rect 20694 16838 20710 16855
rect 19836 16821 20244 16838
rect 18644 16774 20244 16821
rect 20302 16821 20710 16838
rect 21494 16838 21510 16855
rect 22352 16855 23168 16871
rect 22352 16838 22368 16855
rect 21494 16821 21902 16838
rect 20302 16774 21902 16821
rect 21960 16821 22368 16838
rect 23152 16838 23168 16855
rect 24010 16855 24826 16871
rect 24010 16838 24026 16855
rect 23152 16821 23560 16838
rect 21960 16774 23560 16821
rect 23618 16821 24026 16838
rect 24810 16838 24826 16855
rect 25668 16855 26484 16871
rect 25668 16838 25684 16855
rect 24810 16821 25218 16838
rect 23618 16774 25218 16821
rect 25276 16821 25684 16838
rect 26468 16838 26484 16855
rect 27326 16855 28142 16871
rect 27326 16838 27342 16855
rect 26468 16821 26876 16838
rect 25276 16774 26876 16821
rect 26934 16821 27342 16838
rect 28126 16838 28142 16855
rect 28984 16855 29800 16871
rect 28984 16838 29000 16855
rect 28126 16821 28534 16838
rect 26934 16774 28534 16821
rect 28592 16821 29000 16838
rect 29784 16838 29800 16855
rect 30642 16855 31458 16871
rect 30642 16838 30658 16855
rect 29784 16821 30192 16838
rect 28592 16774 30192 16821
rect 30250 16821 30658 16838
rect 31442 16838 31458 16855
rect 32300 16855 33116 16871
rect 32300 16838 32316 16855
rect 31442 16821 31850 16838
rect 30250 16774 31850 16821
rect 31908 16821 32316 16838
rect 33100 16838 33116 16855
rect 33100 16821 33508 16838
rect 31908 16774 33508 16821
rect -32754 15327 -31154 15374
rect -32754 15310 -32346 15327
rect -32362 15293 -32346 15310
rect -31562 15310 -31154 15327
rect -31096 15327 -29496 15374
rect -31096 15310 -30688 15327
rect -31562 15293 -31546 15310
rect -32362 15277 -31546 15293
rect -30704 15293 -30688 15310
rect -29904 15310 -29496 15327
rect -29438 15327 -27838 15374
rect -29438 15310 -29030 15327
rect -29904 15293 -29888 15310
rect -30704 15277 -29888 15293
rect -29046 15293 -29030 15310
rect -28246 15310 -27838 15327
rect -27780 15327 -26180 15374
rect -27780 15310 -27372 15327
rect -28246 15293 -28230 15310
rect -29046 15277 -28230 15293
rect -27388 15293 -27372 15310
rect -26588 15310 -26180 15327
rect -26122 15327 -24522 15374
rect -26122 15310 -25714 15327
rect -26588 15293 -26572 15310
rect -27388 15277 -26572 15293
rect -25730 15293 -25714 15310
rect -24930 15310 -24522 15327
rect -24464 15327 -22864 15374
rect -24464 15310 -24056 15327
rect -24930 15293 -24914 15310
rect -25730 15277 -24914 15293
rect -24072 15293 -24056 15310
rect -23272 15310 -22864 15327
rect -22806 15327 -21206 15374
rect -22806 15310 -22398 15327
rect -23272 15293 -23256 15310
rect -24072 15277 -23256 15293
rect -22414 15293 -22398 15310
rect -21614 15310 -21206 15327
rect -21148 15327 -19548 15374
rect -21148 15310 -20740 15327
rect -21614 15293 -21598 15310
rect -22414 15277 -21598 15293
rect -20756 15293 -20740 15310
rect -19956 15310 -19548 15327
rect -19490 15327 -17890 15374
rect -19490 15310 -19082 15327
rect -19956 15293 -19940 15310
rect -20756 15277 -19940 15293
rect -19098 15293 -19082 15310
rect -18298 15310 -17890 15327
rect -17832 15327 -16232 15374
rect -17832 15310 -17424 15327
rect -18298 15293 -18282 15310
rect -19098 15277 -18282 15293
rect -17440 15293 -17424 15310
rect -16640 15310 -16232 15327
rect -16174 15327 -14574 15374
rect -16174 15310 -15766 15327
rect -16640 15293 -16624 15310
rect -17440 15277 -16624 15293
rect -15782 15293 -15766 15310
rect -14982 15310 -14574 15327
rect -14516 15327 -12916 15374
rect -14516 15310 -14108 15327
rect -14982 15293 -14966 15310
rect -15782 15277 -14966 15293
rect -14124 15293 -14108 15310
rect -13324 15310 -12916 15327
rect -12858 15327 -11258 15374
rect -12858 15310 -12450 15327
rect -13324 15293 -13308 15310
rect -14124 15277 -13308 15293
rect -12466 15293 -12450 15310
rect -11666 15310 -11258 15327
rect -11200 15327 -9600 15374
rect -11200 15310 -10792 15327
rect -11666 15293 -11650 15310
rect -12466 15277 -11650 15293
rect -10808 15293 -10792 15310
rect -10008 15310 -9600 15327
rect -9542 15327 -7942 15374
rect -9542 15310 -9134 15327
rect -10008 15293 -9992 15310
rect -10808 15277 -9992 15293
rect -9150 15293 -9134 15310
rect -8350 15310 -7942 15327
rect -7884 15327 -6284 15374
rect -7884 15310 -7476 15327
rect -8350 15293 -8334 15310
rect -9150 15277 -8334 15293
rect -7492 15293 -7476 15310
rect -6692 15310 -6284 15327
rect -6226 15327 -4626 15374
rect -6226 15310 -5818 15327
rect -6692 15293 -6676 15310
rect -7492 15277 -6676 15293
rect -5834 15293 -5818 15310
rect -5034 15310 -4626 15327
rect -4568 15327 -2968 15374
rect -4568 15310 -4160 15327
rect -5034 15293 -5018 15310
rect -5834 15277 -5018 15293
rect -4176 15293 -4160 15310
rect -3376 15310 -2968 15327
rect -2910 15327 -1310 15374
rect -2910 15310 -2502 15327
rect -3376 15293 -3360 15310
rect -4176 15277 -3360 15293
rect -2518 15293 -2502 15310
rect -1718 15310 -1310 15327
rect -1252 15327 348 15374
rect -1252 15310 -844 15327
rect -1718 15293 -1702 15310
rect -2518 15277 -1702 15293
rect -860 15293 -844 15310
rect -60 15310 348 15327
rect 406 15327 2006 15374
rect 406 15310 814 15327
rect -60 15293 -44 15310
rect -860 15277 -44 15293
rect 798 15293 814 15310
rect 1598 15310 2006 15327
rect 2064 15327 3664 15374
rect 2064 15310 2472 15327
rect 1598 15293 1614 15310
rect 798 15277 1614 15293
rect 2456 15293 2472 15310
rect 3256 15310 3664 15327
rect 3722 15327 5322 15374
rect 3722 15310 4130 15327
rect 3256 15293 3272 15310
rect 2456 15277 3272 15293
rect 4114 15293 4130 15310
rect 4914 15310 5322 15327
rect 5380 15327 6980 15374
rect 5380 15310 5788 15327
rect 4914 15293 4930 15310
rect 4114 15277 4930 15293
rect 5772 15293 5788 15310
rect 6572 15310 6980 15327
rect 7038 15327 8638 15374
rect 7038 15310 7446 15327
rect 6572 15293 6588 15310
rect 5772 15277 6588 15293
rect 7430 15293 7446 15310
rect 8230 15310 8638 15327
rect 8696 15327 10296 15374
rect 8696 15310 9104 15327
rect 8230 15293 8246 15310
rect 7430 15277 8246 15293
rect 9088 15293 9104 15310
rect 9888 15310 10296 15327
rect 10354 15327 11954 15374
rect 10354 15310 10762 15327
rect 9888 15293 9904 15310
rect 9088 15277 9904 15293
rect 10746 15293 10762 15310
rect 11546 15310 11954 15327
rect 12012 15327 13612 15374
rect 12012 15310 12420 15327
rect 11546 15293 11562 15310
rect 10746 15277 11562 15293
rect 12404 15293 12420 15310
rect 13204 15310 13612 15327
rect 13670 15327 15270 15374
rect 13670 15310 14078 15327
rect 13204 15293 13220 15310
rect 12404 15277 13220 15293
rect 14062 15293 14078 15310
rect 14862 15310 15270 15327
rect 15328 15327 16928 15374
rect 15328 15310 15736 15327
rect 14862 15293 14878 15310
rect 14062 15277 14878 15293
rect 15720 15293 15736 15310
rect 16520 15310 16928 15327
rect 16986 15327 18586 15374
rect 16986 15310 17394 15327
rect 16520 15293 16536 15310
rect 15720 15277 16536 15293
rect 17378 15293 17394 15310
rect 18178 15310 18586 15327
rect 18644 15327 20244 15374
rect 18644 15310 19052 15327
rect 18178 15293 18194 15310
rect 17378 15277 18194 15293
rect 19036 15293 19052 15310
rect 19836 15310 20244 15327
rect 20302 15327 21902 15374
rect 20302 15310 20710 15327
rect 19836 15293 19852 15310
rect 19036 15277 19852 15293
rect 20694 15293 20710 15310
rect 21494 15310 21902 15327
rect 21960 15327 23560 15374
rect 21960 15310 22368 15327
rect 21494 15293 21510 15310
rect 20694 15277 21510 15293
rect 22352 15293 22368 15310
rect 23152 15310 23560 15327
rect 23618 15327 25218 15374
rect 23618 15310 24026 15327
rect 23152 15293 23168 15310
rect 22352 15277 23168 15293
rect 24010 15293 24026 15310
rect 24810 15310 25218 15327
rect 25276 15327 26876 15374
rect 25276 15310 25684 15327
rect 24810 15293 24826 15310
rect 24010 15277 24826 15293
rect 25668 15293 25684 15310
rect 26468 15310 26876 15327
rect 26934 15327 28534 15374
rect 26934 15310 27342 15327
rect 26468 15293 26484 15310
rect 25668 15277 26484 15293
rect 27326 15293 27342 15310
rect 28126 15310 28534 15327
rect 28592 15327 30192 15374
rect 28592 15310 29000 15327
rect 28126 15293 28142 15310
rect 27326 15277 28142 15293
rect 28984 15293 29000 15310
rect 29784 15310 30192 15327
rect 30250 15327 31850 15374
rect 30250 15310 30658 15327
rect 29784 15293 29800 15310
rect 28984 15277 29800 15293
rect 30642 15293 30658 15310
rect 31442 15310 31850 15327
rect 31908 15327 33508 15374
rect 31908 15310 32316 15327
rect 31442 15293 31458 15310
rect 30642 15277 31458 15293
rect 32300 15293 32316 15310
rect 33100 15310 33508 15327
rect 33100 15293 33116 15310
rect 32300 15277 33116 15293
rect -32362 15219 -31546 15235
rect -32362 15202 -32346 15219
rect -32754 15185 -32346 15202
rect -31562 15202 -31546 15219
rect -30704 15219 -29888 15235
rect -30704 15202 -30688 15219
rect -31562 15185 -31154 15202
rect -32754 15138 -31154 15185
rect -31096 15185 -30688 15202
rect -29904 15202 -29888 15219
rect -29046 15219 -28230 15235
rect -29046 15202 -29030 15219
rect -29904 15185 -29496 15202
rect -31096 15138 -29496 15185
rect -29438 15185 -29030 15202
rect -28246 15202 -28230 15219
rect -27388 15219 -26572 15235
rect -27388 15202 -27372 15219
rect -28246 15185 -27838 15202
rect -29438 15138 -27838 15185
rect -27780 15185 -27372 15202
rect -26588 15202 -26572 15219
rect -25730 15219 -24914 15235
rect -25730 15202 -25714 15219
rect -26588 15185 -26180 15202
rect -27780 15138 -26180 15185
rect -26122 15185 -25714 15202
rect -24930 15202 -24914 15219
rect -24072 15219 -23256 15235
rect -24072 15202 -24056 15219
rect -24930 15185 -24522 15202
rect -26122 15138 -24522 15185
rect -24464 15185 -24056 15202
rect -23272 15202 -23256 15219
rect -22414 15219 -21598 15235
rect -22414 15202 -22398 15219
rect -23272 15185 -22864 15202
rect -24464 15138 -22864 15185
rect -22806 15185 -22398 15202
rect -21614 15202 -21598 15219
rect -20756 15219 -19940 15235
rect -20756 15202 -20740 15219
rect -21614 15185 -21206 15202
rect -22806 15138 -21206 15185
rect -21148 15185 -20740 15202
rect -19956 15202 -19940 15219
rect -19098 15219 -18282 15235
rect -19098 15202 -19082 15219
rect -19956 15185 -19548 15202
rect -21148 15138 -19548 15185
rect -19490 15185 -19082 15202
rect -18298 15202 -18282 15219
rect -17440 15219 -16624 15235
rect -17440 15202 -17424 15219
rect -18298 15185 -17890 15202
rect -19490 15138 -17890 15185
rect -17832 15185 -17424 15202
rect -16640 15202 -16624 15219
rect -15782 15219 -14966 15235
rect -15782 15202 -15766 15219
rect -16640 15185 -16232 15202
rect -17832 15138 -16232 15185
rect -16174 15185 -15766 15202
rect -14982 15202 -14966 15219
rect -14124 15219 -13308 15235
rect -14124 15202 -14108 15219
rect -14982 15185 -14574 15202
rect -16174 15138 -14574 15185
rect -14516 15185 -14108 15202
rect -13324 15202 -13308 15219
rect -12466 15219 -11650 15235
rect -12466 15202 -12450 15219
rect -13324 15185 -12916 15202
rect -14516 15138 -12916 15185
rect -12858 15185 -12450 15202
rect -11666 15202 -11650 15219
rect -10808 15219 -9992 15235
rect -10808 15202 -10792 15219
rect -11666 15185 -11258 15202
rect -12858 15138 -11258 15185
rect -11200 15185 -10792 15202
rect -10008 15202 -9992 15219
rect -9150 15219 -8334 15235
rect -9150 15202 -9134 15219
rect -10008 15185 -9600 15202
rect -11200 15138 -9600 15185
rect -9542 15185 -9134 15202
rect -8350 15202 -8334 15219
rect -7492 15219 -6676 15235
rect -7492 15202 -7476 15219
rect -8350 15185 -7942 15202
rect -9542 15138 -7942 15185
rect -7884 15185 -7476 15202
rect -6692 15202 -6676 15219
rect -5834 15219 -5018 15235
rect -5834 15202 -5818 15219
rect -6692 15185 -6284 15202
rect -7884 15138 -6284 15185
rect -6226 15185 -5818 15202
rect -5034 15202 -5018 15219
rect -4176 15219 -3360 15235
rect -4176 15202 -4160 15219
rect -5034 15185 -4626 15202
rect -6226 15138 -4626 15185
rect -4568 15185 -4160 15202
rect -3376 15202 -3360 15219
rect -2518 15219 -1702 15235
rect -2518 15202 -2502 15219
rect -3376 15185 -2968 15202
rect -4568 15138 -2968 15185
rect -2910 15185 -2502 15202
rect -1718 15202 -1702 15219
rect -860 15219 -44 15235
rect -860 15202 -844 15219
rect -1718 15185 -1310 15202
rect -2910 15138 -1310 15185
rect -1252 15185 -844 15202
rect -60 15202 -44 15219
rect 798 15219 1614 15235
rect 798 15202 814 15219
rect -60 15185 348 15202
rect -1252 15138 348 15185
rect 406 15185 814 15202
rect 1598 15202 1614 15219
rect 2456 15219 3272 15235
rect 2456 15202 2472 15219
rect 1598 15185 2006 15202
rect 406 15138 2006 15185
rect 2064 15185 2472 15202
rect 3256 15202 3272 15219
rect 4114 15219 4930 15235
rect 4114 15202 4130 15219
rect 3256 15185 3664 15202
rect 2064 15138 3664 15185
rect 3722 15185 4130 15202
rect 4914 15202 4930 15219
rect 5772 15219 6588 15235
rect 5772 15202 5788 15219
rect 4914 15185 5322 15202
rect 3722 15138 5322 15185
rect 5380 15185 5788 15202
rect 6572 15202 6588 15219
rect 7430 15219 8246 15235
rect 7430 15202 7446 15219
rect 6572 15185 6980 15202
rect 5380 15138 6980 15185
rect 7038 15185 7446 15202
rect 8230 15202 8246 15219
rect 9088 15219 9904 15235
rect 9088 15202 9104 15219
rect 8230 15185 8638 15202
rect 7038 15138 8638 15185
rect 8696 15185 9104 15202
rect 9888 15202 9904 15219
rect 10746 15219 11562 15235
rect 10746 15202 10762 15219
rect 9888 15185 10296 15202
rect 8696 15138 10296 15185
rect 10354 15185 10762 15202
rect 11546 15202 11562 15219
rect 12404 15219 13220 15235
rect 12404 15202 12420 15219
rect 11546 15185 11954 15202
rect 10354 15138 11954 15185
rect 12012 15185 12420 15202
rect 13204 15202 13220 15219
rect 14062 15219 14878 15235
rect 14062 15202 14078 15219
rect 13204 15185 13612 15202
rect 12012 15138 13612 15185
rect 13670 15185 14078 15202
rect 14862 15202 14878 15219
rect 15720 15219 16536 15235
rect 15720 15202 15736 15219
rect 14862 15185 15270 15202
rect 13670 15138 15270 15185
rect 15328 15185 15736 15202
rect 16520 15202 16536 15219
rect 17378 15219 18194 15235
rect 17378 15202 17394 15219
rect 16520 15185 16928 15202
rect 15328 15138 16928 15185
rect 16986 15185 17394 15202
rect 18178 15202 18194 15219
rect 19036 15219 19852 15235
rect 19036 15202 19052 15219
rect 18178 15185 18586 15202
rect 16986 15138 18586 15185
rect 18644 15185 19052 15202
rect 19836 15202 19852 15219
rect 20694 15219 21510 15235
rect 20694 15202 20710 15219
rect 19836 15185 20244 15202
rect 18644 15138 20244 15185
rect 20302 15185 20710 15202
rect 21494 15202 21510 15219
rect 22352 15219 23168 15235
rect 22352 15202 22368 15219
rect 21494 15185 21902 15202
rect 20302 15138 21902 15185
rect 21960 15185 22368 15202
rect 23152 15202 23168 15219
rect 24010 15219 24826 15235
rect 24010 15202 24026 15219
rect 23152 15185 23560 15202
rect 21960 15138 23560 15185
rect 23618 15185 24026 15202
rect 24810 15202 24826 15219
rect 25668 15219 26484 15235
rect 25668 15202 25684 15219
rect 24810 15185 25218 15202
rect 23618 15138 25218 15185
rect 25276 15185 25684 15202
rect 26468 15202 26484 15219
rect 27326 15219 28142 15235
rect 27326 15202 27342 15219
rect 26468 15185 26876 15202
rect 25276 15138 26876 15185
rect 26934 15185 27342 15202
rect 28126 15202 28142 15219
rect 28984 15219 29800 15235
rect 28984 15202 29000 15219
rect 28126 15185 28534 15202
rect 26934 15138 28534 15185
rect 28592 15185 29000 15202
rect 29784 15202 29800 15219
rect 30642 15219 31458 15235
rect 30642 15202 30658 15219
rect 29784 15185 30192 15202
rect 28592 15138 30192 15185
rect 30250 15185 30658 15202
rect 31442 15202 31458 15219
rect 32300 15219 33116 15235
rect 32300 15202 32316 15219
rect 31442 15185 31850 15202
rect 30250 15138 31850 15185
rect 31908 15185 32316 15202
rect 33100 15202 33116 15219
rect 33100 15185 33508 15202
rect 31908 15138 33508 15185
rect -32754 13691 -31154 13738
rect -32754 13674 -32346 13691
rect -32362 13657 -32346 13674
rect -31562 13674 -31154 13691
rect -31096 13691 -29496 13738
rect -31096 13674 -30688 13691
rect -31562 13657 -31546 13674
rect -32362 13641 -31546 13657
rect -30704 13657 -30688 13674
rect -29904 13674 -29496 13691
rect -29438 13691 -27838 13738
rect -29438 13674 -29030 13691
rect -29904 13657 -29888 13674
rect -30704 13641 -29888 13657
rect -29046 13657 -29030 13674
rect -28246 13674 -27838 13691
rect -27780 13691 -26180 13738
rect -27780 13674 -27372 13691
rect -28246 13657 -28230 13674
rect -29046 13641 -28230 13657
rect -27388 13657 -27372 13674
rect -26588 13674 -26180 13691
rect -26122 13691 -24522 13738
rect -26122 13674 -25714 13691
rect -26588 13657 -26572 13674
rect -27388 13641 -26572 13657
rect -25730 13657 -25714 13674
rect -24930 13674 -24522 13691
rect -24464 13691 -22864 13738
rect -24464 13674 -24056 13691
rect -24930 13657 -24914 13674
rect -25730 13641 -24914 13657
rect -24072 13657 -24056 13674
rect -23272 13674 -22864 13691
rect -22806 13691 -21206 13738
rect -22806 13674 -22398 13691
rect -23272 13657 -23256 13674
rect -24072 13641 -23256 13657
rect -22414 13657 -22398 13674
rect -21614 13674 -21206 13691
rect -21148 13691 -19548 13738
rect -21148 13674 -20740 13691
rect -21614 13657 -21598 13674
rect -22414 13641 -21598 13657
rect -20756 13657 -20740 13674
rect -19956 13674 -19548 13691
rect -19490 13691 -17890 13738
rect -19490 13674 -19082 13691
rect -19956 13657 -19940 13674
rect -20756 13641 -19940 13657
rect -19098 13657 -19082 13674
rect -18298 13674 -17890 13691
rect -17832 13691 -16232 13738
rect -17832 13674 -17424 13691
rect -18298 13657 -18282 13674
rect -19098 13641 -18282 13657
rect -17440 13657 -17424 13674
rect -16640 13674 -16232 13691
rect -16174 13691 -14574 13738
rect -16174 13674 -15766 13691
rect -16640 13657 -16624 13674
rect -17440 13641 -16624 13657
rect -15782 13657 -15766 13674
rect -14982 13674 -14574 13691
rect -14516 13691 -12916 13738
rect -14516 13674 -14108 13691
rect -14982 13657 -14966 13674
rect -15782 13641 -14966 13657
rect -14124 13657 -14108 13674
rect -13324 13674 -12916 13691
rect -12858 13691 -11258 13738
rect -12858 13674 -12450 13691
rect -13324 13657 -13308 13674
rect -14124 13641 -13308 13657
rect -12466 13657 -12450 13674
rect -11666 13674 -11258 13691
rect -11200 13691 -9600 13738
rect -11200 13674 -10792 13691
rect -11666 13657 -11650 13674
rect -12466 13641 -11650 13657
rect -10808 13657 -10792 13674
rect -10008 13674 -9600 13691
rect -9542 13691 -7942 13738
rect -9542 13674 -9134 13691
rect -10008 13657 -9992 13674
rect -10808 13641 -9992 13657
rect -9150 13657 -9134 13674
rect -8350 13674 -7942 13691
rect -7884 13691 -6284 13738
rect -7884 13674 -7476 13691
rect -8350 13657 -8334 13674
rect -9150 13641 -8334 13657
rect -7492 13657 -7476 13674
rect -6692 13674 -6284 13691
rect -6226 13691 -4626 13738
rect -6226 13674 -5818 13691
rect -6692 13657 -6676 13674
rect -7492 13641 -6676 13657
rect -5834 13657 -5818 13674
rect -5034 13674 -4626 13691
rect -4568 13691 -2968 13738
rect -4568 13674 -4160 13691
rect -5034 13657 -5018 13674
rect -5834 13641 -5018 13657
rect -4176 13657 -4160 13674
rect -3376 13674 -2968 13691
rect -2910 13691 -1310 13738
rect -2910 13674 -2502 13691
rect -3376 13657 -3360 13674
rect -4176 13641 -3360 13657
rect -2518 13657 -2502 13674
rect -1718 13674 -1310 13691
rect -1252 13691 348 13738
rect -1252 13674 -844 13691
rect -1718 13657 -1702 13674
rect -2518 13641 -1702 13657
rect -860 13657 -844 13674
rect -60 13674 348 13691
rect 406 13691 2006 13738
rect 406 13674 814 13691
rect -60 13657 -44 13674
rect -860 13641 -44 13657
rect 798 13657 814 13674
rect 1598 13674 2006 13691
rect 2064 13691 3664 13738
rect 2064 13674 2472 13691
rect 1598 13657 1614 13674
rect 798 13641 1614 13657
rect 2456 13657 2472 13674
rect 3256 13674 3664 13691
rect 3722 13691 5322 13738
rect 3722 13674 4130 13691
rect 3256 13657 3272 13674
rect 2456 13641 3272 13657
rect 4114 13657 4130 13674
rect 4914 13674 5322 13691
rect 5380 13691 6980 13738
rect 5380 13674 5788 13691
rect 4914 13657 4930 13674
rect 4114 13641 4930 13657
rect 5772 13657 5788 13674
rect 6572 13674 6980 13691
rect 7038 13691 8638 13738
rect 7038 13674 7446 13691
rect 6572 13657 6588 13674
rect 5772 13641 6588 13657
rect 7430 13657 7446 13674
rect 8230 13674 8638 13691
rect 8696 13691 10296 13738
rect 8696 13674 9104 13691
rect 8230 13657 8246 13674
rect 7430 13641 8246 13657
rect 9088 13657 9104 13674
rect 9888 13674 10296 13691
rect 10354 13691 11954 13738
rect 10354 13674 10762 13691
rect 9888 13657 9904 13674
rect 9088 13641 9904 13657
rect 10746 13657 10762 13674
rect 11546 13674 11954 13691
rect 12012 13691 13612 13738
rect 12012 13674 12420 13691
rect 11546 13657 11562 13674
rect 10746 13641 11562 13657
rect 12404 13657 12420 13674
rect 13204 13674 13612 13691
rect 13670 13691 15270 13738
rect 13670 13674 14078 13691
rect 13204 13657 13220 13674
rect 12404 13641 13220 13657
rect 14062 13657 14078 13674
rect 14862 13674 15270 13691
rect 15328 13691 16928 13738
rect 15328 13674 15736 13691
rect 14862 13657 14878 13674
rect 14062 13641 14878 13657
rect 15720 13657 15736 13674
rect 16520 13674 16928 13691
rect 16986 13691 18586 13738
rect 16986 13674 17394 13691
rect 16520 13657 16536 13674
rect 15720 13641 16536 13657
rect 17378 13657 17394 13674
rect 18178 13674 18586 13691
rect 18644 13691 20244 13738
rect 18644 13674 19052 13691
rect 18178 13657 18194 13674
rect 17378 13641 18194 13657
rect 19036 13657 19052 13674
rect 19836 13674 20244 13691
rect 20302 13691 21902 13738
rect 20302 13674 20710 13691
rect 19836 13657 19852 13674
rect 19036 13641 19852 13657
rect 20694 13657 20710 13674
rect 21494 13674 21902 13691
rect 21960 13691 23560 13738
rect 21960 13674 22368 13691
rect 21494 13657 21510 13674
rect 20694 13641 21510 13657
rect 22352 13657 22368 13674
rect 23152 13674 23560 13691
rect 23618 13691 25218 13738
rect 23618 13674 24026 13691
rect 23152 13657 23168 13674
rect 22352 13641 23168 13657
rect 24010 13657 24026 13674
rect 24810 13674 25218 13691
rect 25276 13691 26876 13738
rect 25276 13674 25684 13691
rect 24810 13657 24826 13674
rect 24010 13641 24826 13657
rect 25668 13657 25684 13674
rect 26468 13674 26876 13691
rect 26934 13691 28534 13738
rect 26934 13674 27342 13691
rect 26468 13657 26484 13674
rect 25668 13641 26484 13657
rect 27326 13657 27342 13674
rect 28126 13674 28534 13691
rect 28592 13691 30192 13738
rect 28592 13674 29000 13691
rect 28126 13657 28142 13674
rect 27326 13641 28142 13657
rect 28984 13657 29000 13674
rect 29784 13674 30192 13691
rect 30250 13691 31850 13738
rect 30250 13674 30658 13691
rect 29784 13657 29800 13674
rect 28984 13641 29800 13657
rect 30642 13657 30658 13674
rect 31442 13674 31850 13691
rect 31908 13691 33508 13738
rect 31908 13674 32316 13691
rect 31442 13657 31458 13674
rect 30642 13641 31458 13657
rect 32300 13657 32316 13674
rect 33100 13674 33508 13691
rect 33100 13657 33116 13674
rect 32300 13641 33116 13657
rect -32360 13473 -31544 13489
rect -32360 13456 -32344 13473
rect -32752 13439 -32344 13456
rect -31560 13456 -31544 13473
rect -30702 13473 -29886 13489
rect -30702 13456 -30686 13473
rect -31560 13439 -31152 13456
rect -32752 13392 -31152 13439
rect -31094 13439 -30686 13456
rect -29902 13456 -29886 13473
rect -29044 13473 -28228 13489
rect -29044 13456 -29028 13473
rect -29902 13439 -29494 13456
rect -31094 13392 -29494 13439
rect -29436 13439 -29028 13456
rect -28244 13456 -28228 13473
rect -27386 13473 -26570 13489
rect -27386 13456 -27370 13473
rect -28244 13439 -27836 13456
rect -29436 13392 -27836 13439
rect -27778 13439 -27370 13456
rect -26586 13456 -26570 13473
rect -25728 13473 -24912 13489
rect -25728 13456 -25712 13473
rect -26586 13439 -26178 13456
rect -27778 13392 -26178 13439
rect -26120 13439 -25712 13456
rect -24928 13456 -24912 13473
rect -24070 13473 -23254 13489
rect -24070 13456 -24054 13473
rect -24928 13439 -24520 13456
rect -26120 13392 -24520 13439
rect -24462 13439 -24054 13456
rect -23270 13456 -23254 13473
rect -22412 13473 -21596 13489
rect -22412 13456 -22396 13473
rect -23270 13439 -22862 13456
rect -24462 13392 -22862 13439
rect -22804 13439 -22396 13456
rect -21612 13456 -21596 13473
rect -20754 13473 -19938 13489
rect -20754 13456 -20738 13473
rect -21612 13439 -21204 13456
rect -22804 13392 -21204 13439
rect -21146 13439 -20738 13456
rect -19954 13456 -19938 13473
rect -19096 13473 -18280 13489
rect -19096 13456 -19080 13473
rect -19954 13439 -19546 13456
rect -21146 13392 -19546 13439
rect -19488 13439 -19080 13456
rect -18296 13456 -18280 13473
rect -17438 13473 -16622 13489
rect -17438 13456 -17422 13473
rect -18296 13439 -17888 13456
rect -19488 13392 -17888 13439
rect -17830 13439 -17422 13456
rect -16638 13456 -16622 13473
rect -15780 13473 -14964 13489
rect -15780 13456 -15764 13473
rect -16638 13439 -16230 13456
rect -17830 13392 -16230 13439
rect -16172 13439 -15764 13456
rect -14980 13456 -14964 13473
rect -14122 13473 -13306 13489
rect -14122 13456 -14106 13473
rect -14980 13439 -14572 13456
rect -16172 13392 -14572 13439
rect -14514 13439 -14106 13456
rect -13322 13456 -13306 13473
rect -12464 13473 -11648 13489
rect -12464 13456 -12448 13473
rect -13322 13439 -12914 13456
rect -14514 13392 -12914 13439
rect -12856 13439 -12448 13456
rect -11664 13456 -11648 13473
rect -10806 13473 -9990 13489
rect -10806 13456 -10790 13473
rect -11664 13439 -11256 13456
rect -12856 13392 -11256 13439
rect -11198 13439 -10790 13456
rect -10006 13456 -9990 13473
rect -9148 13473 -8332 13489
rect -9148 13456 -9132 13473
rect -10006 13439 -9598 13456
rect -11198 13392 -9598 13439
rect -9540 13439 -9132 13456
rect -8348 13456 -8332 13473
rect -7490 13473 -6674 13489
rect -7490 13456 -7474 13473
rect -8348 13439 -7940 13456
rect -9540 13392 -7940 13439
rect -7882 13439 -7474 13456
rect -6690 13456 -6674 13473
rect -5832 13473 -5016 13489
rect -5832 13456 -5816 13473
rect -6690 13439 -6282 13456
rect -7882 13392 -6282 13439
rect -6224 13439 -5816 13456
rect -5032 13456 -5016 13473
rect -4174 13473 -3358 13489
rect -4174 13456 -4158 13473
rect -5032 13439 -4624 13456
rect -6224 13392 -4624 13439
rect -4566 13439 -4158 13456
rect -3374 13456 -3358 13473
rect -2516 13473 -1700 13489
rect -2516 13456 -2500 13473
rect -3374 13439 -2966 13456
rect -4566 13392 -2966 13439
rect -2908 13439 -2500 13456
rect -1716 13456 -1700 13473
rect -858 13473 -42 13489
rect -858 13456 -842 13473
rect -1716 13439 -1308 13456
rect -2908 13392 -1308 13439
rect -1250 13439 -842 13456
rect -58 13456 -42 13473
rect 800 13473 1616 13489
rect 800 13456 816 13473
rect -58 13439 350 13456
rect -1250 13392 350 13439
rect 408 13439 816 13456
rect 1600 13456 1616 13473
rect 2458 13473 3274 13489
rect 2458 13456 2474 13473
rect 1600 13439 2008 13456
rect 408 13392 2008 13439
rect 2066 13439 2474 13456
rect 3258 13456 3274 13473
rect 4116 13473 4932 13489
rect 4116 13456 4132 13473
rect 3258 13439 3666 13456
rect 2066 13392 3666 13439
rect 3724 13439 4132 13456
rect 4916 13456 4932 13473
rect 5774 13473 6590 13489
rect 5774 13456 5790 13473
rect 4916 13439 5324 13456
rect 3724 13392 5324 13439
rect 5382 13439 5790 13456
rect 6574 13456 6590 13473
rect 7432 13473 8248 13489
rect 7432 13456 7448 13473
rect 6574 13439 6982 13456
rect 5382 13392 6982 13439
rect 7040 13439 7448 13456
rect 8232 13456 8248 13473
rect 9090 13473 9906 13489
rect 9090 13456 9106 13473
rect 8232 13439 8640 13456
rect 7040 13392 8640 13439
rect 8698 13439 9106 13456
rect 9890 13456 9906 13473
rect 10748 13473 11564 13489
rect 10748 13456 10764 13473
rect 9890 13439 10298 13456
rect 8698 13392 10298 13439
rect 10356 13439 10764 13456
rect 11548 13456 11564 13473
rect 12406 13473 13222 13489
rect 12406 13456 12422 13473
rect 11548 13439 11956 13456
rect 10356 13392 11956 13439
rect 12014 13439 12422 13456
rect 13206 13456 13222 13473
rect 14064 13473 14880 13489
rect 14064 13456 14080 13473
rect 13206 13439 13614 13456
rect 12014 13392 13614 13439
rect 13672 13439 14080 13456
rect 14864 13456 14880 13473
rect 15722 13473 16538 13489
rect 15722 13456 15738 13473
rect 14864 13439 15272 13456
rect 13672 13392 15272 13439
rect 15330 13439 15738 13456
rect 16522 13456 16538 13473
rect 17380 13473 18196 13489
rect 17380 13456 17396 13473
rect 16522 13439 16930 13456
rect 15330 13392 16930 13439
rect 16988 13439 17396 13456
rect 18180 13456 18196 13473
rect 19038 13473 19854 13489
rect 19038 13456 19054 13473
rect 18180 13439 18588 13456
rect 16988 13392 18588 13439
rect 18646 13439 19054 13456
rect 19838 13456 19854 13473
rect 20696 13473 21512 13489
rect 20696 13456 20712 13473
rect 19838 13439 20246 13456
rect 18646 13392 20246 13439
rect 20304 13439 20712 13456
rect 21496 13456 21512 13473
rect 22354 13473 23170 13489
rect 22354 13456 22370 13473
rect 21496 13439 21904 13456
rect 20304 13392 21904 13439
rect 21962 13439 22370 13456
rect 23154 13456 23170 13473
rect 24012 13473 24828 13489
rect 24012 13456 24028 13473
rect 23154 13439 23562 13456
rect 21962 13392 23562 13439
rect 23620 13439 24028 13456
rect 24812 13456 24828 13473
rect 25670 13473 26486 13489
rect 25670 13456 25686 13473
rect 24812 13439 25220 13456
rect 23620 13392 25220 13439
rect 25278 13439 25686 13456
rect 26470 13456 26486 13473
rect 27328 13473 28144 13489
rect 27328 13456 27344 13473
rect 26470 13439 26878 13456
rect 25278 13392 26878 13439
rect 26936 13439 27344 13456
rect 28128 13456 28144 13473
rect 28986 13473 29802 13489
rect 28986 13456 29002 13473
rect 28128 13439 28536 13456
rect 26936 13392 28536 13439
rect 28594 13439 29002 13456
rect 29786 13456 29802 13473
rect 30644 13473 31460 13489
rect 30644 13456 30660 13473
rect 29786 13439 30194 13456
rect 28594 13392 30194 13439
rect 30252 13439 30660 13456
rect 31444 13456 31460 13473
rect 32302 13473 33118 13489
rect 32302 13456 32318 13473
rect 31444 13439 31852 13456
rect 30252 13392 31852 13439
rect 31910 13439 32318 13456
rect 33102 13456 33118 13473
rect 33102 13439 33510 13456
rect 31910 13392 33510 13439
rect -32752 11945 -31152 11992
rect -32752 11928 -32344 11945
rect -32360 11911 -32344 11928
rect -31560 11928 -31152 11945
rect -31094 11945 -29494 11992
rect -31094 11928 -30686 11945
rect -31560 11911 -31544 11928
rect -32360 11895 -31544 11911
rect -30702 11911 -30686 11928
rect -29902 11928 -29494 11945
rect -29436 11945 -27836 11992
rect -29436 11928 -29028 11945
rect -29902 11911 -29886 11928
rect -30702 11895 -29886 11911
rect -29044 11911 -29028 11928
rect -28244 11928 -27836 11945
rect -27778 11945 -26178 11992
rect -27778 11928 -27370 11945
rect -28244 11911 -28228 11928
rect -29044 11895 -28228 11911
rect -27386 11911 -27370 11928
rect -26586 11928 -26178 11945
rect -26120 11945 -24520 11992
rect -26120 11928 -25712 11945
rect -26586 11911 -26570 11928
rect -27386 11895 -26570 11911
rect -25728 11911 -25712 11928
rect -24928 11928 -24520 11945
rect -24462 11945 -22862 11992
rect -24462 11928 -24054 11945
rect -24928 11911 -24912 11928
rect -25728 11895 -24912 11911
rect -24070 11911 -24054 11928
rect -23270 11928 -22862 11945
rect -22804 11945 -21204 11992
rect -22804 11928 -22396 11945
rect -23270 11911 -23254 11928
rect -24070 11895 -23254 11911
rect -22412 11911 -22396 11928
rect -21612 11928 -21204 11945
rect -21146 11945 -19546 11992
rect -21146 11928 -20738 11945
rect -21612 11911 -21596 11928
rect -22412 11895 -21596 11911
rect -20754 11911 -20738 11928
rect -19954 11928 -19546 11945
rect -19488 11945 -17888 11992
rect -19488 11928 -19080 11945
rect -19954 11911 -19938 11928
rect -20754 11895 -19938 11911
rect -19096 11911 -19080 11928
rect -18296 11928 -17888 11945
rect -17830 11945 -16230 11992
rect -17830 11928 -17422 11945
rect -18296 11911 -18280 11928
rect -19096 11895 -18280 11911
rect -17438 11911 -17422 11928
rect -16638 11928 -16230 11945
rect -16172 11945 -14572 11992
rect -16172 11928 -15764 11945
rect -16638 11911 -16622 11928
rect -17438 11895 -16622 11911
rect -15780 11911 -15764 11928
rect -14980 11928 -14572 11945
rect -14514 11945 -12914 11992
rect -14514 11928 -14106 11945
rect -14980 11911 -14964 11928
rect -15780 11895 -14964 11911
rect -14122 11911 -14106 11928
rect -13322 11928 -12914 11945
rect -12856 11945 -11256 11992
rect -12856 11928 -12448 11945
rect -13322 11911 -13306 11928
rect -14122 11895 -13306 11911
rect -12464 11911 -12448 11928
rect -11664 11928 -11256 11945
rect -11198 11945 -9598 11992
rect -11198 11928 -10790 11945
rect -11664 11911 -11648 11928
rect -12464 11895 -11648 11911
rect -10806 11911 -10790 11928
rect -10006 11928 -9598 11945
rect -9540 11945 -7940 11992
rect -9540 11928 -9132 11945
rect -10006 11911 -9990 11928
rect -10806 11895 -9990 11911
rect -9148 11911 -9132 11928
rect -8348 11928 -7940 11945
rect -7882 11945 -6282 11992
rect -7882 11928 -7474 11945
rect -8348 11911 -8332 11928
rect -9148 11895 -8332 11911
rect -7490 11911 -7474 11928
rect -6690 11928 -6282 11945
rect -6224 11945 -4624 11992
rect -6224 11928 -5816 11945
rect -6690 11911 -6674 11928
rect -7490 11895 -6674 11911
rect -5832 11911 -5816 11928
rect -5032 11928 -4624 11945
rect -4566 11945 -2966 11992
rect -4566 11928 -4158 11945
rect -5032 11911 -5016 11928
rect -5832 11895 -5016 11911
rect -4174 11911 -4158 11928
rect -3374 11928 -2966 11945
rect -2908 11945 -1308 11992
rect -2908 11928 -2500 11945
rect -3374 11911 -3358 11928
rect -4174 11895 -3358 11911
rect -2516 11911 -2500 11928
rect -1716 11928 -1308 11945
rect -1250 11945 350 11992
rect -1250 11928 -842 11945
rect -1716 11911 -1700 11928
rect -2516 11895 -1700 11911
rect -858 11911 -842 11928
rect -58 11928 350 11945
rect 408 11945 2008 11992
rect 408 11928 816 11945
rect -58 11911 -42 11928
rect -858 11895 -42 11911
rect 800 11911 816 11928
rect 1600 11928 2008 11945
rect 2066 11945 3666 11992
rect 2066 11928 2474 11945
rect 1600 11911 1616 11928
rect 800 11895 1616 11911
rect 2458 11911 2474 11928
rect 3258 11928 3666 11945
rect 3724 11945 5324 11992
rect 3724 11928 4132 11945
rect 3258 11911 3274 11928
rect 2458 11895 3274 11911
rect 4116 11911 4132 11928
rect 4916 11928 5324 11945
rect 5382 11945 6982 11992
rect 5382 11928 5790 11945
rect 4916 11911 4932 11928
rect 4116 11895 4932 11911
rect 5774 11911 5790 11928
rect 6574 11928 6982 11945
rect 7040 11945 8640 11992
rect 7040 11928 7448 11945
rect 6574 11911 6590 11928
rect 5774 11895 6590 11911
rect 7432 11911 7448 11928
rect 8232 11928 8640 11945
rect 8698 11945 10298 11992
rect 8698 11928 9106 11945
rect 8232 11911 8248 11928
rect 7432 11895 8248 11911
rect 9090 11911 9106 11928
rect 9890 11928 10298 11945
rect 10356 11945 11956 11992
rect 10356 11928 10764 11945
rect 9890 11911 9906 11928
rect 9090 11895 9906 11911
rect 10748 11911 10764 11928
rect 11548 11928 11956 11945
rect 12014 11945 13614 11992
rect 12014 11928 12422 11945
rect 11548 11911 11564 11928
rect 10748 11895 11564 11911
rect 12406 11911 12422 11928
rect 13206 11928 13614 11945
rect 13672 11945 15272 11992
rect 13672 11928 14080 11945
rect 13206 11911 13222 11928
rect 12406 11895 13222 11911
rect 14064 11911 14080 11928
rect 14864 11928 15272 11945
rect 15330 11945 16930 11992
rect 15330 11928 15738 11945
rect 14864 11911 14880 11928
rect 14064 11895 14880 11911
rect 15722 11911 15738 11928
rect 16522 11928 16930 11945
rect 16988 11945 18588 11992
rect 16988 11928 17396 11945
rect 16522 11911 16538 11928
rect 15722 11895 16538 11911
rect 17380 11911 17396 11928
rect 18180 11928 18588 11945
rect 18646 11945 20246 11992
rect 18646 11928 19054 11945
rect 18180 11911 18196 11928
rect 17380 11895 18196 11911
rect 19038 11911 19054 11928
rect 19838 11928 20246 11945
rect 20304 11945 21904 11992
rect 20304 11928 20712 11945
rect 19838 11911 19854 11928
rect 19038 11895 19854 11911
rect 20696 11911 20712 11928
rect 21496 11928 21904 11945
rect 21962 11945 23562 11992
rect 21962 11928 22370 11945
rect 21496 11911 21512 11928
rect 20696 11895 21512 11911
rect 22354 11911 22370 11928
rect 23154 11928 23562 11945
rect 23620 11945 25220 11992
rect 23620 11928 24028 11945
rect 23154 11911 23170 11928
rect 22354 11895 23170 11911
rect 24012 11911 24028 11928
rect 24812 11928 25220 11945
rect 25278 11945 26878 11992
rect 25278 11928 25686 11945
rect 24812 11911 24828 11928
rect 24012 11895 24828 11911
rect 25670 11911 25686 11928
rect 26470 11928 26878 11945
rect 26936 11945 28536 11992
rect 26936 11928 27344 11945
rect 26470 11911 26486 11928
rect 25670 11895 26486 11911
rect 27328 11911 27344 11928
rect 28128 11928 28536 11945
rect 28594 11945 30194 11992
rect 28594 11928 29002 11945
rect 28128 11911 28144 11928
rect 27328 11895 28144 11911
rect 28986 11911 29002 11928
rect 29786 11928 30194 11945
rect 30252 11945 31852 11992
rect 30252 11928 30660 11945
rect 29786 11911 29802 11928
rect 28986 11895 29802 11911
rect 30644 11911 30660 11928
rect 31444 11928 31852 11945
rect 31910 11945 33510 11992
rect 31910 11928 32318 11945
rect 31444 11911 31460 11928
rect 30644 11895 31460 11911
rect 32302 11911 32318 11928
rect 33102 11928 33510 11945
rect 33102 11911 33118 11928
rect 32302 11895 33118 11911
rect -32360 11837 -31544 11853
rect -32360 11820 -32344 11837
rect -32752 11803 -32344 11820
rect -31560 11820 -31544 11837
rect -30702 11837 -29886 11853
rect -30702 11820 -30686 11837
rect -31560 11803 -31152 11820
rect -32752 11756 -31152 11803
rect -31094 11803 -30686 11820
rect -29902 11820 -29886 11837
rect -29044 11837 -28228 11853
rect -29044 11820 -29028 11837
rect -29902 11803 -29494 11820
rect -31094 11756 -29494 11803
rect -29436 11803 -29028 11820
rect -28244 11820 -28228 11837
rect -27386 11837 -26570 11853
rect -27386 11820 -27370 11837
rect -28244 11803 -27836 11820
rect -29436 11756 -27836 11803
rect -27778 11803 -27370 11820
rect -26586 11820 -26570 11837
rect -25728 11837 -24912 11853
rect -25728 11820 -25712 11837
rect -26586 11803 -26178 11820
rect -27778 11756 -26178 11803
rect -26120 11803 -25712 11820
rect -24928 11820 -24912 11837
rect -24070 11837 -23254 11853
rect -24070 11820 -24054 11837
rect -24928 11803 -24520 11820
rect -26120 11756 -24520 11803
rect -24462 11803 -24054 11820
rect -23270 11820 -23254 11837
rect -22412 11837 -21596 11853
rect -22412 11820 -22396 11837
rect -23270 11803 -22862 11820
rect -24462 11756 -22862 11803
rect -22804 11803 -22396 11820
rect -21612 11820 -21596 11837
rect -20754 11837 -19938 11853
rect -20754 11820 -20738 11837
rect -21612 11803 -21204 11820
rect -22804 11756 -21204 11803
rect -21146 11803 -20738 11820
rect -19954 11820 -19938 11837
rect -19096 11837 -18280 11853
rect -19096 11820 -19080 11837
rect -19954 11803 -19546 11820
rect -21146 11756 -19546 11803
rect -19488 11803 -19080 11820
rect -18296 11820 -18280 11837
rect -17438 11837 -16622 11853
rect -17438 11820 -17422 11837
rect -18296 11803 -17888 11820
rect -19488 11756 -17888 11803
rect -17830 11803 -17422 11820
rect -16638 11820 -16622 11837
rect -15780 11837 -14964 11853
rect -15780 11820 -15764 11837
rect -16638 11803 -16230 11820
rect -17830 11756 -16230 11803
rect -16172 11803 -15764 11820
rect -14980 11820 -14964 11837
rect -14122 11837 -13306 11853
rect -14122 11820 -14106 11837
rect -14980 11803 -14572 11820
rect -16172 11756 -14572 11803
rect -14514 11803 -14106 11820
rect -13322 11820 -13306 11837
rect -12464 11837 -11648 11853
rect -12464 11820 -12448 11837
rect -13322 11803 -12914 11820
rect -14514 11756 -12914 11803
rect -12856 11803 -12448 11820
rect -11664 11820 -11648 11837
rect -10806 11837 -9990 11853
rect -10806 11820 -10790 11837
rect -11664 11803 -11256 11820
rect -12856 11756 -11256 11803
rect -11198 11803 -10790 11820
rect -10006 11820 -9990 11837
rect -9148 11837 -8332 11853
rect -9148 11820 -9132 11837
rect -10006 11803 -9598 11820
rect -11198 11756 -9598 11803
rect -9540 11803 -9132 11820
rect -8348 11820 -8332 11837
rect -7490 11837 -6674 11853
rect -7490 11820 -7474 11837
rect -8348 11803 -7940 11820
rect -9540 11756 -7940 11803
rect -7882 11803 -7474 11820
rect -6690 11820 -6674 11837
rect -5832 11837 -5016 11853
rect -5832 11820 -5816 11837
rect -6690 11803 -6282 11820
rect -7882 11756 -6282 11803
rect -6224 11803 -5816 11820
rect -5032 11820 -5016 11837
rect -4174 11837 -3358 11853
rect -4174 11820 -4158 11837
rect -5032 11803 -4624 11820
rect -6224 11756 -4624 11803
rect -4566 11803 -4158 11820
rect -3374 11820 -3358 11837
rect -2516 11837 -1700 11853
rect -2516 11820 -2500 11837
rect -3374 11803 -2966 11820
rect -4566 11756 -2966 11803
rect -2908 11803 -2500 11820
rect -1716 11820 -1700 11837
rect -858 11837 -42 11853
rect -858 11820 -842 11837
rect -1716 11803 -1308 11820
rect -2908 11756 -1308 11803
rect -1250 11803 -842 11820
rect -58 11820 -42 11837
rect 800 11837 1616 11853
rect 800 11820 816 11837
rect -58 11803 350 11820
rect -1250 11756 350 11803
rect 408 11803 816 11820
rect 1600 11820 1616 11837
rect 2458 11837 3274 11853
rect 2458 11820 2474 11837
rect 1600 11803 2008 11820
rect 408 11756 2008 11803
rect 2066 11803 2474 11820
rect 3258 11820 3274 11837
rect 4116 11837 4932 11853
rect 4116 11820 4132 11837
rect 3258 11803 3666 11820
rect 2066 11756 3666 11803
rect 3724 11803 4132 11820
rect 4916 11820 4932 11837
rect 5774 11837 6590 11853
rect 5774 11820 5790 11837
rect 4916 11803 5324 11820
rect 3724 11756 5324 11803
rect 5382 11803 5790 11820
rect 6574 11820 6590 11837
rect 7432 11837 8248 11853
rect 7432 11820 7448 11837
rect 6574 11803 6982 11820
rect 5382 11756 6982 11803
rect 7040 11803 7448 11820
rect 8232 11820 8248 11837
rect 9090 11837 9906 11853
rect 9090 11820 9106 11837
rect 8232 11803 8640 11820
rect 7040 11756 8640 11803
rect 8698 11803 9106 11820
rect 9890 11820 9906 11837
rect 10748 11837 11564 11853
rect 10748 11820 10764 11837
rect 9890 11803 10298 11820
rect 8698 11756 10298 11803
rect 10356 11803 10764 11820
rect 11548 11820 11564 11837
rect 12406 11837 13222 11853
rect 12406 11820 12422 11837
rect 11548 11803 11956 11820
rect 10356 11756 11956 11803
rect 12014 11803 12422 11820
rect 13206 11820 13222 11837
rect 14064 11837 14880 11853
rect 14064 11820 14080 11837
rect 13206 11803 13614 11820
rect 12014 11756 13614 11803
rect 13672 11803 14080 11820
rect 14864 11820 14880 11837
rect 15722 11837 16538 11853
rect 15722 11820 15738 11837
rect 14864 11803 15272 11820
rect 13672 11756 15272 11803
rect 15330 11803 15738 11820
rect 16522 11820 16538 11837
rect 17380 11837 18196 11853
rect 17380 11820 17396 11837
rect 16522 11803 16930 11820
rect 15330 11756 16930 11803
rect 16988 11803 17396 11820
rect 18180 11820 18196 11837
rect 19038 11837 19854 11853
rect 19038 11820 19054 11837
rect 18180 11803 18588 11820
rect 16988 11756 18588 11803
rect 18646 11803 19054 11820
rect 19838 11820 19854 11837
rect 20696 11837 21512 11853
rect 20696 11820 20712 11837
rect 19838 11803 20246 11820
rect 18646 11756 20246 11803
rect 20304 11803 20712 11820
rect 21496 11820 21512 11837
rect 22354 11837 23170 11853
rect 22354 11820 22370 11837
rect 21496 11803 21904 11820
rect 20304 11756 21904 11803
rect 21962 11803 22370 11820
rect 23154 11820 23170 11837
rect 24012 11837 24828 11853
rect 24012 11820 24028 11837
rect 23154 11803 23562 11820
rect 21962 11756 23562 11803
rect 23620 11803 24028 11820
rect 24812 11820 24828 11837
rect 25670 11837 26486 11853
rect 25670 11820 25686 11837
rect 24812 11803 25220 11820
rect 23620 11756 25220 11803
rect 25278 11803 25686 11820
rect 26470 11820 26486 11837
rect 27328 11837 28144 11853
rect 27328 11820 27344 11837
rect 26470 11803 26878 11820
rect 25278 11756 26878 11803
rect 26936 11803 27344 11820
rect 28128 11820 28144 11837
rect 28986 11837 29802 11853
rect 28986 11820 29002 11837
rect 28128 11803 28536 11820
rect 26936 11756 28536 11803
rect 28594 11803 29002 11820
rect 29786 11820 29802 11837
rect 30644 11837 31460 11853
rect 30644 11820 30660 11837
rect 29786 11803 30194 11820
rect 28594 11756 30194 11803
rect 30252 11803 30660 11820
rect 31444 11820 31460 11837
rect 32302 11837 33118 11853
rect 32302 11820 32318 11837
rect 31444 11803 31852 11820
rect 30252 11756 31852 11803
rect 31910 11803 32318 11820
rect 33102 11820 33118 11837
rect 33102 11803 33510 11820
rect 31910 11756 33510 11803
rect -32752 10309 -31152 10356
rect -32752 10292 -32344 10309
rect -32360 10275 -32344 10292
rect -31560 10292 -31152 10309
rect -31094 10309 -29494 10356
rect -31094 10292 -30686 10309
rect -31560 10275 -31544 10292
rect -32360 10259 -31544 10275
rect -30702 10275 -30686 10292
rect -29902 10292 -29494 10309
rect -29436 10309 -27836 10356
rect -29436 10292 -29028 10309
rect -29902 10275 -29886 10292
rect -30702 10259 -29886 10275
rect -29044 10275 -29028 10292
rect -28244 10292 -27836 10309
rect -27778 10309 -26178 10356
rect -27778 10292 -27370 10309
rect -28244 10275 -28228 10292
rect -29044 10259 -28228 10275
rect -27386 10275 -27370 10292
rect -26586 10292 -26178 10309
rect -26120 10309 -24520 10356
rect -26120 10292 -25712 10309
rect -26586 10275 -26570 10292
rect -27386 10259 -26570 10275
rect -25728 10275 -25712 10292
rect -24928 10292 -24520 10309
rect -24462 10309 -22862 10356
rect -24462 10292 -24054 10309
rect -24928 10275 -24912 10292
rect -25728 10259 -24912 10275
rect -24070 10275 -24054 10292
rect -23270 10292 -22862 10309
rect -22804 10309 -21204 10356
rect -22804 10292 -22396 10309
rect -23270 10275 -23254 10292
rect -24070 10259 -23254 10275
rect -22412 10275 -22396 10292
rect -21612 10292 -21204 10309
rect -21146 10309 -19546 10356
rect -21146 10292 -20738 10309
rect -21612 10275 -21596 10292
rect -22412 10259 -21596 10275
rect -20754 10275 -20738 10292
rect -19954 10292 -19546 10309
rect -19488 10309 -17888 10356
rect -19488 10292 -19080 10309
rect -19954 10275 -19938 10292
rect -20754 10259 -19938 10275
rect -19096 10275 -19080 10292
rect -18296 10292 -17888 10309
rect -17830 10309 -16230 10356
rect -17830 10292 -17422 10309
rect -18296 10275 -18280 10292
rect -19096 10259 -18280 10275
rect -17438 10275 -17422 10292
rect -16638 10292 -16230 10309
rect -16172 10309 -14572 10356
rect -16172 10292 -15764 10309
rect -16638 10275 -16622 10292
rect -17438 10259 -16622 10275
rect -15780 10275 -15764 10292
rect -14980 10292 -14572 10309
rect -14514 10309 -12914 10356
rect -14514 10292 -14106 10309
rect -14980 10275 -14964 10292
rect -15780 10259 -14964 10275
rect -14122 10275 -14106 10292
rect -13322 10292 -12914 10309
rect -12856 10309 -11256 10356
rect -12856 10292 -12448 10309
rect -13322 10275 -13306 10292
rect -14122 10259 -13306 10275
rect -12464 10275 -12448 10292
rect -11664 10292 -11256 10309
rect -11198 10309 -9598 10356
rect -11198 10292 -10790 10309
rect -11664 10275 -11648 10292
rect -12464 10259 -11648 10275
rect -10806 10275 -10790 10292
rect -10006 10292 -9598 10309
rect -9540 10309 -7940 10356
rect -9540 10292 -9132 10309
rect -10006 10275 -9990 10292
rect -10806 10259 -9990 10275
rect -9148 10275 -9132 10292
rect -8348 10292 -7940 10309
rect -7882 10309 -6282 10356
rect -7882 10292 -7474 10309
rect -8348 10275 -8332 10292
rect -9148 10259 -8332 10275
rect -7490 10275 -7474 10292
rect -6690 10292 -6282 10309
rect -6224 10309 -4624 10356
rect -6224 10292 -5816 10309
rect -6690 10275 -6674 10292
rect -7490 10259 -6674 10275
rect -5832 10275 -5816 10292
rect -5032 10292 -4624 10309
rect -4566 10309 -2966 10356
rect -4566 10292 -4158 10309
rect -5032 10275 -5016 10292
rect -5832 10259 -5016 10275
rect -4174 10275 -4158 10292
rect -3374 10292 -2966 10309
rect -2908 10309 -1308 10356
rect -2908 10292 -2500 10309
rect -3374 10275 -3358 10292
rect -4174 10259 -3358 10275
rect -2516 10275 -2500 10292
rect -1716 10292 -1308 10309
rect -1250 10309 350 10356
rect -1250 10292 -842 10309
rect -1716 10275 -1700 10292
rect -2516 10259 -1700 10275
rect -858 10275 -842 10292
rect -58 10292 350 10309
rect 408 10309 2008 10356
rect 408 10292 816 10309
rect -58 10275 -42 10292
rect -858 10259 -42 10275
rect 800 10275 816 10292
rect 1600 10292 2008 10309
rect 2066 10309 3666 10356
rect 2066 10292 2474 10309
rect 1600 10275 1616 10292
rect 800 10259 1616 10275
rect 2458 10275 2474 10292
rect 3258 10292 3666 10309
rect 3724 10309 5324 10356
rect 3724 10292 4132 10309
rect 3258 10275 3274 10292
rect 2458 10259 3274 10275
rect 4116 10275 4132 10292
rect 4916 10292 5324 10309
rect 5382 10309 6982 10356
rect 5382 10292 5790 10309
rect 4916 10275 4932 10292
rect 4116 10259 4932 10275
rect 5774 10275 5790 10292
rect 6574 10292 6982 10309
rect 7040 10309 8640 10356
rect 7040 10292 7448 10309
rect 6574 10275 6590 10292
rect 5774 10259 6590 10275
rect 7432 10275 7448 10292
rect 8232 10292 8640 10309
rect 8698 10309 10298 10356
rect 8698 10292 9106 10309
rect 8232 10275 8248 10292
rect 7432 10259 8248 10275
rect 9090 10275 9106 10292
rect 9890 10292 10298 10309
rect 10356 10309 11956 10356
rect 10356 10292 10764 10309
rect 9890 10275 9906 10292
rect 9090 10259 9906 10275
rect 10748 10275 10764 10292
rect 11548 10292 11956 10309
rect 12014 10309 13614 10356
rect 12014 10292 12422 10309
rect 11548 10275 11564 10292
rect 10748 10259 11564 10275
rect 12406 10275 12422 10292
rect 13206 10292 13614 10309
rect 13672 10309 15272 10356
rect 13672 10292 14080 10309
rect 13206 10275 13222 10292
rect 12406 10259 13222 10275
rect 14064 10275 14080 10292
rect 14864 10292 15272 10309
rect 15330 10309 16930 10356
rect 15330 10292 15738 10309
rect 14864 10275 14880 10292
rect 14064 10259 14880 10275
rect 15722 10275 15738 10292
rect 16522 10292 16930 10309
rect 16988 10309 18588 10356
rect 16988 10292 17396 10309
rect 16522 10275 16538 10292
rect 15722 10259 16538 10275
rect 17380 10275 17396 10292
rect 18180 10292 18588 10309
rect 18646 10309 20246 10356
rect 18646 10292 19054 10309
rect 18180 10275 18196 10292
rect 17380 10259 18196 10275
rect 19038 10275 19054 10292
rect 19838 10292 20246 10309
rect 20304 10309 21904 10356
rect 20304 10292 20712 10309
rect 19838 10275 19854 10292
rect 19038 10259 19854 10275
rect 20696 10275 20712 10292
rect 21496 10292 21904 10309
rect 21962 10309 23562 10356
rect 21962 10292 22370 10309
rect 21496 10275 21512 10292
rect 20696 10259 21512 10275
rect 22354 10275 22370 10292
rect 23154 10292 23562 10309
rect 23620 10309 25220 10356
rect 23620 10292 24028 10309
rect 23154 10275 23170 10292
rect 22354 10259 23170 10275
rect 24012 10275 24028 10292
rect 24812 10292 25220 10309
rect 25278 10309 26878 10356
rect 25278 10292 25686 10309
rect 24812 10275 24828 10292
rect 24012 10259 24828 10275
rect 25670 10275 25686 10292
rect 26470 10292 26878 10309
rect 26936 10309 28536 10356
rect 26936 10292 27344 10309
rect 26470 10275 26486 10292
rect 25670 10259 26486 10275
rect 27328 10275 27344 10292
rect 28128 10292 28536 10309
rect 28594 10309 30194 10356
rect 28594 10292 29002 10309
rect 28128 10275 28144 10292
rect 27328 10259 28144 10275
rect 28986 10275 29002 10292
rect 29786 10292 30194 10309
rect 30252 10309 31852 10356
rect 30252 10292 30660 10309
rect 29786 10275 29802 10292
rect 28986 10259 29802 10275
rect 30644 10275 30660 10292
rect 31444 10292 31852 10309
rect 31910 10309 33510 10356
rect 31910 10292 32318 10309
rect 31444 10275 31460 10292
rect 30644 10259 31460 10275
rect 32302 10275 32318 10292
rect 33102 10292 33510 10309
rect 33102 10275 33118 10292
rect 32302 10259 33118 10275
rect -32360 10201 -31544 10217
rect -32360 10184 -32344 10201
rect -32752 10167 -32344 10184
rect -31560 10184 -31544 10201
rect -30702 10201 -29886 10217
rect -30702 10184 -30686 10201
rect -31560 10167 -31152 10184
rect -32752 10120 -31152 10167
rect -31094 10167 -30686 10184
rect -29902 10184 -29886 10201
rect -29044 10201 -28228 10217
rect -29044 10184 -29028 10201
rect -29902 10167 -29494 10184
rect -31094 10120 -29494 10167
rect -29436 10167 -29028 10184
rect -28244 10184 -28228 10201
rect -27386 10201 -26570 10217
rect -27386 10184 -27370 10201
rect -28244 10167 -27836 10184
rect -29436 10120 -27836 10167
rect -27778 10167 -27370 10184
rect -26586 10184 -26570 10201
rect -25728 10201 -24912 10217
rect -25728 10184 -25712 10201
rect -26586 10167 -26178 10184
rect -27778 10120 -26178 10167
rect -26120 10167 -25712 10184
rect -24928 10184 -24912 10201
rect -24070 10201 -23254 10217
rect -24070 10184 -24054 10201
rect -24928 10167 -24520 10184
rect -26120 10120 -24520 10167
rect -24462 10167 -24054 10184
rect -23270 10184 -23254 10201
rect -22412 10201 -21596 10217
rect -22412 10184 -22396 10201
rect -23270 10167 -22862 10184
rect -24462 10120 -22862 10167
rect -22804 10167 -22396 10184
rect -21612 10184 -21596 10201
rect -20754 10201 -19938 10217
rect -20754 10184 -20738 10201
rect -21612 10167 -21204 10184
rect -22804 10120 -21204 10167
rect -21146 10167 -20738 10184
rect -19954 10184 -19938 10201
rect -19096 10201 -18280 10217
rect -19096 10184 -19080 10201
rect -19954 10167 -19546 10184
rect -21146 10120 -19546 10167
rect -19488 10167 -19080 10184
rect -18296 10184 -18280 10201
rect -17438 10201 -16622 10217
rect -17438 10184 -17422 10201
rect -18296 10167 -17888 10184
rect -19488 10120 -17888 10167
rect -17830 10167 -17422 10184
rect -16638 10184 -16622 10201
rect -15780 10201 -14964 10217
rect -15780 10184 -15764 10201
rect -16638 10167 -16230 10184
rect -17830 10120 -16230 10167
rect -16172 10167 -15764 10184
rect -14980 10184 -14964 10201
rect -14122 10201 -13306 10217
rect -14122 10184 -14106 10201
rect -14980 10167 -14572 10184
rect -16172 10120 -14572 10167
rect -14514 10167 -14106 10184
rect -13322 10184 -13306 10201
rect -12464 10201 -11648 10217
rect -12464 10184 -12448 10201
rect -13322 10167 -12914 10184
rect -14514 10120 -12914 10167
rect -12856 10167 -12448 10184
rect -11664 10184 -11648 10201
rect -10806 10201 -9990 10217
rect -10806 10184 -10790 10201
rect -11664 10167 -11256 10184
rect -12856 10120 -11256 10167
rect -11198 10167 -10790 10184
rect -10006 10184 -9990 10201
rect -9148 10201 -8332 10217
rect -9148 10184 -9132 10201
rect -10006 10167 -9598 10184
rect -11198 10120 -9598 10167
rect -9540 10167 -9132 10184
rect -8348 10184 -8332 10201
rect -7490 10201 -6674 10217
rect -7490 10184 -7474 10201
rect -8348 10167 -7940 10184
rect -9540 10120 -7940 10167
rect -7882 10167 -7474 10184
rect -6690 10184 -6674 10201
rect -5832 10201 -5016 10217
rect -5832 10184 -5816 10201
rect -6690 10167 -6282 10184
rect -7882 10120 -6282 10167
rect -6224 10167 -5816 10184
rect -5032 10184 -5016 10201
rect -4174 10201 -3358 10217
rect -4174 10184 -4158 10201
rect -5032 10167 -4624 10184
rect -6224 10120 -4624 10167
rect -4566 10167 -4158 10184
rect -3374 10184 -3358 10201
rect -2516 10201 -1700 10217
rect -2516 10184 -2500 10201
rect -3374 10167 -2966 10184
rect -4566 10120 -2966 10167
rect -2908 10167 -2500 10184
rect -1716 10184 -1700 10201
rect -858 10201 -42 10217
rect -858 10184 -842 10201
rect -1716 10167 -1308 10184
rect -2908 10120 -1308 10167
rect -1250 10167 -842 10184
rect -58 10184 -42 10201
rect 800 10201 1616 10217
rect 800 10184 816 10201
rect -58 10167 350 10184
rect -1250 10120 350 10167
rect 408 10167 816 10184
rect 1600 10184 1616 10201
rect 2458 10201 3274 10217
rect 2458 10184 2474 10201
rect 1600 10167 2008 10184
rect 408 10120 2008 10167
rect 2066 10167 2474 10184
rect 3258 10184 3274 10201
rect 4116 10201 4932 10217
rect 4116 10184 4132 10201
rect 3258 10167 3666 10184
rect 2066 10120 3666 10167
rect 3724 10167 4132 10184
rect 4916 10184 4932 10201
rect 5774 10201 6590 10217
rect 5774 10184 5790 10201
rect 4916 10167 5324 10184
rect 3724 10120 5324 10167
rect 5382 10167 5790 10184
rect 6574 10184 6590 10201
rect 7432 10201 8248 10217
rect 7432 10184 7448 10201
rect 6574 10167 6982 10184
rect 5382 10120 6982 10167
rect 7040 10167 7448 10184
rect 8232 10184 8248 10201
rect 9090 10201 9906 10217
rect 9090 10184 9106 10201
rect 8232 10167 8640 10184
rect 7040 10120 8640 10167
rect 8698 10167 9106 10184
rect 9890 10184 9906 10201
rect 10748 10201 11564 10217
rect 10748 10184 10764 10201
rect 9890 10167 10298 10184
rect 8698 10120 10298 10167
rect 10356 10167 10764 10184
rect 11548 10184 11564 10201
rect 12406 10201 13222 10217
rect 12406 10184 12422 10201
rect 11548 10167 11956 10184
rect 10356 10120 11956 10167
rect 12014 10167 12422 10184
rect 13206 10184 13222 10201
rect 14064 10201 14880 10217
rect 14064 10184 14080 10201
rect 13206 10167 13614 10184
rect 12014 10120 13614 10167
rect 13672 10167 14080 10184
rect 14864 10184 14880 10201
rect 15722 10201 16538 10217
rect 15722 10184 15738 10201
rect 14864 10167 15272 10184
rect 13672 10120 15272 10167
rect 15330 10167 15738 10184
rect 16522 10184 16538 10201
rect 17380 10201 18196 10217
rect 17380 10184 17396 10201
rect 16522 10167 16930 10184
rect 15330 10120 16930 10167
rect 16988 10167 17396 10184
rect 18180 10184 18196 10201
rect 19038 10201 19854 10217
rect 19038 10184 19054 10201
rect 18180 10167 18588 10184
rect 16988 10120 18588 10167
rect 18646 10167 19054 10184
rect 19838 10184 19854 10201
rect 20696 10201 21512 10217
rect 20696 10184 20712 10201
rect 19838 10167 20246 10184
rect 18646 10120 20246 10167
rect 20304 10167 20712 10184
rect 21496 10184 21512 10201
rect 22354 10201 23170 10217
rect 22354 10184 22370 10201
rect 21496 10167 21904 10184
rect 20304 10120 21904 10167
rect 21962 10167 22370 10184
rect 23154 10184 23170 10201
rect 24012 10201 24828 10217
rect 24012 10184 24028 10201
rect 23154 10167 23562 10184
rect 21962 10120 23562 10167
rect 23620 10167 24028 10184
rect 24812 10184 24828 10201
rect 25670 10201 26486 10217
rect 25670 10184 25686 10201
rect 24812 10167 25220 10184
rect 23620 10120 25220 10167
rect 25278 10167 25686 10184
rect 26470 10184 26486 10201
rect 27328 10201 28144 10217
rect 27328 10184 27344 10201
rect 26470 10167 26878 10184
rect 25278 10120 26878 10167
rect 26936 10167 27344 10184
rect 28128 10184 28144 10201
rect 28986 10201 29802 10217
rect 28986 10184 29002 10201
rect 28128 10167 28536 10184
rect 26936 10120 28536 10167
rect 28594 10167 29002 10184
rect 29786 10184 29802 10201
rect 30644 10201 31460 10217
rect 30644 10184 30660 10201
rect 29786 10167 30194 10184
rect 28594 10120 30194 10167
rect 30252 10167 30660 10184
rect 31444 10184 31460 10201
rect 32302 10201 33118 10217
rect 32302 10184 32318 10201
rect 31444 10167 31852 10184
rect 30252 10120 31852 10167
rect 31910 10167 32318 10184
rect 33102 10184 33118 10201
rect 33102 10167 33510 10184
rect 31910 10120 33510 10167
rect -32752 8673 -31152 8720
rect -32752 8656 -32344 8673
rect -32360 8639 -32344 8656
rect -31560 8656 -31152 8673
rect -31094 8673 -29494 8720
rect -31094 8656 -30686 8673
rect -31560 8639 -31544 8656
rect -32360 8623 -31544 8639
rect -30702 8639 -30686 8656
rect -29902 8656 -29494 8673
rect -29436 8673 -27836 8720
rect -29436 8656 -29028 8673
rect -29902 8639 -29886 8656
rect -30702 8623 -29886 8639
rect -29044 8639 -29028 8656
rect -28244 8656 -27836 8673
rect -27778 8673 -26178 8720
rect -27778 8656 -27370 8673
rect -28244 8639 -28228 8656
rect -29044 8623 -28228 8639
rect -27386 8639 -27370 8656
rect -26586 8656 -26178 8673
rect -26120 8673 -24520 8720
rect -26120 8656 -25712 8673
rect -26586 8639 -26570 8656
rect -27386 8623 -26570 8639
rect -25728 8639 -25712 8656
rect -24928 8656 -24520 8673
rect -24462 8673 -22862 8720
rect -24462 8656 -24054 8673
rect -24928 8639 -24912 8656
rect -25728 8623 -24912 8639
rect -24070 8639 -24054 8656
rect -23270 8656 -22862 8673
rect -22804 8673 -21204 8720
rect -22804 8656 -22396 8673
rect -23270 8639 -23254 8656
rect -24070 8623 -23254 8639
rect -22412 8639 -22396 8656
rect -21612 8656 -21204 8673
rect -21146 8673 -19546 8720
rect -21146 8656 -20738 8673
rect -21612 8639 -21596 8656
rect -22412 8623 -21596 8639
rect -20754 8639 -20738 8656
rect -19954 8656 -19546 8673
rect -19488 8673 -17888 8720
rect -19488 8656 -19080 8673
rect -19954 8639 -19938 8656
rect -20754 8623 -19938 8639
rect -19096 8639 -19080 8656
rect -18296 8656 -17888 8673
rect -17830 8673 -16230 8720
rect -17830 8656 -17422 8673
rect -18296 8639 -18280 8656
rect -19096 8623 -18280 8639
rect -17438 8639 -17422 8656
rect -16638 8656 -16230 8673
rect -16172 8673 -14572 8720
rect -16172 8656 -15764 8673
rect -16638 8639 -16622 8656
rect -17438 8623 -16622 8639
rect -15780 8639 -15764 8656
rect -14980 8656 -14572 8673
rect -14514 8673 -12914 8720
rect -14514 8656 -14106 8673
rect -14980 8639 -14964 8656
rect -15780 8623 -14964 8639
rect -14122 8639 -14106 8656
rect -13322 8656 -12914 8673
rect -12856 8673 -11256 8720
rect -12856 8656 -12448 8673
rect -13322 8639 -13306 8656
rect -14122 8623 -13306 8639
rect -12464 8639 -12448 8656
rect -11664 8656 -11256 8673
rect -11198 8673 -9598 8720
rect -11198 8656 -10790 8673
rect -11664 8639 -11648 8656
rect -12464 8623 -11648 8639
rect -10806 8639 -10790 8656
rect -10006 8656 -9598 8673
rect -9540 8673 -7940 8720
rect -9540 8656 -9132 8673
rect -10006 8639 -9990 8656
rect -10806 8623 -9990 8639
rect -9148 8639 -9132 8656
rect -8348 8656 -7940 8673
rect -7882 8673 -6282 8720
rect -7882 8656 -7474 8673
rect -8348 8639 -8332 8656
rect -9148 8623 -8332 8639
rect -7490 8639 -7474 8656
rect -6690 8656 -6282 8673
rect -6224 8673 -4624 8720
rect -6224 8656 -5816 8673
rect -6690 8639 -6674 8656
rect -7490 8623 -6674 8639
rect -5832 8639 -5816 8656
rect -5032 8656 -4624 8673
rect -4566 8673 -2966 8720
rect -4566 8656 -4158 8673
rect -5032 8639 -5016 8656
rect -5832 8623 -5016 8639
rect -4174 8639 -4158 8656
rect -3374 8656 -2966 8673
rect -2908 8673 -1308 8720
rect -2908 8656 -2500 8673
rect -3374 8639 -3358 8656
rect -4174 8623 -3358 8639
rect -2516 8639 -2500 8656
rect -1716 8656 -1308 8673
rect -1250 8673 350 8720
rect -1250 8656 -842 8673
rect -1716 8639 -1700 8656
rect -2516 8623 -1700 8639
rect -858 8639 -842 8656
rect -58 8656 350 8673
rect 408 8673 2008 8720
rect 408 8656 816 8673
rect -58 8639 -42 8656
rect -858 8623 -42 8639
rect 800 8639 816 8656
rect 1600 8656 2008 8673
rect 2066 8673 3666 8720
rect 2066 8656 2474 8673
rect 1600 8639 1616 8656
rect 800 8623 1616 8639
rect 2458 8639 2474 8656
rect 3258 8656 3666 8673
rect 3724 8673 5324 8720
rect 3724 8656 4132 8673
rect 3258 8639 3274 8656
rect 2458 8623 3274 8639
rect 4116 8639 4132 8656
rect 4916 8656 5324 8673
rect 5382 8673 6982 8720
rect 5382 8656 5790 8673
rect 4916 8639 4932 8656
rect 4116 8623 4932 8639
rect 5774 8639 5790 8656
rect 6574 8656 6982 8673
rect 7040 8673 8640 8720
rect 7040 8656 7448 8673
rect 6574 8639 6590 8656
rect 5774 8623 6590 8639
rect 7432 8639 7448 8656
rect 8232 8656 8640 8673
rect 8698 8673 10298 8720
rect 8698 8656 9106 8673
rect 8232 8639 8248 8656
rect 7432 8623 8248 8639
rect 9090 8639 9106 8656
rect 9890 8656 10298 8673
rect 10356 8673 11956 8720
rect 10356 8656 10764 8673
rect 9890 8639 9906 8656
rect 9090 8623 9906 8639
rect 10748 8639 10764 8656
rect 11548 8656 11956 8673
rect 12014 8673 13614 8720
rect 12014 8656 12422 8673
rect 11548 8639 11564 8656
rect 10748 8623 11564 8639
rect 12406 8639 12422 8656
rect 13206 8656 13614 8673
rect 13672 8673 15272 8720
rect 13672 8656 14080 8673
rect 13206 8639 13222 8656
rect 12406 8623 13222 8639
rect 14064 8639 14080 8656
rect 14864 8656 15272 8673
rect 15330 8673 16930 8720
rect 15330 8656 15738 8673
rect 14864 8639 14880 8656
rect 14064 8623 14880 8639
rect 15722 8639 15738 8656
rect 16522 8656 16930 8673
rect 16988 8673 18588 8720
rect 16988 8656 17396 8673
rect 16522 8639 16538 8656
rect 15722 8623 16538 8639
rect 17380 8639 17396 8656
rect 18180 8656 18588 8673
rect 18646 8673 20246 8720
rect 18646 8656 19054 8673
rect 18180 8639 18196 8656
rect 17380 8623 18196 8639
rect 19038 8639 19054 8656
rect 19838 8656 20246 8673
rect 20304 8673 21904 8720
rect 20304 8656 20712 8673
rect 19838 8639 19854 8656
rect 19038 8623 19854 8639
rect 20696 8639 20712 8656
rect 21496 8656 21904 8673
rect 21962 8673 23562 8720
rect 21962 8656 22370 8673
rect 21496 8639 21512 8656
rect 20696 8623 21512 8639
rect 22354 8639 22370 8656
rect 23154 8656 23562 8673
rect 23620 8673 25220 8720
rect 23620 8656 24028 8673
rect 23154 8639 23170 8656
rect 22354 8623 23170 8639
rect 24012 8639 24028 8656
rect 24812 8656 25220 8673
rect 25278 8673 26878 8720
rect 25278 8656 25686 8673
rect 24812 8639 24828 8656
rect 24012 8623 24828 8639
rect 25670 8639 25686 8656
rect 26470 8656 26878 8673
rect 26936 8673 28536 8720
rect 26936 8656 27344 8673
rect 26470 8639 26486 8656
rect 25670 8623 26486 8639
rect 27328 8639 27344 8656
rect 28128 8656 28536 8673
rect 28594 8673 30194 8720
rect 28594 8656 29002 8673
rect 28128 8639 28144 8656
rect 27328 8623 28144 8639
rect 28986 8639 29002 8656
rect 29786 8656 30194 8673
rect 30252 8673 31852 8720
rect 30252 8656 30660 8673
rect 29786 8639 29802 8656
rect 28986 8623 29802 8639
rect 30644 8639 30660 8656
rect 31444 8656 31852 8673
rect 31910 8673 33510 8720
rect 31910 8656 32318 8673
rect 31444 8639 31460 8656
rect 30644 8623 31460 8639
rect 32302 8639 32318 8656
rect 33102 8656 33510 8673
rect 33102 8639 33118 8656
rect 32302 8623 33118 8639
rect -32360 8565 -31544 8581
rect -32360 8548 -32344 8565
rect -32752 8531 -32344 8548
rect -31560 8548 -31544 8565
rect -30702 8565 -29886 8581
rect -30702 8548 -30686 8565
rect -31560 8531 -31152 8548
rect -32752 8484 -31152 8531
rect -31094 8531 -30686 8548
rect -29902 8548 -29886 8565
rect -29044 8565 -28228 8581
rect -29044 8548 -29028 8565
rect -29902 8531 -29494 8548
rect -31094 8484 -29494 8531
rect -29436 8531 -29028 8548
rect -28244 8548 -28228 8565
rect -27386 8565 -26570 8581
rect -27386 8548 -27370 8565
rect -28244 8531 -27836 8548
rect -29436 8484 -27836 8531
rect -27778 8531 -27370 8548
rect -26586 8548 -26570 8565
rect -25728 8565 -24912 8581
rect -25728 8548 -25712 8565
rect -26586 8531 -26178 8548
rect -27778 8484 -26178 8531
rect -26120 8531 -25712 8548
rect -24928 8548 -24912 8565
rect -24070 8565 -23254 8581
rect -24070 8548 -24054 8565
rect -24928 8531 -24520 8548
rect -26120 8484 -24520 8531
rect -24462 8531 -24054 8548
rect -23270 8548 -23254 8565
rect -22412 8565 -21596 8581
rect -22412 8548 -22396 8565
rect -23270 8531 -22862 8548
rect -24462 8484 -22862 8531
rect -22804 8531 -22396 8548
rect -21612 8548 -21596 8565
rect -20754 8565 -19938 8581
rect -20754 8548 -20738 8565
rect -21612 8531 -21204 8548
rect -22804 8484 -21204 8531
rect -21146 8531 -20738 8548
rect -19954 8548 -19938 8565
rect -19096 8565 -18280 8581
rect -19096 8548 -19080 8565
rect -19954 8531 -19546 8548
rect -21146 8484 -19546 8531
rect -19488 8531 -19080 8548
rect -18296 8548 -18280 8565
rect -17438 8565 -16622 8581
rect -17438 8548 -17422 8565
rect -18296 8531 -17888 8548
rect -19488 8484 -17888 8531
rect -17830 8531 -17422 8548
rect -16638 8548 -16622 8565
rect -15780 8565 -14964 8581
rect -15780 8548 -15764 8565
rect -16638 8531 -16230 8548
rect -17830 8484 -16230 8531
rect -16172 8531 -15764 8548
rect -14980 8548 -14964 8565
rect -14122 8565 -13306 8581
rect -14122 8548 -14106 8565
rect -14980 8531 -14572 8548
rect -16172 8484 -14572 8531
rect -14514 8531 -14106 8548
rect -13322 8548 -13306 8565
rect -12464 8565 -11648 8581
rect -12464 8548 -12448 8565
rect -13322 8531 -12914 8548
rect -14514 8484 -12914 8531
rect -12856 8531 -12448 8548
rect -11664 8548 -11648 8565
rect -10806 8565 -9990 8581
rect -10806 8548 -10790 8565
rect -11664 8531 -11256 8548
rect -12856 8484 -11256 8531
rect -11198 8531 -10790 8548
rect -10006 8548 -9990 8565
rect -9148 8565 -8332 8581
rect -9148 8548 -9132 8565
rect -10006 8531 -9598 8548
rect -11198 8484 -9598 8531
rect -9540 8531 -9132 8548
rect -8348 8548 -8332 8565
rect -7490 8565 -6674 8581
rect -7490 8548 -7474 8565
rect -8348 8531 -7940 8548
rect -9540 8484 -7940 8531
rect -7882 8531 -7474 8548
rect -6690 8548 -6674 8565
rect -5832 8565 -5016 8581
rect -5832 8548 -5816 8565
rect -6690 8531 -6282 8548
rect -7882 8484 -6282 8531
rect -6224 8531 -5816 8548
rect -5032 8548 -5016 8565
rect -4174 8565 -3358 8581
rect -4174 8548 -4158 8565
rect -5032 8531 -4624 8548
rect -6224 8484 -4624 8531
rect -4566 8531 -4158 8548
rect -3374 8548 -3358 8565
rect -2516 8565 -1700 8581
rect -2516 8548 -2500 8565
rect -3374 8531 -2966 8548
rect -4566 8484 -2966 8531
rect -2908 8531 -2500 8548
rect -1716 8548 -1700 8565
rect -858 8565 -42 8581
rect -858 8548 -842 8565
rect -1716 8531 -1308 8548
rect -2908 8484 -1308 8531
rect -1250 8531 -842 8548
rect -58 8548 -42 8565
rect 800 8565 1616 8581
rect 800 8548 816 8565
rect -58 8531 350 8548
rect -1250 8484 350 8531
rect 408 8531 816 8548
rect 1600 8548 1616 8565
rect 2458 8565 3274 8581
rect 2458 8548 2474 8565
rect 1600 8531 2008 8548
rect 408 8484 2008 8531
rect 2066 8531 2474 8548
rect 3258 8548 3274 8565
rect 4116 8565 4932 8581
rect 4116 8548 4132 8565
rect 3258 8531 3666 8548
rect 2066 8484 3666 8531
rect 3724 8531 4132 8548
rect 4916 8548 4932 8565
rect 5774 8565 6590 8581
rect 5774 8548 5790 8565
rect 4916 8531 5324 8548
rect 3724 8484 5324 8531
rect 5382 8531 5790 8548
rect 6574 8548 6590 8565
rect 7432 8565 8248 8581
rect 7432 8548 7448 8565
rect 6574 8531 6982 8548
rect 5382 8484 6982 8531
rect 7040 8531 7448 8548
rect 8232 8548 8248 8565
rect 9090 8565 9906 8581
rect 9090 8548 9106 8565
rect 8232 8531 8640 8548
rect 7040 8484 8640 8531
rect 8698 8531 9106 8548
rect 9890 8548 9906 8565
rect 10748 8565 11564 8581
rect 10748 8548 10764 8565
rect 9890 8531 10298 8548
rect 8698 8484 10298 8531
rect 10356 8531 10764 8548
rect 11548 8548 11564 8565
rect 12406 8565 13222 8581
rect 12406 8548 12422 8565
rect 11548 8531 11956 8548
rect 10356 8484 11956 8531
rect 12014 8531 12422 8548
rect 13206 8548 13222 8565
rect 14064 8565 14880 8581
rect 14064 8548 14080 8565
rect 13206 8531 13614 8548
rect 12014 8484 13614 8531
rect 13672 8531 14080 8548
rect 14864 8548 14880 8565
rect 15722 8565 16538 8581
rect 15722 8548 15738 8565
rect 14864 8531 15272 8548
rect 13672 8484 15272 8531
rect 15330 8531 15738 8548
rect 16522 8548 16538 8565
rect 17380 8565 18196 8581
rect 17380 8548 17396 8565
rect 16522 8531 16930 8548
rect 15330 8484 16930 8531
rect 16988 8531 17396 8548
rect 18180 8548 18196 8565
rect 19038 8565 19854 8581
rect 19038 8548 19054 8565
rect 18180 8531 18588 8548
rect 16988 8484 18588 8531
rect 18646 8531 19054 8548
rect 19838 8548 19854 8565
rect 20696 8565 21512 8581
rect 20696 8548 20712 8565
rect 19838 8531 20246 8548
rect 18646 8484 20246 8531
rect 20304 8531 20712 8548
rect 21496 8548 21512 8565
rect 22354 8565 23170 8581
rect 22354 8548 22370 8565
rect 21496 8531 21904 8548
rect 20304 8484 21904 8531
rect 21962 8531 22370 8548
rect 23154 8548 23170 8565
rect 24012 8565 24828 8581
rect 24012 8548 24028 8565
rect 23154 8531 23562 8548
rect 21962 8484 23562 8531
rect 23620 8531 24028 8548
rect 24812 8548 24828 8565
rect 25670 8565 26486 8581
rect 25670 8548 25686 8565
rect 24812 8531 25220 8548
rect 23620 8484 25220 8531
rect 25278 8531 25686 8548
rect 26470 8548 26486 8565
rect 27328 8565 28144 8581
rect 27328 8548 27344 8565
rect 26470 8531 26878 8548
rect 25278 8484 26878 8531
rect 26936 8531 27344 8548
rect 28128 8548 28144 8565
rect 28986 8565 29802 8581
rect 28986 8548 29002 8565
rect 28128 8531 28536 8548
rect 26936 8484 28536 8531
rect 28594 8531 29002 8548
rect 29786 8548 29802 8565
rect 30644 8565 31460 8581
rect 30644 8548 30660 8565
rect 29786 8531 30194 8548
rect 28594 8484 30194 8531
rect 30252 8531 30660 8548
rect 31444 8548 31460 8565
rect 32302 8565 33118 8581
rect 32302 8548 32318 8565
rect 31444 8531 31852 8548
rect 30252 8484 31852 8531
rect 31910 8531 32318 8548
rect 33102 8548 33118 8565
rect 33102 8531 33510 8548
rect 31910 8484 33510 8531
rect -32752 7037 -31152 7084
rect -32752 7020 -32344 7037
rect -32360 7003 -32344 7020
rect -31560 7020 -31152 7037
rect -31094 7037 -29494 7084
rect -31094 7020 -30686 7037
rect -31560 7003 -31544 7020
rect -32360 6987 -31544 7003
rect -30702 7003 -30686 7020
rect -29902 7020 -29494 7037
rect -29436 7037 -27836 7084
rect -29436 7020 -29028 7037
rect -29902 7003 -29886 7020
rect -30702 6987 -29886 7003
rect -29044 7003 -29028 7020
rect -28244 7020 -27836 7037
rect -27778 7037 -26178 7084
rect -27778 7020 -27370 7037
rect -28244 7003 -28228 7020
rect -29044 6987 -28228 7003
rect -27386 7003 -27370 7020
rect -26586 7020 -26178 7037
rect -26120 7037 -24520 7084
rect -26120 7020 -25712 7037
rect -26586 7003 -26570 7020
rect -27386 6987 -26570 7003
rect -25728 7003 -25712 7020
rect -24928 7020 -24520 7037
rect -24462 7037 -22862 7084
rect -24462 7020 -24054 7037
rect -24928 7003 -24912 7020
rect -25728 6987 -24912 7003
rect -24070 7003 -24054 7020
rect -23270 7020 -22862 7037
rect -22804 7037 -21204 7084
rect -22804 7020 -22396 7037
rect -23270 7003 -23254 7020
rect -24070 6987 -23254 7003
rect -22412 7003 -22396 7020
rect -21612 7020 -21204 7037
rect -21146 7037 -19546 7084
rect -21146 7020 -20738 7037
rect -21612 7003 -21596 7020
rect -22412 6987 -21596 7003
rect -20754 7003 -20738 7020
rect -19954 7020 -19546 7037
rect -19488 7037 -17888 7084
rect -19488 7020 -19080 7037
rect -19954 7003 -19938 7020
rect -20754 6987 -19938 7003
rect -19096 7003 -19080 7020
rect -18296 7020 -17888 7037
rect -17830 7037 -16230 7084
rect -17830 7020 -17422 7037
rect -18296 7003 -18280 7020
rect -19096 6987 -18280 7003
rect -17438 7003 -17422 7020
rect -16638 7020 -16230 7037
rect -16172 7037 -14572 7084
rect -16172 7020 -15764 7037
rect -16638 7003 -16622 7020
rect -17438 6987 -16622 7003
rect -15780 7003 -15764 7020
rect -14980 7020 -14572 7037
rect -14514 7037 -12914 7084
rect -14514 7020 -14106 7037
rect -14980 7003 -14964 7020
rect -15780 6987 -14964 7003
rect -14122 7003 -14106 7020
rect -13322 7020 -12914 7037
rect -12856 7037 -11256 7084
rect -12856 7020 -12448 7037
rect -13322 7003 -13306 7020
rect -14122 6987 -13306 7003
rect -12464 7003 -12448 7020
rect -11664 7020 -11256 7037
rect -11198 7037 -9598 7084
rect -11198 7020 -10790 7037
rect -11664 7003 -11648 7020
rect -12464 6987 -11648 7003
rect -10806 7003 -10790 7020
rect -10006 7020 -9598 7037
rect -9540 7037 -7940 7084
rect -9540 7020 -9132 7037
rect -10006 7003 -9990 7020
rect -10806 6987 -9990 7003
rect -9148 7003 -9132 7020
rect -8348 7020 -7940 7037
rect -7882 7037 -6282 7084
rect -7882 7020 -7474 7037
rect -8348 7003 -8332 7020
rect -9148 6987 -8332 7003
rect -7490 7003 -7474 7020
rect -6690 7020 -6282 7037
rect -6224 7037 -4624 7084
rect -6224 7020 -5816 7037
rect -6690 7003 -6674 7020
rect -7490 6987 -6674 7003
rect -5832 7003 -5816 7020
rect -5032 7020 -4624 7037
rect -4566 7037 -2966 7084
rect -4566 7020 -4158 7037
rect -5032 7003 -5016 7020
rect -5832 6987 -5016 7003
rect -4174 7003 -4158 7020
rect -3374 7020 -2966 7037
rect -2908 7037 -1308 7084
rect -2908 7020 -2500 7037
rect -3374 7003 -3358 7020
rect -4174 6987 -3358 7003
rect -2516 7003 -2500 7020
rect -1716 7020 -1308 7037
rect -1250 7037 350 7084
rect -1250 7020 -842 7037
rect -1716 7003 -1700 7020
rect -2516 6987 -1700 7003
rect -858 7003 -842 7020
rect -58 7020 350 7037
rect 408 7037 2008 7084
rect 408 7020 816 7037
rect -58 7003 -42 7020
rect -858 6987 -42 7003
rect 800 7003 816 7020
rect 1600 7020 2008 7037
rect 2066 7037 3666 7084
rect 2066 7020 2474 7037
rect 1600 7003 1616 7020
rect 800 6987 1616 7003
rect 2458 7003 2474 7020
rect 3258 7020 3666 7037
rect 3724 7037 5324 7084
rect 3724 7020 4132 7037
rect 3258 7003 3274 7020
rect 2458 6987 3274 7003
rect 4116 7003 4132 7020
rect 4916 7020 5324 7037
rect 5382 7037 6982 7084
rect 5382 7020 5790 7037
rect 4916 7003 4932 7020
rect 4116 6987 4932 7003
rect 5774 7003 5790 7020
rect 6574 7020 6982 7037
rect 7040 7037 8640 7084
rect 7040 7020 7448 7037
rect 6574 7003 6590 7020
rect 5774 6987 6590 7003
rect 7432 7003 7448 7020
rect 8232 7020 8640 7037
rect 8698 7037 10298 7084
rect 8698 7020 9106 7037
rect 8232 7003 8248 7020
rect 7432 6987 8248 7003
rect 9090 7003 9106 7020
rect 9890 7020 10298 7037
rect 10356 7037 11956 7084
rect 10356 7020 10764 7037
rect 9890 7003 9906 7020
rect 9090 6987 9906 7003
rect 10748 7003 10764 7020
rect 11548 7020 11956 7037
rect 12014 7037 13614 7084
rect 12014 7020 12422 7037
rect 11548 7003 11564 7020
rect 10748 6987 11564 7003
rect 12406 7003 12422 7020
rect 13206 7020 13614 7037
rect 13672 7037 15272 7084
rect 13672 7020 14080 7037
rect 13206 7003 13222 7020
rect 12406 6987 13222 7003
rect 14064 7003 14080 7020
rect 14864 7020 15272 7037
rect 15330 7037 16930 7084
rect 15330 7020 15738 7037
rect 14864 7003 14880 7020
rect 14064 6987 14880 7003
rect 15722 7003 15738 7020
rect 16522 7020 16930 7037
rect 16988 7037 18588 7084
rect 16988 7020 17396 7037
rect 16522 7003 16538 7020
rect 15722 6987 16538 7003
rect 17380 7003 17396 7020
rect 18180 7020 18588 7037
rect 18646 7037 20246 7084
rect 18646 7020 19054 7037
rect 18180 7003 18196 7020
rect 17380 6987 18196 7003
rect 19038 7003 19054 7020
rect 19838 7020 20246 7037
rect 20304 7037 21904 7084
rect 20304 7020 20712 7037
rect 19838 7003 19854 7020
rect 19038 6987 19854 7003
rect 20696 7003 20712 7020
rect 21496 7020 21904 7037
rect 21962 7037 23562 7084
rect 21962 7020 22370 7037
rect 21496 7003 21512 7020
rect 20696 6987 21512 7003
rect 22354 7003 22370 7020
rect 23154 7020 23562 7037
rect 23620 7037 25220 7084
rect 23620 7020 24028 7037
rect 23154 7003 23170 7020
rect 22354 6987 23170 7003
rect 24012 7003 24028 7020
rect 24812 7020 25220 7037
rect 25278 7037 26878 7084
rect 25278 7020 25686 7037
rect 24812 7003 24828 7020
rect 24012 6987 24828 7003
rect 25670 7003 25686 7020
rect 26470 7020 26878 7037
rect 26936 7037 28536 7084
rect 26936 7020 27344 7037
rect 26470 7003 26486 7020
rect 25670 6987 26486 7003
rect 27328 7003 27344 7020
rect 28128 7020 28536 7037
rect 28594 7037 30194 7084
rect 28594 7020 29002 7037
rect 28128 7003 28144 7020
rect 27328 6987 28144 7003
rect 28986 7003 29002 7020
rect 29786 7020 30194 7037
rect 30252 7037 31852 7084
rect 30252 7020 30660 7037
rect 29786 7003 29802 7020
rect 28986 6987 29802 7003
rect 30644 7003 30660 7020
rect 31444 7020 31852 7037
rect 31910 7037 33510 7084
rect 31910 7020 32318 7037
rect 31444 7003 31460 7020
rect 30644 6987 31460 7003
rect 32302 7003 32318 7020
rect 33102 7020 33510 7037
rect 33102 7003 33118 7020
rect 32302 6987 33118 7003
rect -32360 6927 -31544 6943
rect -32360 6910 -32344 6927
rect -32752 6893 -32344 6910
rect -31560 6910 -31544 6927
rect -30702 6927 -29886 6943
rect -30702 6910 -30686 6927
rect -31560 6893 -31152 6910
rect -32752 6846 -31152 6893
rect -31094 6893 -30686 6910
rect -29902 6910 -29886 6927
rect -29044 6927 -28228 6943
rect -29044 6910 -29028 6927
rect -29902 6893 -29494 6910
rect -31094 6846 -29494 6893
rect -29436 6893 -29028 6910
rect -28244 6910 -28228 6927
rect -27386 6927 -26570 6943
rect -27386 6910 -27370 6927
rect -28244 6893 -27836 6910
rect -29436 6846 -27836 6893
rect -27778 6893 -27370 6910
rect -26586 6910 -26570 6927
rect -25728 6927 -24912 6943
rect -25728 6910 -25712 6927
rect -26586 6893 -26178 6910
rect -27778 6846 -26178 6893
rect -26120 6893 -25712 6910
rect -24928 6910 -24912 6927
rect -24070 6927 -23254 6943
rect -24070 6910 -24054 6927
rect -24928 6893 -24520 6910
rect -26120 6846 -24520 6893
rect -24462 6893 -24054 6910
rect -23270 6910 -23254 6927
rect -22412 6927 -21596 6943
rect -22412 6910 -22396 6927
rect -23270 6893 -22862 6910
rect -24462 6846 -22862 6893
rect -22804 6893 -22396 6910
rect -21612 6910 -21596 6927
rect -20754 6927 -19938 6943
rect -20754 6910 -20738 6927
rect -21612 6893 -21204 6910
rect -22804 6846 -21204 6893
rect -21146 6893 -20738 6910
rect -19954 6910 -19938 6927
rect -19096 6927 -18280 6943
rect -19096 6910 -19080 6927
rect -19954 6893 -19546 6910
rect -21146 6846 -19546 6893
rect -19488 6893 -19080 6910
rect -18296 6910 -18280 6927
rect -17438 6927 -16622 6943
rect -17438 6910 -17422 6927
rect -18296 6893 -17888 6910
rect -19488 6846 -17888 6893
rect -17830 6893 -17422 6910
rect -16638 6910 -16622 6927
rect -15780 6927 -14964 6943
rect -15780 6910 -15764 6927
rect -16638 6893 -16230 6910
rect -17830 6846 -16230 6893
rect -16172 6893 -15764 6910
rect -14980 6910 -14964 6927
rect -14122 6927 -13306 6943
rect -14122 6910 -14106 6927
rect -14980 6893 -14572 6910
rect -16172 6846 -14572 6893
rect -14514 6893 -14106 6910
rect -13322 6910 -13306 6927
rect -12464 6927 -11648 6943
rect -12464 6910 -12448 6927
rect -13322 6893 -12914 6910
rect -14514 6846 -12914 6893
rect -12856 6893 -12448 6910
rect -11664 6910 -11648 6927
rect -10806 6927 -9990 6943
rect -10806 6910 -10790 6927
rect -11664 6893 -11256 6910
rect -12856 6846 -11256 6893
rect -11198 6893 -10790 6910
rect -10006 6910 -9990 6927
rect -9148 6927 -8332 6943
rect -9148 6910 -9132 6927
rect -10006 6893 -9598 6910
rect -11198 6846 -9598 6893
rect -9540 6893 -9132 6910
rect -8348 6910 -8332 6927
rect -7490 6927 -6674 6943
rect -7490 6910 -7474 6927
rect -8348 6893 -7940 6910
rect -9540 6846 -7940 6893
rect -7882 6893 -7474 6910
rect -6690 6910 -6674 6927
rect -5832 6927 -5016 6943
rect -5832 6910 -5816 6927
rect -6690 6893 -6282 6910
rect -7882 6846 -6282 6893
rect -6224 6893 -5816 6910
rect -5032 6910 -5016 6927
rect -4174 6927 -3358 6943
rect -4174 6910 -4158 6927
rect -5032 6893 -4624 6910
rect -6224 6846 -4624 6893
rect -4566 6893 -4158 6910
rect -3374 6910 -3358 6927
rect -2516 6927 -1700 6943
rect -2516 6910 -2500 6927
rect -3374 6893 -2966 6910
rect -4566 6846 -2966 6893
rect -2908 6893 -2500 6910
rect -1716 6910 -1700 6927
rect -858 6927 -42 6943
rect -858 6910 -842 6927
rect -1716 6893 -1308 6910
rect -2908 6846 -1308 6893
rect -1250 6893 -842 6910
rect -58 6910 -42 6927
rect 800 6927 1616 6943
rect 800 6910 816 6927
rect -58 6893 350 6910
rect -1250 6846 350 6893
rect 408 6893 816 6910
rect 1600 6910 1616 6927
rect 2458 6927 3274 6943
rect 2458 6910 2474 6927
rect 1600 6893 2008 6910
rect 408 6846 2008 6893
rect 2066 6893 2474 6910
rect 3258 6910 3274 6927
rect 4116 6927 4932 6943
rect 4116 6910 4132 6927
rect 3258 6893 3666 6910
rect 2066 6846 3666 6893
rect 3724 6893 4132 6910
rect 4916 6910 4932 6927
rect 5774 6927 6590 6943
rect 5774 6910 5790 6927
rect 4916 6893 5324 6910
rect 3724 6846 5324 6893
rect 5382 6893 5790 6910
rect 6574 6910 6590 6927
rect 7432 6927 8248 6943
rect 7432 6910 7448 6927
rect 6574 6893 6982 6910
rect 5382 6846 6982 6893
rect 7040 6893 7448 6910
rect 8232 6910 8248 6927
rect 9090 6927 9906 6943
rect 9090 6910 9106 6927
rect 8232 6893 8640 6910
rect 7040 6846 8640 6893
rect 8698 6893 9106 6910
rect 9890 6910 9906 6927
rect 10748 6927 11564 6943
rect 10748 6910 10764 6927
rect 9890 6893 10298 6910
rect 8698 6846 10298 6893
rect 10356 6893 10764 6910
rect 11548 6910 11564 6927
rect 12406 6927 13222 6943
rect 12406 6910 12422 6927
rect 11548 6893 11956 6910
rect 10356 6846 11956 6893
rect 12014 6893 12422 6910
rect 13206 6910 13222 6927
rect 14064 6927 14880 6943
rect 14064 6910 14080 6927
rect 13206 6893 13614 6910
rect 12014 6846 13614 6893
rect 13672 6893 14080 6910
rect 14864 6910 14880 6927
rect 15722 6927 16538 6943
rect 15722 6910 15738 6927
rect 14864 6893 15272 6910
rect 13672 6846 15272 6893
rect 15330 6893 15738 6910
rect 16522 6910 16538 6927
rect 17380 6927 18196 6943
rect 17380 6910 17396 6927
rect 16522 6893 16930 6910
rect 15330 6846 16930 6893
rect 16988 6893 17396 6910
rect 18180 6910 18196 6927
rect 19038 6927 19854 6943
rect 19038 6910 19054 6927
rect 18180 6893 18588 6910
rect 16988 6846 18588 6893
rect 18646 6893 19054 6910
rect 19838 6910 19854 6927
rect 20696 6927 21512 6943
rect 20696 6910 20712 6927
rect 19838 6893 20246 6910
rect 18646 6846 20246 6893
rect 20304 6893 20712 6910
rect 21496 6910 21512 6927
rect 22354 6927 23170 6943
rect 22354 6910 22370 6927
rect 21496 6893 21904 6910
rect 20304 6846 21904 6893
rect 21962 6893 22370 6910
rect 23154 6910 23170 6927
rect 24012 6927 24828 6943
rect 24012 6910 24028 6927
rect 23154 6893 23562 6910
rect 21962 6846 23562 6893
rect 23620 6893 24028 6910
rect 24812 6910 24828 6927
rect 25670 6927 26486 6943
rect 25670 6910 25686 6927
rect 24812 6893 25220 6910
rect 23620 6846 25220 6893
rect 25278 6893 25686 6910
rect 26470 6910 26486 6927
rect 27328 6927 28144 6943
rect 27328 6910 27344 6927
rect 26470 6893 26878 6910
rect 25278 6846 26878 6893
rect 26936 6893 27344 6910
rect 28128 6910 28144 6927
rect 28986 6927 29802 6943
rect 28986 6910 29002 6927
rect 28128 6893 28536 6910
rect 26936 6846 28536 6893
rect 28594 6893 29002 6910
rect 29786 6910 29802 6927
rect 30644 6927 31460 6943
rect 30644 6910 30660 6927
rect 29786 6893 30194 6910
rect 28594 6846 30194 6893
rect 30252 6893 30660 6910
rect 31444 6910 31460 6927
rect 32302 6927 33118 6943
rect 32302 6910 32318 6927
rect 31444 6893 31852 6910
rect 30252 6846 31852 6893
rect 31910 6893 32318 6910
rect 33102 6910 33118 6927
rect 33102 6893 33510 6910
rect 31910 6846 33510 6893
rect -32752 5399 -31152 5446
rect -32752 5382 -32344 5399
rect -32360 5365 -32344 5382
rect -31560 5382 -31152 5399
rect -31094 5399 -29494 5446
rect -31094 5382 -30686 5399
rect -31560 5365 -31544 5382
rect -32360 5349 -31544 5365
rect -30702 5365 -30686 5382
rect -29902 5382 -29494 5399
rect -29436 5399 -27836 5446
rect -29436 5382 -29028 5399
rect -29902 5365 -29886 5382
rect -30702 5349 -29886 5365
rect -29044 5365 -29028 5382
rect -28244 5382 -27836 5399
rect -27778 5399 -26178 5446
rect -27778 5382 -27370 5399
rect -28244 5365 -28228 5382
rect -29044 5349 -28228 5365
rect -27386 5365 -27370 5382
rect -26586 5382 -26178 5399
rect -26120 5399 -24520 5446
rect -26120 5382 -25712 5399
rect -26586 5365 -26570 5382
rect -27386 5349 -26570 5365
rect -25728 5365 -25712 5382
rect -24928 5382 -24520 5399
rect -24462 5399 -22862 5446
rect -24462 5382 -24054 5399
rect -24928 5365 -24912 5382
rect -25728 5349 -24912 5365
rect -24070 5365 -24054 5382
rect -23270 5382 -22862 5399
rect -22804 5399 -21204 5446
rect -22804 5382 -22396 5399
rect -23270 5365 -23254 5382
rect -24070 5349 -23254 5365
rect -22412 5365 -22396 5382
rect -21612 5382 -21204 5399
rect -21146 5399 -19546 5446
rect -21146 5382 -20738 5399
rect -21612 5365 -21596 5382
rect -22412 5349 -21596 5365
rect -20754 5365 -20738 5382
rect -19954 5382 -19546 5399
rect -19488 5399 -17888 5446
rect -19488 5382 -19080 5399
rect -19954 5365 -19938 5382
rect -20754 5349 -19938 5365
rect -19096 5365 -19080 5382
rect -18296 5382 -17888 5399
rect -17830 5399 -16230 5446
rect -17830 5382 -17422 5399
rect -18296 5365 -18280 5382
rect -19096 5349 -18280 5365
rect -17438 5365 -17422 5382
rect -16638 5382 -16230 5399
rect -16172 5399 -14572 5446
rect -16172 5382 -15764 5399
rect -16638 5365 -16622 5382
rect -17438 5349 -16622 5365
rect -15780 5365 -15764 5382
rect -14980 5382 -14572 5399
rect -14514 5399 -12914 5446
rect -14514 5382 -14106 5399
rect -14980 5365 -14964 5382
rect -15780 5349 -14964 5365
rect -14122 5365 -14106 5382
rect -13322 5382 -12914 5399
rect -12856 5399 -11256 5446
rect -12856 5382 -12448 5399
rect -13322 5365 -13306 5382
rect -14122 5349 -13306 5365
rect -12464 5365 -12448 5382
rect -11664 5382 -11256 5399
rect -11198 5399 -9598 5446
rect -11198 5382 -10790 5399
rect -11664 5365 -11648 5382
rect -12464 5349 -11648 5365
rect -10806 5365 -10790 5382
rect -10006 5382 -9598 5399
rect -9540 5399 -7940 5446
rect -9540 5382 -9132 5399
rect -10006 5365 -9990 5382
rect -10806 5349 -9990 5365
rect -9148 5365 -9132 5382
rect -8348 5382 -7940 5399
rect -7882 5399 -6282 5446
rect -7882 5382 -7474 5399
rect -8348 5365 -8332 5382
rect -9148 5349 -8332 5365
rect -7490 5365 -7474 5382
rect -6690 5382 -6282 5399
rect -6224 5399 -4624 5446
rect -6224 5382 -5816 5399
rect -6690 5365 -6674 5382
rect -7490 5349 -6674 5365
rect -5832 5365 -5816 5382
rect -5032 5382 -4624 5399
rect -4566 5399 -2966 5446
rect -4566 5382 -4158 5399
rect -5032 5365 -5016 5382
rect -5832 5349 -5016 5365
rect -4174 5365 -4158 5382
rect -3374 5382 -2966 5399
rect -2908 5399 -1308 5446
rect -2908 5382 -2500 5399
rect -3374 5365 -3358 5382
rect -4174 5349 -3358 5365
rect -2516 5365 -2500 5382
rect -1716 5382 -1308 5399
rect -1250 5399 350 5446
rect -1250 5382 -842 5399
rect -1716 5365 -1700 5382
rect -2516 5349 -1700 5365
rect -858 5365 -842 5382
rect -58 5382 350 5399
rect 408 5399 2008 5446
rect 408 5382 816 5399
rect -58 5365 -42 5382
rect -858 5349 -42 5365
rect 800 5365 816 5382
rect 1600 5382 2008 5399
rect 2066 5399 3666 5446
rect 2066 5382 2474 5399
rect 1600 5365 1616 5382
rect 800 5349 1616 5365
rect 2458 5365 2474 5382
rect 3258 5382 3666 5399
rect 3724 5399 5324 5446
rect 3724 5382 4132 5399
rect 3258 5365 3274 5382
rect 2458 5349 3274 5365
rect 4116 5365 4132 5382
rect 4916 5382 5324 5399
rect 5382 5399 6982 5446
rect 5382 5382 5790 5399
rect 4916 5365 4932 5382
rect 4116 5349 4932 5365
rect 5774 5365 5790 5382
rect 6574 5382 6982 5399
rect 7040 5399 8640 5446
rect 7040 5382 7448 5399
rect 6574 5365 6590 5382
rect 5774 5349 6590 5365
rect 7432 5365 7448 5382
rect 8232 5382 8640 5399
rect 8698 5399 10298 5446
rect 8698 5382 9106 5399
rect 8232 5365 8248 5382
rect 7432 5349 8248 5365
rect 9090 5365 9106 5382
rect 9890 5382 10298 5399
rect 10356 5399 11956 5446
rect 10356 5382 10764 5399
rect 9890 5365 9906 5382
rect 9090 5349 9906 5365
rect 10748 5365 10764 5382
rect 11548 5382 11956 5399
rect 12014 5399 13614 5446
rect 12014 5382 12422 5399
rect 11548 5365 11564 5382
rect 10748 5349 11564 5365
rect 12406 5365 12422 5382
rect 13206 5382 13614 5399
rect 13672 5399 15272 5446
rect 13672 5382 14080 5399
rect 13206 5365 13222 5382
rect 12406 5349 13222 5365
rect 14064 5365 14080 5382
rect 14864 5382 15272 5399
rect 15330 5399 16930 5446
rect 15330 5382 15738 5399
rect 14864 5365 14880 5382
rect 14064 5349 14880 5365
rect 15722 5365 15738 5382
rect 16522 5382 16930 5399
rect 16988 5399 18588 5446
rect 16988 5382 17396 5399
rect 16522 5365 16538 5382
rect 15722 5349 16538 5365
rect 17380 5365 17396 5382
rect 18180 5382 18588 5399
rect 18646 5399 20246 5446
rect 18646 5382 19054 5399
rect 18180 5365 18196 5382
rect 17380 5349 18196 5365
rect 19038 5365 19054 5382
rect 19838 5382 20246 5399
rect 20304 5399 21904 5446
rect 20304 5382 20712 5399
rect 19838 5365 19854 5382
rect 19038 5349 19854 5365
rect 20696 5365 20712 5382
rect 21496 5382 21904 5399
rect 21962 5399 23562 5446
rect 21962 5382 22370 5399
rect 21496 5365 21512 5382
rect 20696 5349 21512 5365
rect 22354 5365 22370 5382
rect 23154 5382 23562 5399
rect 23620 5399 25220 5446
rect 23620 5382 24028 5399
rect 23154 5365 23170 5382
rect 22354 5349 23170 5365
rect 24012 5365 24028 5382
rect 24812 5382 25220 5399
rect 25278 5399 26878 5446
rect 25278 5382 25686 5399
rect 24812 5365 24828 5382
rect 24012 5349 24828 5365
rect 25670 5365 25686 5382
rect 26470 5382 26878 5399
rect 26936 5399 28536 5446
rect 26936 5382 27344 5399
rect 26470 5365 26486 5382
rect 25670 5349 26486 5365
rect 27328 5365 27344 5382
rect 28128 5382 28536 5399
rect 28594 5399 30194 5446
rect 28594 5382 29002 5399
rect 28128 5365 28144 5382
rect 27328 5349 28144 5365
rect 28986 5365 29002 5382
rect 29786 5382 30194 5399
rect 30252 5399 31852 5446
rect 30252 5382 30660 5399
rect 29786 5365 29802 5382
rect 28986 5349 29802 5365
rect 30644 5365 30660 5382
rect 31444 5382 31852 5399
rect 31910 5399 33510 5446
rect 31910 5382 32318 5399
rect 31444 5365 31460 5382
rect 30644 5349 31460 5365
rect 32302 5365 32318 5382
rect 33102 5382 33510 5399
rect 33102 5365 33118 5382
rect 32302 5349 33118 5365
rect -32360 5291 -31544 5307
rect -32360 5274 -32344 5291
rect -32752 5257 -32344 5274
rect -31560 5274 -31544 5291
rect -30702 5291 -29886 5307
rect -30702 5274 -30686 5291
rect -31560 5257 -31152 5274
rect -32752 5210 -31152 5257
rect -31094 5257 -30686 5274
rect -29902 5274 -29886 5291
rect -29044 5291 -28228 5307
rect -29044 5274 -29028 5291
rect -29902 5257 -29494 5274
rect -31094 5210 -29494 5257
rect -29436 5257 -29028 5274
rect -28244 5274 -28228 5291
rect -27386 5291 -26570 5307
rect -27386 5274 -27370 5291
rect -28244 5257 -27836 5274
rect -29436 5210 -27836 5257
rect -27778 5257 -27370 5274
rect -26586 5274 -26570 5291
rect -25728 5291 -24912 5307
rect -25728 5274 -25712 5291
rect -26586 5257 -26178 5274
rect -27778 5210 -26178 5257
rect -26120 5257 -25712 5274
rect -24928 5274 -24912 5291
rect -24070 5291 -23254 5307
rect -24070 5274 -24054 5291
rect -24928 5257 -24520 5274
rect -26120 5210 -24520 5257
rect -24462 5257 -24054 5274
rect -23270 5274 -23254 5291
rect -22412 5291 -21596 5307
rect -22412 5274 -22396 5291
rect -23270 5257 -22862 5274
rect -24462 5210 -22862 5257
rect -22804 5257 -22396 5274
rect -21612 5274 -21596 5291
rect -20754 5291 -19938 5307
rect -20754 5274 -20738 5291
rect -21612 5257 -21204 5274
rect -22804 5210 -21204 5257
rect -21146 5257 -20738 5274
rect -19954 5274 -19938 5291
rect -19096 5291 -18280 5307
rect -19096 5274 -19080 5291
rect -19954 5257 -19546 5274
rect -21146 5210 -19546 5257
rect -19488 5257 -19080 5274
rect -18296 5274 -18280 5291
rect -17438 5291 -16622 5307
rect -17438 5274 -17422 5291
rect -18296 5257 -17888 5274
rect -19488 5210 -17888 5257
rect -17830 5257 -17422 5274
rect -16638 5274 -16622 5291
rect -15780 5291 -14964 5307
rect -15780 5274 -15764 5291
rect -16638 5257 -16230 5274
rect -17830 5210 -16230 5257
rect -16172 5257 -15764 5274
rect -14980 5274 -14964 5291
rect -14122 5291 -13306 5307
rect -14122 5274 -14106 5291
rect -14980 5257 -14572 5274
rect -16172 5210 -14572 5257
rect -14514 5257 -14106 5274
rect -13322 5274 -13306 5291
rect -12464 5291 -11648 5307
rect -12464 5274 -12448 5291
rect -13322 5257 -12914 5274
rect -14514 5210 -12914 5257
rect -12856 5257 -12448 5274
rect -11664 5274 -11648 5291
rect -10806 5291 -9990 5307
rect -10806 5274 -10790 5291
rect -11664 5257 -11256 5274
rect -12856 5210 -11256 5257
rect -11198 5257 -10790 5274
rect -10006 5274 -9990 5291
rect -9148 5291 -8332 5307
rect -9148 5274 -9132 5291
rect -10006 5257 -9598 5274
rect -11198 5210 -9598 5257
rect -9540 5257 -9132 5274
rect -8348 5274 -8332 5291
rect -7490 5291 -6674 5307
rect -7490 5274 -7474 5291
rect -8348 5257 -7940 5274
rect -9540 5210 -7940 5257
rect -7882 5257 -7474 5274
rect -6690 5274 -6674 5291
rect -5832 5291 -5016 5307
rect -5832 5274 -5816 5291
rect -6690 5257 -6282 5274
rect -7882 5210 -6282 5257
rect -6224 5257 -5816 5274
rect -5032 5274 -5016 5291
rect -4174 5291 -3358 5307
rect -4174 5274 -4158 5291
rect -5032 5257 -4624 5274
rect -6224 5210 -4624 5257
rect -4566 5257 -4158 5274
rect -3374 5274 -3358 5291
rect -2516 5291 -1700 5307
rect -2516 5274 -2500 5291
rect -3374 5257 -2966 5274
rect -4566 5210 -2966 5257
rect -2908 5257 -2500 5274
rect -1716 5274 -1700 5291
rect -858 5291 -42 5307
rect -858 5274 -842 5291
rect -1716 5257 -1308 5274
rect -2908 5210 -1308 5257
rect -1250 5257 -842 5274
rect -58 5274 -42 5291
rect 800 5291 1616 5307
rect 800 5274 816 5291
rect -58 5257 350 5274
rect -1250 5210 350 5257
rect 408 5257 816 5274
rect 1600 5274 1616 5291
rect 2458 5291 3274 5307
rect 2458 5274 2474 5291
rect 1600 5257 2008 5274
rect 408 5210 2008 5257
rect 2066 5257 2474 5274
rect 3258 5274 3274 5291
rect 4116 5291 4932 5307
rect 4116 5274 4132 5291
rect 3258 5257 3666 5274
rect 2066 5210 3666 5257
rect 3724 5257 4132 5274
rect 4916 5274 4932 5291
rect 5774 5291 6590 5307
rect 5774 5274 5790 5291
rect 4916 5257 5324 5274
rect 3724 5210 5324 5257
rect 5382 5257 5790 5274
rect 6574 5274 6590 5291
rect 7432 5291 8248 5307
rect 7432 5274 7448 5291
rect 6574 5257 6982 5274
rect 5382 5210 6982 5257
rect 7040 5257 7448 5274
rect 8232 5274 8248 5291
rect 9090 5291 9906 5307
rect 9090 5274 9106 5291
rect 8232 5257 8640 5274
rect 7040 5210 8640 5257
rect 8698 5257 9106 5274
rect 9890 5274 9906 5291
rect 10748 5291 11564 5307
rect 10748 5274 10764 5291
rect 9890 5257 10298 5274
rect 8698 5210 10298 5257
rect 10356 5257 10764 5274
rect 11548 5274 11564 5291
rect 12406 5291 13222 5307
rect 12406 5274 12422 5291
rect 11548 5257 11956 5274
rect 10356 5210 11956 5257
rect 12014 5257 12422 5274
rect 13206 5274 13222 5291
rect 14064 5291 14880 5307
rect 14064 5274 14080 5291
rect 13206 5257 13614 5274
rect 12014 5210 13614 5257
rect 13672 5257 14080 5274
rect 14864 5274 14880 5291
rect 15722 5291 16538 5307
rect 15722 5274 15738 5291
rect 14864 5257 15272 5274
rect 13672 5210 15272 5257
rect 15330 5257 15738 5274
rect 16522 5274 16538 5291
rect 17380 5291 18196 5307
rect 17380 5274 17396 5291
rect 16522 5257 16930 5274
rect 15330 5210 16930 5257
rect 16988 5257 17396 5274
rect 18180 5274 18196 5291
rect 19038 5291 19854 5307
rect 19038 5274 19054 5291
rect 18180 5257 18588 5274
rect 16988 5210 18588 5257
rect 18646 5257 19054 5274
rect 19838 5274 19854 5291
rect 20696 5291 21512 5307
rect 20696 5274 20712 5291
rect 19838 5257 20246 5274
rect 18646 5210 20246 5257
rect 20304 5257 20712 5274
rect 21496 5274 21512 5291
rect 22354 5291 23170 5307
rect 22354 5274 22370 5291
rect 21496 5257 21904 5274
rect 20304 5210 21904 5257
rect 21962 5257 22370 5274
rect 23154 5274 23170 5291
rect 24012 5291 24828 5307
rect 24012 5274 24028 5291
rect 23154 5257 23562 5274
rect 21962 5210 23562 5257
rect 23620 5257 24028 5274
rect 24812 5274 24828 5291
rect 25670 5291 26486 5307
rect 25670 5274 25686 5291
rect 24812 5257 25220 5274
rect 23620 5210 25220 5257
rect 25278 5257 25686 5274
rect 26470 5274 26486 5291
rect 27328 5291 28144 5307
rect 27328 5274 27344 5291
rect 26470 5257 26878 5274
rect 25278 5210 26878 5257
rect 26936 5257 27344 5274
rect 28128 5274 28144 5291
rect 28986 5291 29802 5307
rect 28986 5274 29002 5291
rect 28128 5257 28536 5274
rect 26936 5210 28536 5257
rect 28594 5257 29002 5274
rect 29786 5274 29802 5291
rect 30644 5291 31460 5307
rect 30644 5274 30660 5291
rect 29786 5257 30194 5274
rect 28594 5210 30194 5257
rect 30252 5257 30660 5274
rect 31444 5274 31460 5291
rect 32302 5291 33118 5307
rect 32302 5274 32318 5291
rect 31444 5257 31852 5274
rect 30252 5210 31852 5257
rect 31910 5257 32318 5274
rect 33102 5274 33118 5291
rect 33102 5257 33510 5274
rect 31910 5210 33510 5257
rect -32752 3763 -31152 3810
rect -32752 3746 -32344 3763
rect -32360 3729 -32344 3746
rect -31560 3746 -31152 3763
rect -31094 3763 -29494 3810
rect -31094 3746 -30686 3763
rect -31560 3729 -31544 3746
rect -32360 3713 -31544 3729
rect -30702 3729 -30686 3746
rect -29902 3746 -29494 3763
rect -29436 3763 -27836 3810
rect -29436 3746 -29028 3763
rect -29902 3729 -29886 3746
rect -30702 3713 -29886 3729
rect -29044 3729 -29028 3746
rect -28244 3746 -27836 3763
rect -27778 3763 -26178 3810
rect -27778 3746 -27370 3763
rect -28244 3729 -28228 3746
rect -29044 3713 -28228 3729
rect -27386 3729 -27370 3746
rect -26586 3746 -26178 3763
rect -26120 3763 -24520 3810
rect -26120 3746 -25712 3763
rect -26586 3729 -26570 3746
rect -27386 3713 -26570 3729
rect -25728 3729 -25712 3746
rect -24928 3746 -24520 3763
rect -24462 3763 -22862 3810
rect -24462 3746 -24054 3763
rect -24928 3729 -24912 3746
rect -25728 3713 -24912 3729
rect -24070 3729 -24054 3746
rect -23270 3746 -22862 3763
rect -22804 3763 -21204 3810
rect -22804 3746 -22396 3763
rect -23270 3729 -23254 3746
rect -24070 3713 -23254 3729
rect -22412 3729 -22396 3746
rect -21612 3746 -21204 3763
rect -21146 3763 -19546 3810
rect -21146 3746 -20738 3763
rect -21612 3729 -21596 3746
rect -22412 3713 -21596 3729
rect -20754 3729 -20738 3746
rect -19954 3746 -19546 3763
rect -19488 3763 -17888 3810
rect -19488 3746 -19080 3763
rect -19954 3729 -19938 3746
rect -20754 3713 -19938 3729
rect -19096 3729 -19080 3746
rect -18296 3746 -17888 3763
rect -17830 3763 -16230 3810
rect -17830 3746 -17422 3763
rect -18296 3729 -18280 3746
rect -19096 3713 -18280 3729
rect -17438 3729 -17422 3746
rect -16638 3746 -16230 3763
rect -16172 3763 -14572 3810
rect -16172 3746 -15764 3763
rect -16638 3729 -16622 3746
rect -17438 3713 -16622 3729
rect -15780 3729 -15764 3746
rect -14980 3746 -14572 3763
rect -14514 3763 -12914 3810
rect -14514 3746 -14106 3763
rect -14980 3729 -14964 3746
rect -15780 3713 -14964 3729
rect -14122 3729 -14106 3746
rect -13322 3746 -12914 3763
rect -12856 3763 -11256 3810
rect -12856 3746 -12448 3763
rect -13322 3729 -13306 3746
rect -14122 3713 -13306 3729
rect -12464 3729 -12448 3746
rect -11664 3746 -11256 3763
rect -11198 3763 -9598 3810
rect -11198 3746 -10790 3763
rect -11664 3729 -11648 3746
rect -12464 3713 -11648 3729
rect -10806 3729 -10790 3746
rect -10006 3746 -9598 3763
rect -9540 3763 -7940 3810
rect -9540 3746 -9132 3763
rect -10006 3729 -9990 3746
rect -10806 3713 -9990 3729
rect -9148 3729 -9132 3746
rect -8348 3746 -7940 3763
rect -7882 3763 -6282 3810
rect -7882 3746 -7474 3763
rect -8348 3729 -8332 3746
rect -9148 3713 -8332 3729
rect -7490 3729 -7474 3746
rect -6690 3746 -6282 3763
rect -6224 3763 -4624 3810
rect -6224 3746 -5816 3763
rect -6690 3729 -6674 3746
rect -7490 3713 -6674 3729
rect -5832 3729 -5816 3746
rect -5032 3746 -4624 3763
rect -4566 3763 -2966 3810
rect -4566 3746 -4158 3763
rect -5032 3729 -5016 3746
rect -5832 3713 -5016 3729
rect -4174 3729 -4158 3746
rect -3374 3746 -2966 3763
rect -2908 3763 -1308 3810
rect -2908 3746 -2500 3763
rect -3374 3729 -3358 3746
rect -4174 3713 -3358 3729
rect -2516 3729 -2500 3746
rect -1716 3746 -1308 3763
rect -1250 3763 350 3810
rect -1250 3746 -842 3763
rect -1716 3729 -1700 3746
rect -2516 3713 -1700 3729
rect -858 3729 -842 3746
rect -58 3746 350 3763
rect 408 3763 2008 3810
rect 408 3746 816 3763
rect -58 3729 -42 3746
rect -858 3713 -42 3729
rect 800 3729 816 3746
rect 1600 3746 2008 3763
rect 2066 3763 3666 3810
rect 2066 3746 2474 3763
rect 1600 3729 1616 3746
rect 800 3713 1616 3729
rect 2458 3729 2474 3746
rect 3258 3746 3666 3763
rect 3724 3763 5324 3810
rect 3724 3746 4132 3763
rect 3258 3729 3274 3746
rect 2458 3713 3274 3729
rect 4116 3729 4132 3746
rect 4916 3746 5324 3763
rect 5382 3763 6982 3810
rect 5382 3746 5790 3763
rect 4916 3729 4932 3746
rect 4116 3713 4932 3729
rect 5774 3729 5790 3746
rect 6574 3746 6982 3763
rect 7040 3763 8640 3810
rect 7040 3746 7448 3763
rect 6574 3729 6590 3746
rect 5774 3713 6590 3729
rect 7432 3729 7448 3746
rect 8232 3746 8640 3763
rect 8698 3763 10298 3810
rect 8698 3746 9106 3763
rect 8232 3729 8248 3746
rect 7432 3713 8248 3729
rect 9090 3729 9106 3746
rect 9890 3746 10298 3763
rect 10356 3763 11956 3810
rect 10356 3746 10764 3763
rect 9890 3729 9906 3746
rect 9090 3713 9906 3729
rect 10748 3729 10764 3746
rect 11548 3746 11956 3763
rect 12014 3763 13614 3810
rect 12014 3746 12422 3763
rect 11548 3729 11564 3746
rect 10748 3713 11564 3729
rect 12406 3729 12422 3746
rect 13206 3746 13614 3763
rect 13672 3763 15272 3810
rect 13672 3746 14080 3763
rect 13206 3729 13222 3746
rect 12406 3713 13222 3729
rect 14064 3729 14080 3746
rect 14864 3746 15272 3763
rect 15330 3763 16930 3810
rect 15330 3746 15738 3763
rect 14864 3729 14880 3746
rect 14064 3713 14880 3729
rect 15722 3729 15738 3746
rect 16522 3746 16930 3763
rect 16988 3763 18588 3810
rect 16988 3746 17396 3763
rect 16522 3729 16538 3746
rect 15722 3713 16538 3729
rect 17380 3729 17396 3746
rect 18180 3746 18588 3763
rect 18646 3763 20246 3810
rect 18646 3746 19054 3763
rect 18180 3729 18196 3746
rect 17380 3713 18196 3729
rect 19038 3729 19054 3746
rect 19838 3746 20246 3763
rect 20304 3763 21904 3810
rect 20304 3746 20712 3763
rect 19838 3729 19854 3746
rect 19038 3713 19854 3729
rect 20696 3729 20712 3746
rect 21496 3746 21904 3763
rect 21962 3763 23562 3810
rect 21962 3746 22370 3763
rect 21496 3729 21512 3746
rect 20696 3713 21512 3729
rect 22354 3729 22370 3746
rect 23154 3746 23562 3763
rect 23620 3763 25220 3810
rect 23620 3746 24028 3763
rect 23154 3729 23170 3746
rect 22354 3713 23170 3729
rect 24012 3729 24028 3746
rect 24812 3746 25220 3763
rect 25278 3763 26878 3810
rect 25278 3746 25686 3763
rect 24812 3729 24828 3746
rect 24012 3713 24828 3729
rect 25670 3729 25686 3746
rect 26470 3746 26878 3763
rect 26936 3763 28536 3810
rect 26936 3746 27344 3763
rect 26470 3729 26486 3746
rect 25670 3713 26486 3729
rect 27328 3729 27344 3746
rect 28128 3746 28536 3763
rect 28594 3763 30194 3810
rect 28594 3746 29002 3763
rect 28128 3729 28144 3746
rect 27328 3713 28144 3729
rect 28986 3729 29002 3746
rect 29786 3746 30194 3763
rect 30252 3763 31852 3810
rect 30252 3746 30660 3763
rect 29786 3729 29802 3746
rect 28986 3713 29802 3729
rect 30644 3729 30660 3746
rect 31444 3746 31852 3763
rect 31910 3763 33510 3810
rect 31910 3746 32318 3763
rect 31444 3729 31460 3746
rect 30644 3713 31460 3729
rect 32302 3729 32318 3746
rect 33102 3746 33510 3763
rect 33102 3729 33118 3746
rect 32302 3713 33118 3729
rect -32360 3655 -31544 3671
rect -32360 3638 -32344 3655
rect -32752 3621 -32344 3638
rect -31560 3638 -31544 3655
rect -30702 3655 -29886 3671
rect -30702 3638 -30686 3655
rect -31560 3621 -31152 3638
rect -32752 3574 -31152 3621
rect -31094 3621 -30686 3638
rect -29902 3638 -29886 3655
rect -29044 3655 -28228 3671
rect -29044 3638 -29028 3655
rect -29902 3621 -29494 3638
rect -31094 3574 -29494 3621
rect -29436 3621 -29028 3638
rect -28244 3638 -28228 3655
rect -27386 3655 -26570 3671
rect -27386 3638 -27370 3655
rect -28244 3621 -27836 3638
rect -29436 3574 -27836 3621
rect -27778 3621 -27370 3638
rect -26586 3638 -26570 3655
rect -25728 3655 -24912 3671
rect -25728 3638 -25712 3655
rect -26586 3621 -26178 3638
rect -27778 3574 -26178 3621
rect -26120 3621 -25712 3638
rect -24928 3638 -24912 3655
rect -24070 3655 -23254 3671
rect -24070 3638 -24054 3655
rect -24928 3621 -24520 3638
rect -26120 3574 -24520 3621
rect -24462 3621 -24054 3638
rect -23270 3638 -23254 3655
rect -22412 3655 -21596 3671
rect -22412 3638 -22396 3655
rect -23270 3621 -22862 3638
rect -24462 3574 -22862 3621
rect -22804 3621 -22396 3638
rect -21612 3638 -21596 3655
rect -20754 3655 -19938 3671
rect -20754 3638 -20738 3655
rect -21612 3621 -21204 3638
rect -22804 3574 -21204 3621
rect -21146 3621 -20738 3638
rect -19954 3638 -19938 3655
rect -19096 3655 -18280 3671
rect -19096 3638 -19080 3655
rect -19954 3621 -19546 3638
rect -21146 3574 -19546 3621
rect -19488 3621 -19080 3638
rect -18296 3638 -18280 3655
rect -17438 3655 -16622 3671
rect -17438 3638 -17422 3655
rect -18296 3621 -17888 3638
rect -19488 3574 -17888 3621
rect -17830 3621 -17422 3638
rect -16638 3638 -16622 3655
rect -15780 3655 -14964 3671
rect -15780 3638 -15764 3655
rect -16638 3621 -16230 3638
rect -17830 3574 -16230 3621
rect -16172 3621 -15764 3638
rect -14980 3638 -14964 3655
rect -14122 3655 -13306 3671
rect -14122 3638 -14106 3655
rect -14980 3621 -14572 3638
rect -16172 3574 -14572 3621
rect -14514 3621 -14106 3638
rect -13322 3638 -13306 3655
rect -12464 3655 -11648 3671
rect -12464 3638 -12448 3655
rect -13322 3621 -12914 3638
rect -14514 3574 -12914 3621
rect -12856 3621 -12448 3638
rect -11664 3638 -11648 3655
rect -10806 3655 -9990 3671
rect -10806 3638 -10790 3655
rect -11664 3621 -11256 3638
rect -12856 3574 -11256 3621
rect -11198 3621 -10790 3638
rect -10006 3638 -9990 3655
rect -9148 3655 -8332 3671
rect -9148 3638 -9132 3655
rect -10006 3621 -9598 3638
rect -11198 3574 -9598 3621
rect -9540 3621 -9132 3638
rect -8348 3638 -8332 3655
rect -7490 3655 -6674 3671
rect -7490 3638 -7474 3655
rect -8348 3621 -7940 3638
rect -9540 3574 -7940 3621
rect -7882 3621 -7474 3638
rect -6690 3638 -6674 3655
rect -5832 3655 -5016 3671
rect -5832 3638 -5816 3655
rect -6690 3621 -6282 3638
rect -7882 3574 -6282 3621
rect -6224 3621 -5816 3638
rect -5032 3638 -5016 3655
rect -4174 3655 -3358 3671
rect -4174 3638 -4158 3655
rect -5032 3621 -4624 3638
rect -6224 3574 -4624 3621
rect -4566 3621 -4158 3638
rect -3374 3638 -3358 3655
rect -2516 3655 -1700 3671
rect -2516 3638 -2500 3655
rect -3374 3621 -2966 3638
rect -4566 3574 -2966 3621
rect -2908 3621 -2500 3638
rect -1716 3638 -1700 3655
rect -858 3655 -42 3671
rect -858 3638 -842 3655
rect -1716 3621 -1308 3638
rect -2908 3574 -1308 3621
rect -1250 3621 -842 3638
rect -58 3638 -42 3655
rect 800 3655 1616 3671
rect 800 3638 816 3655
rect -58 3621 350 3638
rect -1250 3574 350 3621
rect 408 3621 816 3638
rect 1600 3638 1616 3655
rect 2458 3655 3274 3671
rect 2458 3638 2474 3655
rect 1600 3621 2008 3638
rect 408 3574 2008 3621
rect 2066 3621 2474 3638
rect 3258 3638 3274 3655
rect 4116 3655 4932 3671
rect 4116 3638 4132 3655
rect 3258 3621 3666 3638
rect 2066 3574 3666 3621
rect 3724 3621 4132 3638
rect 4916 3638 4932 3655
rect 5774 3655 6590 3671
rect 5774 3638 5790 3655
rect 4916 3621 5324 3638
rect 3724 3574 5324 3621
rect 5382 3621 5790 3638
rect 6574 3638 6590 3655
rect 7432 3655 8248 3671
rect 7432 3638 7448 3655
rect 6574 3621 6982 3638
rect 5382 3574 6982 3621
rect 7040 3621 7448 3638
rect 8232 3638 8248 3655
rect 9090 3655 9906 3671
rect 9090 3638 9106 3655
rect 8232 3621 8640 3638
rect 7040 3574 8640 3621
rect 8698 3621 9106 3638
rect 9890 3638 9906 3655
rect 10748 3655 11564 3671
rect 10748 3638 10764 3655
rect 9890 3621 10298 3638
rect 8698 3574 10298 3621
rect 10356 3621 10764 3638
rect 11548 3638 11564 3655
rect 12406 3655 13222 3671
rect 12406 3638 12422 3655
rect 11548 3621 11956 3638
rect 10356 3574 11956 3621
rect 12014 3621 12422 3638
rect 13206 3638 13222 3655
rect 14064 3655 14880 3671
rect 14064 3638 14080 3655
rect 13206 3621 13614 3638
rect 12014 3574 13614 3621
rect 13672 3621 14080 3638
rect 14864 3638 14880 3655
rect 15722 3655 16538 3671
rect 15722 3638 15738 3655
rect 14864 3621 15272 3638
rect 13672 3574 15272 3621
rect 15330 3621 15738 3638
rect 16522 3638 16538 3655
rect 17380 3655 18196 3671
rect 17380 3638 17396 3655
rect 16522 3621 16930 3638
rect 15330 3574 16930 3621
rect 16988 3621 17396 3638
rect 18180 3638 18196 3655
rect 19038 3655 19854 3671
rect 19038 3638 19054 3655
rect 18180 3621 18588 3638
rect 16988 3574 18588 3621
rect 18646 3621 19054 3638
rect 19838 3638 19854 3655
rect 20696 3655 21512 3671
rect 20696 3638 20712 3655
rect 19838 3621 20246 3638
rect 18646 3574 20246 3621
rect 20304 3621 20712 3638
rect 21496 3638 21512 3655
rect 22354 3655 23170 3671
rect 22354 3638 22370 3655
rect 21496 3621 21904 3638
rect 20304 3574 21904 3621
rect 21962 3621 22370 3638
rect 23154 3638 23170 3655
rect 24012 3655 24828 3671
rect 24012 3638 24028 3655
rect 23154 3621 23562 3638
rect 21962 3574 23562 3621
rect 23620 3621 24028 3638
rect 24812 3638 24828 3655
rect 25670 3655 26486 3671
rect 25670 3638 25686 3655
rect 24812 3621 25220 3638
rect 23620 3574 25220 3621
rect 25278 3621 25686 3638
rect 26470 3638 26486 3655
rect 27328 3655 28144 3671
rect 27328 3638 27344 3655
rect 26470 3621 26878 3638
rect 25278 3574 26878 3621
rect 26936 3621 27344 3638
rect 28128 3638 28144 3655
rect 28986 3655 29802 3671
rect 28986 3638 29002 3655
rect 28128 3621 28536 3638
rect 26936 3574 28536 3621
rect 28594 3621 29002 3638
rect 29786 3638 29802 3655
rect 30644 3655 31460 3671
rect 30644 3638 30660 3655
rect 29786 3621 30194 3638
rect 28594 3574 30194 3621
rect 30252 3621 30660 3638
rect 31444 3638 31460 3655
rect 32302 3655 33118 3671
rect 32302 3638 32318 3655
rect 31444 3621 31852 3638
rect 30252 3574 31852 3621
rect 31910 3621 32318 3638
rect 33102 3638 33118 3655
rect 33102 3621 33510 3638
rect 31910 3574 33510 3621
rect -32752 2127 -31152 2174
rect -32752 2110 -32344 2127
rect -32360 2093 -32344 2110
rect -31560 2110 -31152 2127
rect -31094 2127 -29494 2174
rect -31094 2110 -30686 2127
rect -31560 2093 -31544 2110
rect -32360 2077 -31544 2093
rect -30702 2093 -30686 2110
rect -29902 2110 -29494 2127
rect -29436 2127 -27836 2174
rect -29436 2110 -29028 2127
rect -29902 2093 -29886 2110
rect -30702 2077 -29886 2093
rect -29044 2093 -29028 2110
rect -28244 2110 -27836 2127
rect -27778 2127 -26178 2174
rect -27778 2110 -27370 2127
rect -28244 2093 -28228 2110
rect -29044 2077 -28228 2093
rect -27386 2093 -27370 2110
rect -26586 2110 -26178 2127
rect -26120 2127 -24520 2174
rect -26120 2110 -25712 2127
rect -26586 2093 -26570 2110
rect -27386 2077 -26570 2093
rect -25728 2093 -25712 2110
rect -24928 2110 -24520 2127
rect -24462 2127 -22862 2174
rect -24462 2110 -24054 2127
rect -24928 2093 -24912 2110
rect -25728 2077 -24912 2093
rect -24070 2093 -24054 2110
rect -23270 2110 -22862 2127
rect -22804 2127 -21204 2174
rect -22804 2110 -22396 2127
rect -23270 2093 -23254 2110
rect -24070 2077 -23254 2093
rect -22412 2093 -22396 2110
rect -21612 2110 -21204 2127
rect -21146 2127 -19546 2174
rect -21146 2110 -20738 2127
rect -21612 2093 -21596 2110
rect -22412 2077 -21596 2093
rect -20754 2093 -20738 2110
rect -19954 2110 -19546 2127
rect -19488 2127 -17888 2174
rect -19488 2110 -19080 2127
rect -19954 2093 -19938 2110
rect -20754 2077 -19938 2093
rect -19096 2093 -19080 2110
rect -18296 2110 -17888 2127
rect -17830 2127 -16230 2174
rect -17830 2110 -17422 2127
rect -18296 2093 -18280 2110
rect -19096 2077 -18280 2093
rect -17438 2093 -17422 2110
rect -16638 2110 -16230 2127
rect -16172 2127 -14572 2174
rect -16172 2110 -15764 2127
rect -16638 2093 -16622 2110
rect -17438 2077 -16622 2093
rect -15780 2093 -15764 2110
rect -14980 2110 -14572 2127
rect -14514 2127 -12914 2174
rect -14514 2110 -14106 2127
rect -14980 2093 -14964 2110
rect -15780 2077 -14964 2093
rect -14122 2093 -14106 2110
rect -13322 2110 -12914 2127
rect -12856 2127 -11256 2174
rect -12856 2110 -12448 2127
rect -13322 2093 -13306 2110
rect -14122 2077 -13306 2093
rect -12464 2093 -12448 2110
rect -11664 2110 -11256 2127
rect -11198 2127 -9598 2174
rect -11198 2110 -10790 2127
rect -11664 2093 -11648 2110
rect -12464 2077 -11648 2093
rect -10806 2093 -10790 2110
rect -10006 2110 -9598 2127
rect -9540 2127 -7940 2174
rect -9540 2110 -9132 2127
rect -10006 2093 -9990 2110
rect -10806 2077 -9990 2093
rect -9148 2093 -9132 2110
rect -8348 2110 -7940 2127
rect -7882 2127 -6282 2174
rect -7882 2110 -7474 2127
rect -8348 2093 -8332 2110
rect -9148 2077 -8332 2093
rect -7490 2093 -7474 2110
rect -6690 2110 -6282 2127
rect -6224 2127 -4624 2174
rect -6224 2110 -5816 2127
rect -6690 2093 -6674 2110
rect -7490 2077 -6674 2093
rect -5832 2093 -5816 2110
rect -5032 2110 -4624 2127
rect -4566 2127 -2966 2174
rect -4566 2110 -4158 2127
rect -5032 2093 -5016 2110
rect -5832 2077 -5016 2093
rect -4174 2093 -4158 2110
rect -3374 2110 -2966 2127
rect -2908 2127 -1308 2174
rect -2908 2110 -2500 2127
rect -3374 2093 -3358 2110
rect -4174 2077 -3358 2093
rect -2516 2093 -2500 2110
rect -1716 2110 -1308 2127
rect -1250 2127 350 2174
rect -1250 2110 -842 2127
rect -1716 2093 -1700 2110
rect -2516 2077 -1700 2093
rect -858 2093 -842 2110
rect -58 2110 350 2127
rect 408 2127 2008 2174
rect 408 2110 816 2127
rect -58 2093 -42 2110
rect -858 2077 -42 2093
rect 800 2093 816 2110
rect 1600 2110 2008 2127
rect 2066 2127 3666 2174
rect 2066 2110 2474 2127
rect 1600 2093 1616 2110
rect 800 2077 1616 2093
rect 2458 2093 2474 2110
rect 3258 2110 3666 2127
rect 3724 2127 5324 2174
rect 3724 2110 4132 2127
rect 3258 2093 3274 2110
rect 2458 2077 3274 2093
rect 4116 2093 4132 2110
rect 4916 2110 5324 2127
rect 5382 2127 6982 2174
rect 5382 2110 5790 2127
rect 4916 2093 4932 2110
rect 4116 2077 4932 2093
rect 5774 2093 5790 2110
rect 6574 2110 6982 2127
rect 7040 2127 8640 2174
rect 7040 2110 7448 2127
rect 6574 2093 6590 2110
rect 5774 2077 6590 2093
rect 7432 2093 7448 2110
rect 8232 2110 8640 2127
rect 8698 2127 10298 2174
rect 8698 2110 9106 2127
rect 8232 2093 8248 2110
rect 7432 2077 8248 2093
rect 9090 2093 9106 2110
rect 9890 2110 10298 2127
rect 10356 2127 11956 2174
rect 10356 2110 10764 2127
rect 9890 2093 9906 2110
rect 9090 2077 9906 2093
rect 10748 2093 10764 2110
rect 11548 2110 11956 2127
rect 12014 2127 13614 2174
rect 12014 2110 12422 2127
rect 11548 2093 11564 2110
rect 10748 2077 11564 2093
rect 12406 2093 12422 2110
rect 13206 2110 13614 2127
rect 13672 2127 15272 2174
rect 13672 2110 14080 2127
rect 13206 2093 13222 2110
rect 12406 2077 13222 2093
rect 14064 2093 14080 2110
rect 14864 2110 15272 2127
rect 15330 2127 16930 2174
rect 15330 2110 15738 2127
rect 14864 2093 14880 2110
rect 14064 2077 14880 2093
rect 15722 2093 15738 2110
rect 16522 2110 16930 2127
rect 16988 2127 18588 2174
rect 16988 2110 17396 2127
rect 16522 2093 16538 2110
rect 15722 2077 16538 2093
rect 17380 2093 17396 2110
rect 18180 2110 18588 2127
rect 18646 2127 20246 2174
rect 18646 2110 19054 2127
rect 18180 2093 18196 2110
rect 17380 2077 18196 2093
rect 19038 2093 19054 2110
rect 19838 2110 20246 2127
rect 20304 2127 21904 2174
rect 20304 2110 20712 2127
rect 19838 2093 19854 2110
rect 19038 2077 19854 2093
rect 20696 2093 20712 2110
rect 21496 2110 21904 2127
rect 21962 2127 23562 2174
rect 21962 2110 22370 2127
rect 21496 2093 21512 2110
rect 20696 2077 21512 2093
rect 22354 2093 22370 2110
rect 23154 2110 23562 2127
rect 23620 2127 25220 2174
rect 23620 2110 24028 2127
rect 23154 2093 23170 2110
rect 22354 2077 23170 2093
rect 24012 2093 24028 2110
rect 24812 2110 25220 2127
rect 25278 2127 26878 2174
rect 25278 2110 25686 2127
rect 24812 2093 24828 2110
rect 24012 2077 24828 2093
rect 25670 2093 25686 2110
rect 26470 2110 26878 2127
rect 26936 2127 28536 2174
rect 26936 2110 27344 2127
rect 26470 2093 26486 2110
rect 25670 2077 26486 2093
rect 27328 2093 27344 2110
rect 28128 2110 28536 2127
rect 28594 2127 30194 2174
rect 28594 2110 29002 2127
rect 28128 2093 28144 2110
rect 27328 2077 28144 2093
rect 28986 2093 29002 2110
rect 29786 2110 30194 2127
rect 30252 2127 31852 2174
rect 30252 2110 30660 2127
rect 29786 2093 29802 2110
rect 28986 2077 29802 2093
rect 30644 2093 30660 2110
rect 31444 2110 31852 2127
rect 31910 2127 33510 2174
rect 31910 2110 32318 2127
rect 31444 2093 31460 2110
rect 30644 2077 31460 2093
rect 32302 2093 32318 2110
rect 33102 2110 33510 2127
rect 33102 2093 33118 2110
rect 32302 2077 33118 2093
rect -32360 2019 -31544 2035
rect -32360 2002 -32344 2019
rect -32752 1985 -32344 2002
rect -31560 2002 -31544 2019
rect -30702 2019 -29886 2035
rect -30702 2002 -30686 2019
rect -31560 1985 -31152 2002
rect -32752 1938 -31152 1985
rect -31094 1985 -30686 2002
rect -29902 2002 -29886 2019
rect -29044 2019 -28228 2035
rect -29044 2002 -29028 2019
rect -29902 1985 -29494 2002
rect -31094 1938 -29494 1985
rect -29436 1985 -29028 2002
rect -28244 2002 -28228 2019
rect -27386 2019 -26570 2035
rect -27386 2002 -27370 2019
rect -28244 1985 -27836 2002
rect -29436 1938 -27836 1985
rect -27778 1985 -27370 2002
rect -26586 2002 -26570 2019
rect -25728 2019 -24912 2035
rect -25728 2002 -25712 2019
rect -26586 1985 -26178 2002
rect -27778 1938 -26178 1985
rect -26120 1985 -25712 2002
rect -24928 2002 -24912 2019
rect -24070 2019 -23254 2035
rect -24070 2002 -24054 2019
rect -24928 1985 -24520 2002
rect -26120 1938 -24520 1985
rect -24462 1985 -24054 2002
rect -23270 2002 -23254 2019
rect -22412 2019 -21596 2035
rect -22412 2002 -22396 2019
rect -23270 1985 -22862 2002
rect -24462 1938 -22862 1985
rect -22804 1985 -22396 2002
rect -21612 2002 -21596 2019
rect -20754 2019 -19938 2035
rect -20754 2002 -20738 2019
rect -21612 1985 -21204 2002
rect -22804 1938 -21204 1985
rect -21146 1985 -20738 2002
rect -19954 2002 -19938 2019
rect -19096 2019 -18280 2035
rect -19096 2002 -19080 2019
rect -19954 1985 -19546 2002
rect -21146 1938 -19546 1985
rect -19488 1985 -19080 2002
rect -18296 2002 -18280 2019
rect -17438 2019 -16622 2035
rect -17438 2002 -17422 2019
rect -18296 1985 -17888 2002
rect -19488 1938 -17888 1985
rect -17830 1985 -17422 2002
rect -16638 2002 -16622 2019
rect -15780 2019 -14964 2035
rect -15780 2002 -15764 2019
rect -16638 1985 -16230 2002
rect -17830 1938 -16230 1985
rect -16172 1985 -15764 2002
rect -14980 2002 -14964 2019
rect -14122 2019 -13306 2035
rect -14122 2002 -14106 2019
rect -14980 1985 -14572 2002
rect -16172 1938 -14572 1985
rect -14514 1985 -14106 2002
rect -13322 2002 -13306 2019
rect -12464 2019 -11648 2035
rect -12464 2002 -12448 2019
rect -13322 1985 -12914 2002
rect -14514 1938 -12914 1985
rect -12856 1985 -12448 2002
rect -11664 2002 -11648 2019
rect -10806 2019 -9990 2035
rect -10806 2002 -10790 2019
rect -11664 1985 -11256 2002
rect -12856 1938 -11256 1985
rect -11198 1985 -10790 2002
rect -10006 2002 -9990 2019
rect -9148 2019 -8332 2035
rect -9148 2002 -9132 2019
rect -10006 1985 -9598 2002
rect -11198 1938 -9598 1985
rect -9540 1985 -9132 2002
rect -8348 2002 -8332 2019
rect -7490 2019 -6674 2035
rect -7490 2002 -7474 2019
rect -8348 1985 -7940 2002
rect -9540 1938 -7940 1985
rect -7882 1985 -7474 2002
rect -6690 2002 -6674 2019
rect -5832 2019 -5016 2035
rect -5832 2002 -5816 2019
rect -6690 1985 -6282 2002
rect -7882 1938 -6282 1985
rect -6224 1985 -5816 2002
rect -5032 2002 -5016 2019
rect -4174 2019 -3358 2035
rect -4174 2002 -4158 2019
rect -5032 1985 -4624 2002
rect -6224 1938 -4624 1985
rect -4566 1985 -4158 2002
rect -3374 2002 -3358 2019
rect -2516 2019 -1700 2035
rect -2516 2002 -2500 2019
rect -3374 1985 -2966 2002
rect -4566 1938 -2966 1985
rect -2908 1985 -2500 2002
rect -1716 2002 -1700 2019
rect -858 2019 -42 2035
rect -858 2002 -842 2019
rect -1716 1985 -1308 2002
rect -2908 1938 -1308 1985
rect -1250 1985 -842 2002
rect -58 2002 -42 2019
rect 800 2019 1616 2035
rect 800 2002 816 2019
rect -58 1985 350 2002
rect -1250 1938 350 1985
rect 408 1985 816 2002
rect 1600 2002 1616 2019
rect 2458 2019 3274 2035
rect 2458 2002 2474 2019
rect 1600 1985 2008 2002
rect 408 1938 2008 1985
rect 2066 1985 2474 2002
rect 3258 2002 3274 2019
rect 4116 2019 4932 2035
rect 4116 2002 4132 2019
rect 3258 1985 3666 2002
rect 2066 1938 3666 1985
rect 3724 1985 4132 2002
rect 4916 2002 4932 2019
rect 5774 2019 6590 2035
rect 5774 2002 5790 2019
rect 4916 1985 5324 2002
rect 3724 1938 5324 1985
rect 5382 1985 5790 2002
rect 6574 2002 6590 2019
rect 7432 2019 8248 2035
rect 7432 2002 7448 2019
rect 6574 1985 6982 2002
rect 5382 1938 6982 1985
rect 7040 1985 7448 2002
rect 8232 2002 8248 2019
rect 9090 2019 9906 2035
rect 9090 2002 9106 2019
rect 8232 1985 8640 2002
rect 7040 1938 8640 1985
rect 8698 1985 9106 2002
rect 9890 2002 9906 2019
rect 10748 2019 11564 2035
rect 10748 2002 10764 2019
rect 9890 1985 10298 2002
rect 8698 1938 10298 1985
rect 10356 1985 10764 2002
rect 11548 2002 11564 2019
rect 12406 2019 13222 2035
rect 12406 2002 12422 2019
rect 11548 1985 11956 2002
rect 10356 1938 11956 1985
rect 12014 1985 12422 2002
rect 13206 2002 13222 2019
rect 14064 2019 14880 2035
rect 14064 2002 14080 2019
rect 13206 1985 13614 2002
rect 12014 1938 13614 1985
rect 13672 1985 14080 2002
rect 14864 2002 14880 2019
rect 15722 2019 16538 2035
rect 15722 2002 15738 2019
rect 14864 1985 15272 2002
rect 13672 1938 15272 1985
rect 15330 1985 15738 2002
rect 16522 2002 16538 2019
rect 17380 2019 18196 2035
rect 17380 2002 17396 2019
rect 16522 1985 16930 2002
rect 15330 1938 16930 1985
rect 16988 1985 17396 2002
rect 18180 2002 18196 2019
rect 19038 2019 19854 2035
rect 19038 2002 19054 2019
rect 18180 1985 18588 2002
rect 16988 1938 18588 1985
rect 18646 1985 19054 2002
rect 19838 2002 19854 2019
rect 20696 2019 21512 2035
rect 20696 2002 20712 2019
rect 19838 1985 20246 2002
rect 18646 1938 20246 1985
rect 20304 1985 20712 2002
rect 21496 2002 21512 2019
rect 22354 2019 23170 2035
rect 22354 2002 22370 2019
rect 21496 1985 21904 2002
rect 20304 1938 21904 1985
rect 21962 1985 22370 2002
rect 23154 2002 23170 2019
rect 24012 2019 24828 2035
rect 24012 2002 24028 2019
rect 23154 1985 23562 2002
rect 21962 1938 23562 1985
rect 23620 1985 24028 2002
rect 24812 2002 24828 2019
rect 25670 2019 26486 2035
rect 25670 2002 25686 2019
rect 24812 1985 25220 2002
rect 23620 1938 25220 1985
rect 25278 1985 25686 2002
rect 26470 2002 26486 2019
rect 27328 2019 28144 2035
rect 27328 2002 27344 2019
rect 26470 1985 26878 2002
rect 25278 1938 26878 1985
rect 26936 1985 27344 2002
rect 28128 2002 28144 2019
rect 28986 2019 29802 2035
rect 28986 2002 29002 2019
rect 28128 1985 28536 2002
rect 26936 1938 28536 1985
rect 28594 1985 29002 2002
rect 29786 2002 29802 2019
rect 30644 2019 31460 2035
rect 30644 2002 30660 2019
rect 29786 1985 30194 2002
rect 28594 1938 30194 1985
rect 30252 1985 30660 2002
rect 31444 2002 31460 2019
rect 32302 2019 33118 2035
rect 32302 2002 32318 2019
rect 31444 1985 31852 2002
rect 30252 1938 31852 1985
rect 31910 1985 32318 2002
rect 33102 2002 33118 2019
rect 33102 1985 33510 2002
rect 31910 1938 33510 1985
rect -32752 491 -31152 538
rect -32752 474 -32344 491
rect -32360 457 -32344 474
rect -31560 474 -31152 491
rect -31094 491 -29494 538
rect -31094 474 -30686 491
rect -31560 457 -31544 474
rect -32360 441 -31544 457
rect -30702 457 -30686 474
rect -29902 474 -29494 491
rect -29436 491 -27836 538
rect -29436 474 -29028 491
rect -29902 457 -29886 474
rect -30702 441 -29886 457
rect -29044 457 -29028 474
rect -28244 474 -27836 491
rect -27778 491 -26178 538
rect -27778 474 -27370 491
rect -28244 457 -28228 474
rect -29044 441 -28228 457
rect -27386 457 -27370 474
rect -26586 474 -26178 491
rect -26120 491 -24520 538
rect -26120 474 -25712 491
rect -26586 457 -26570 474
rect -27386 441 -26570 457
rect -25728 457 -25712 474
rect -24928 474 -24520 491
rect -24462 491 -22862 538
rect -24462 474 -24054 491
rect -24928 457 -24912 474
rect -25728 441 -24912 457
rect -24070 457 -24054 474
rect -23270 474 -22862 491
rect -22804 491 -21204 538
rect -22804 474 -22396 491
rect -23270 457 -23254 474
rect -24070 441 -23254 457
rect -22412 457 -22396 474
rect -21612 474 -21204 491
rect -21146 491 -19546 538
rect -21146 474 -20738 491
rect -21612 457 -21596 474
rect -22412 441 -21596 457
rect -20754 457 -20738 474
rect -19954 474 -19546 491
rect -19488 491 -17888 538
rect -19488 474 -19080 491
rect -19954 457 -19938 474
rect -20754 441 -19938 457
rect -19096 457 -19080 474
rect -18296 474 -17888 491
rect -17830 491 -16230 538
rect -17830 474 -17422 491
rect -18296 457 -18280 474
rect -19096 441 -18280 457
rect -17438 457 -17422 474
rect -16638 474 -16230 491
rect -16172 491 -14572 538
rect -16172 474 -15764 491
rect -16638 457 -16622 474
rect -17438 441 -16622 457
rect -15780 457 -15764 474
rect -14980 474 -14572 491
rect -14514 491 -12914 538
rect -14514 474 -14106 491
rect -14980 457 -14964 474
rect -15780 441 -14964 457
rect -14122 457 -14106 474
rect -13322 474 -12914 491
rect -12856 491 -11256 538
rect -12856 474 -12448 491
rect -13322 457 -13306 474
rect -14122 441 -13306 457
rect -12464 457 -12448 474
rect -11664 474 -11256 491
rect -11198 491 -9598 538
rect -11198 474 -10790 491
rect -11664 457 -11648 474
rect -12464 441 -11648 457
rect -10806 457 -10790 474
rect -10006 474 -9598 491
rect -9540 491 -7940 538
rect -9540 474 -9132 491
rect -10006 457 -9990 474
rect -10806 441 -9990 457
rect -9148 457 -9132 474
rect -8348 474 -7940 491
rect -7882 491 -6282 538
rect -7882 474 -7474 491
rect -8348 457 -8332 474
rect -9148 441 -8332 457
rect -7490 457 -7474 474
rect -6690 474 -6282 491
rect -6224 491 -4624 538
rect -6224 474 -5816 491
rect -6690 457 -6674 474
rect -7490 441 -6674 457
rect -5832 457 -5816 474
rect -5032 474 -4624 491
rect -4566 491 -2966 538
rect -4566 474 -4158 491
rect -5032 457 -5016 474
rect -5832 441 -5016 457
rect -4174 457 -4158 474
rect -3374 474 -2966 491
rect -2908 491 -1308 538
rect -2908 474 -2500 491
rect -3374 457 -3358 474
rect -4174 441 -3358 457
rect -2516 457 -2500 474
rect -1716 474 -1308 491
rect -1250 491 350 538
rect -1250 474 -842 491
rect -1716 457 -1700 474
rect -2516 441 -1700 457
rect -858 457 -842 474
rect -58 474 350 491
rect 408 491 2008 538
rect 408 474 816 491
rect -58 457 -42 474
rect -858 441 -42 457
rect 800 457 816 474
rect 1600 474 2008 491
rect 2066 491 3666 538
rect 2066 474 2474 491
rect 1600 457 1616 474
rect 800 441 1616 457
rect 2458 457 2474 474
rect 3258 474 3666 491
rect 3724 491 5324 538
rect 3724 474 4132 491
rect 3258 457 3274 474
rect 2458 441 3274 457
rect 4116 457 4132 474
rect 4916 474 5324 491
rect 5382 491 6982 538
rect 5382 474 5790 491
rect 4916 457 4932 474
rect 4116 441 4932 457
rect 5774 457 5790 474
rect 6574 474 6982 491
rect 7040 491 8640 538
rect 7040 474 7448 491
rect 6574 457 6590 474
rect 5774 441 6590 457
rect 7432 457 7448 474
rect 8232 474 8640 491
rect 8698 491 10298 538
rect 8698 474 9106 491
rect 8232 457 8248 474
rect 7432 441 8248 457
rect 9090 457 9106 474
rect 9890 474 10298 491
rect 10356 491 11956 538
rect 10356 474 10764 491
rect 9890 457 9906 474
rect 9090 441 9906 457
rect 10748 457 10764 474
rect 11548 474 11956 491
rect 12014 491 13614 538
rect 12014 474 12422 491
rect 11548 457 11564 474
rect 10748 441 11564 457
rect 12406 457 12422 474
rect 13206 474 13614 491
rect 13672 491 15272 538
rect 13672 474 14080 491
rect 13206 457 13222 474
rect 12406 441 13222 457
rect 14064 457 14080 474
rect 14864 474 15272 491
rect 15330 491 16930 538
rect 15330 474 15738 491
rect 14864 457 14880 474
rect 14064 441 14880 457
rect 15722 457 15738 474
rect 16522 474 16930 491
rect 16988 491 18588 538
rect 16988 474 17396 491
rect 16522 457 16538 474
rect 15722 441 16538 457
rect 17380 457 17396 474
rect 18180 474 18588 491
rect 18646 491 20246 538
rect 18646 474 19054 491
rect 18180 457 18196 474
rect 17380 441 18196 457
rect 19038 457 19054 474
rect 19838 474 20246 491
rect 20304 491 21904 538
rect 20304 474 20712 491
rect 19838 457 19854 474
rect 19038 441 19854 457
rect 20696 457 20712 474
rect 21496 474 21904 491
rect 21962 491 23562 538
rect 21962 474 22370 491
rect 21496 457 21512 474
rect 20696 441 21512 457
rect 22354 457 22370 474
rect 23154 474 23562 491
rect 23620 491 25220 538
rect 23620 474 24028 491
rect 23154 457 23170 474
rect 22354 441 23170 457
rect 24012 457 24028 474
rect 24812 474 25220 491
rect 25278 491 26878 538
rect 25278 474 25686 491
rect 24812 457 24828 474
rect 24012 441 24828 457
rect 25670 457 25686 474
rect 26470 474 26878 491
rect 26936 491 28536 538
rect 26936 474 27344 491
rect 26470 457 26486 474
rect 25670 441 26486 457
rect 27328 457 27344 474
rect 28128 474 28536 491
rect 28594 491 30194 538
rect 28594 474 29002 491
rect 28128 457 28144 474
rect 27328 441 28144 457
rect 28986 457 29002 474
rect 29786 474 30194 491
rect 30252 491 31852 538
rect 30252 474 30660 491
rect 29786 457 29802 474
rect 28986 441 29802 457
rect 30644 457 30660 474
rect 31444 474 31852 491
rect 31910 491 33510 538
rect 31910 474 32318 491
rect 31444 457 31460 474
rect 30644 441 31460 457
rect 32302 457 32318 474
rect 33102 474 33510 491
rect 33102 457 33118 474
rect 32302 441 33118 457
rect 168 177 234 193
rect 168 143 184 177
rect 218 143 234 177
rect 168 127 234 143
rect 360 177 426 193
rect 360 143 376 177
rect 410 143 426 177
rect 360 127 426 143
rect 90 96 120 122
rect 186 96 216 127
rect 282 96 312 122
rect 378 96 408 127
rect 90 -335 120 -304
rect 186 -330 216 -304
rect 282 -335 312 -304
rect 378 -330 408 -304
rect 72 -351 138 -335
rect 72 -385 88 -351
rect 122 -385 138 -351
rect 72 -401 138 -385
rect 264 -351 330 -335
rect 264 -385 280 -351
rect 314 -385 330 -351
rect 264 -401 330 -385
rect 120 -476 186 -460
rect 120 -510 136 -476
rect 170 -510 186 -476
rect 42 -548 72 -522
rect 120 -526 186 -510
rect 312 -476 378 -460
rect 312 -510 328 -476
rect 362 -510 378 -476
rect 138 -548 168 -526
rect 234 -548 264 -522
rect 312 -526 378 -510
rect 330 -548 360 -526
rect 42 -770 72 -748
rect 24 -786 90 -770
rect 138 -774 168 -748
rect 234 -770 264 -748
rect 24 -820 40 -786
rect 74 -820 90 -786
rect 24 -836 90 -820
rect 216 -786 282 -770
rect 330 -774 360 -748
rect 216 -820 232 -786
rect 266 -820 282 -786
rect 216 -836 282 -820
<< polycont >>
rect -32346 16821 -31562 16855
rect -30688 16821 -29904 16855
rect -29030 16821 -28246 16855
rect -27372 16821 -26588 16855
rect -25714 16821 -24930 16855
rect -24056 16821 -23272 16855
rect -22398 16821 -21614 16855
rect -20740 16821 -19956 16855
rect -19082 16821 -18298 16855
rect -17424 16821 -16640 16855
rect -15766 16821 -14982 16855
rect -14108 16821 -13324 16855
rect -12450 16821 -11666 16855
rect -10792 16821 -10008 16855
rect -9134 16821 -8350 16855
rect -7476 16821 -6692 16855
rect -5818 16821 -5034 16855
rect -4160 16821 -3376 16855
rect -2502 16821 -1718 16855
rect -844 16821 -60 16855
rect 814 16821 1598 16855
rect 2472 16821 3256 16855
rect 4130 16821 4914 16855
rect 5788 16821 6572 16855
rect 7446 16821 8230 16855
rect 9104 16821 9888 16855
rect 10762 16821 11546 16855
rect 12420 16821 13204 16855
rect 14078 16821 14862 16855
rect 15736 16821 16520 16855
rect 17394 16821 18178 16855
rect 19052 16821 19836 16855
rect 20710 16821 21494 16855
rect 22368 16821 23152 16855
rect 24026 16821 24810 16855
rect 25684 16821 26468 16855
rect 27342 16821 28126 16855
rect 29000 16821 29784 16855
rect 30658 16821 31442 16855
rect 32316 16821 33100 16855
rect -32346 15293 -31562 15327
rect -30688 15293 -29904 15327
rect -29030 15293 -28246 15327
rect -27372 15293 -26588 15327
rect -25714 15293 -24930 15327
rect -24056 15293 -23272 15327
rect -22398 15293 -21614 15327
rect -20740 15293 -19956 15327
rect -19082 15293 -18298 15327
rect -17424 15293 -16640 15327
rect -15766 15293 -14982 15327
rect -14108 15293 -13324 15327
rect -12450 15293 -11666 15327
rect -10792 15293 -10008 15327
rect -9134 15293 -8350 15327
rect -7476 15293 -6692 15327
rect -5818 15293 -5034 15327
rect -4160 15293 -3376 15327
rect -2502 15293 -1718 15327
rect -844 15293 -60 15327
rect 814 15293 1598 15327
rect 2472 15293 3256 15327
rect 4130 15293 4914 15327
rect 5788 15293 6572 15327
rect 7446 15293 8230 15327
rect 9104 15293 9888 15327
rect 10762 15293 11546 15327
rect 12420 15293 13204 15327
rect 14078 15293 14862 15327
rect 15736 15293 16520 15327
rect 17394 15293 18178 15327
rect 19052 15293 19836 15327
rect 20710 15293 21494 15327
rect 22368 15293 23152 15327
rect 24026 15293 24810 15327
rect 25684 15293 26468 15327
rect 27342 15293 28126 15327
rect 29000 15293 29784 15327
rect 30658 15293 31442 15327
rect 32316 15293 33100 15327
rect -32346 15185 -31562 15219
rect -30688 15185 -29904 15219
rect -29030 15185 -28246 15219
rect -27372 15185 -26588 15219
rect -25714 15185 -24930 15219
rect -24056 15185 -23272 15219
rect -22398 15185 -21614 15219
rect -20740 15185 -19956 15219
rect -19082 15185 -18298 15219
rect -17424 15185 -16640 15219
rect -15766 15185 -14982 15219
rect -14108 15185 -13324 15219
rect -12450 15185 -11666 15219
rect -10792 15185 -10008 15219
rect -9134 15185 -8350 15219
rect -7476 15185 -6692 15219
rect -5818 15185 -5034 15219
rect -4160 15185 -3376 15219
rect -2502 15185 -1718 15219
rect -844 15185 -60 15219
rect 814 15185 1598 15219
rect 2472 15185 3256 15219
rect 4130 15185 4914 15219
rect 5788 15185 6572 15219
rect 7446 15185 8230 15219
rect 9104 15185 9888 15219
rect 10762 15185 11546 15219
rect 12420 15185 13204 15219
rect 14078 15185 14862 15219
rect 15736 15185 16520 15219
rect 17394 15185 18178 15219
rect 19052 15185 19836 15219
rect 20710 15185 21494 15219
rect 22368 15185 23152 15219
rect 24026 15185 24810 15219
rect 25684 15185 26468 15219
rect 27342 15185 28126 15219
rect 29000 15185 29784 15219
rect 30658 15185 31442 15219
rect 32316 15185 33100 15219
rect -32346 13657 -31562 13691
rect -30688 13657 -29904 13691
rect -29030 13657 -28246 13691
rect -27372 13657 -26588 13691
rect -25714 13657 -24930 13691
rect -24056 13657 -23272 13691
rect -22398 13657 -21614 13691
rect -20740 13657 -19956 13691
rect -19082 13657 -18298 13691
rect -17424 13657 -16640 13691
rect -15766 13657 -14982 13691
rect -14108 13657 -13324 13691
rect -12450 13657 -11666 13691
rect -10792 13657 -10008 13691
rect -9134 13657 -8350 13691
rect -7476 13657 -6692 13691
rect -5818 13657 -5034 13691
rect -4160 13657 -3376 13691
rect -2502 13657 -1718 13691
rect -844 13657 -60 13691
rect 814 13657 1598 13691
rect 2472 13657 3256 13691
rect 4130 13657 4914 13691
rect 5788 13657 6572 13691
rect 7446 13657 8230 13691
rect 9104 13657 9888 13691
rect 10762 13657 11546 13691
rect 12420 13657 13204 13691
rect 14078 13657 14862 13691
rect 15736 13657 16520 13691
rect 17394 13657 18178 13691
rect 19052 13657 19836 13691
rect 20710 13657 21494 13691
rect 22368 13657 23152 13691
rect 24026 13657 24810 13691
rect 25684 13657 26468 13691
rect 27342 13657 28126 13691
rect 29000 13657 29784 13691
rect 30658 13657 31442 13691
rect 32316 13657 33100 13691
rect -32344 13439 -31560 13473
rect -30686 13439 -29902 13473
rect -29028 13439 -28244 13473
rect -27370 13439 -26586 13473
rect -25712 13439 -24928 13473
rect -24054 13439 -23270 13473
rect -22396 13439 -21612 13473
rect -20738 13439 -19954 13473
rect -19080 13439 -18296 13473
rect -17422 13439 -16638 13473
rect -15764 13439 -14980 13473
rect -14106 13439 -13322 13473
rect -12448 13439 -11664 13473
rect -10790 13439 -10006 13473
rect -9132 13439 -8348 13473
rect -7474 13439 -6690 13473
rect -5816 13439 -5032 13473
rect -4158 13439 -3374 13473
rect -2500 13439 -1716 13473
rect -842 13439 -58 13473
rect 816 13439 1600 13473
rect 2474 13439 3258 13473
rect 4132 13439 4916 13473
rect 5790 13439 6574 13473
rect 7448 13439 8232 13473
rect 9106 13439 9890 13473
rect 10764 13439 11548 13473
rect 12422 13439 13206 13473
rect 14080 13439 14864 13473
rect 15738 13439 16522 13473
rect 17396 13439 18180 13473
rect 19054 13439 19838 13473
rect 20712 13439 21496 13473
rect 22370 13439 23154 13473
rect 24028 13439 24812 13473
rect 25686 13439 26470 13473
rect 27344 13439 28128 13473
rect 29002 13439 29786 13473
rect 30660 13439 31444 13473
rect 32318 13439 33102 13473
rect -32344 11911 -31560 11945
rect -30686 11911 -29902 11945
rect -29028 11911 -28244 11945
rect -27370 11911 -26586 11945
rect -25712 11911 -24928 11945
rect -24054 11911 -23270 11945
rect -22396 11911 -21612 11945
rect -20738 11911 -19954 11945
rect -19080 11911 -18296 11945
rect -17422 11911 -16638 11945
rect -15764 11911 -14980 11945
rect -14106 11911 -13322 11945
rect -12448 11911 -11664 11945
rect -10790 11911 -10006 11945
rect -9132 11911 -8348 11945
rect -7474 11911 -6690 11945
rect -5816 11911 -5032 11945
rect -4158 11911 -3374 11945
rect -2500 11911 -1716 11945
rect -842 11911 -58 11945
rect 816 11911 1600 11945
rect 2474 11911 3258 11945
rect 4132 11911 4916 11945
rect 5790 11911 6574 11945
rect 7448 11911 8232 11945
rect 9106 11911 9890 11945
rect 10764 11911 11548 11945
rect 12422 11911 13206 11945
rect 14080 11911 14864 11945
rect 15738 11911 16522 11945
rect 17396 11911 18180 11945
rect 19054 11911 19838 11945
rect 20712 11911 21496 11945
rect 22370 11911 23154 11945
rect 24028 11911 24812 11945
rect 25686 11911 26470 11945
rect 27344 11911 28128 11945
rect 29002 11911 29786 11945
rect 30660 11911 31444 11945
rect 32318 11911 33102 11945
rect -32344 11803 -31560 11837
rect -30686 11803 -29902 11837
rect -29028 11803 -28244 11837
rect -27370 11803 -26586 11837
rect -25712 11803 -24928 11837
rect -24054 11803 -23270 11837
rect -22396 11803 -21612 11837
rect -20738 11803 -19954 11837
rect -19080 11803 -18296 11837
rect -17422 11803 -16638 11837
rect -15764 11803 -14980 11837
rect -14106 11803 -13322 11837
rect -12448 11803 -11664 11837
rect -10790 11803 -10006 11837
rect -9132 11803 -8348 11837
rect -7474 11803 -6690 11837
rect -5816 11803 -5032 11837
rect -4158 11803 -3374 11837
rect -2500 11803 -1716 11837
rect -842 11803 -58 11837
rect 816 11803 1600 11837
rect 2474 11803 3258 11837
rect 4132 11803 4916 11837
rect 5790 11803 6574 11837
rect 7448 11803 8232 11837
rect 9106 11803 9890 11837
rect 10764 11803 11548 11837
rect 12422 11803 13206 11837
rect 14080 11803 14864 11837
rect 15738 11803 16522 11837
rect 17396 11803 18180 11837
rect 19054 11803 19838 11837
rect 20712 11803 21496 11837
rect 22370 11803 23154 11837
rect 24028 11803 24812 11837
rect 25686 11803 26470 11837
rect 27344 11803 28128 11837
rect 29002 11803 29786 11837
rect 30660 11803 31444 11837
rect 32318 11803 33102 11837
rect -32344 10275 -31560 10309
rect -30686 10275 -29902 10309
rect -29028 10275 -28244 10309
rect -27370 10275 -26586 10309
rect -25712 10275 -24928 10309
rect -24054 10275 -23270 10309
rect -22396 10275 -21612 10309
rect -20738 10275 -19954 10309
rect -19080 10275 -18296 10309
rect -17422 10275 -16638 10309
rect -15764 10275 -14980 10309
rect -14106 10275 -13322 10309
rect -12448 10275 -11664 10309
rect -10790 10275 -10006 10309
rect -9132 10275 -8348 10309
rect -7474 10275 -6690 10309
rect -5816 10275 -5032 10309
rect -4158 10275 -3374 10309
rect -2500 10275 -1716 10309
rect -842 10275 -58 10309
rect 816 10275 1600 10309
rect 2474 10275 3258 10309
rect 4132 10275 4916 10309
rect 5790 10275 6574 10309
rect 7448 10275 8232 10309
rect 9106 10275 9890 10309
rect 10764 10275 11548 10309
rect 12422 10275 13206 10309
rect 14080 10275 14864 10309
rect 15738 10275 16522 10309
rect 17396 10275 18180 10309
rect 19054 10275 19838 10309
rect 20712 10275 21496 10309
rect 22370 10275 23154 10309
rect 24028 10275 24812 10309
rect 25686 10275 26470 10309
rect 27344 10275 28128 10309
rect 29002 10275 29786 10309
rect 30660 10275 31444 10309
rect 32318 10275 33102 10309
rect -32344 10167 -31560 10201
rect -30686 10167 -29902 10201
rect -29028 10167 -28244 10201
rect -27370 10167 -26586 10201
rect -25712 10167 -24928 10201
rect -24054 10167 -23270 10201
rect -22396 10167 -21612 10201
rect -20738 10167 -19954 10201
rect -19080 10167 -18296 10201
rect -17422 10167 -16638 10201
rect -15764 10167 -14980 10201
rect -14106 10167 -13322 10201
rect -12448 10167 -11664 10201
rect -10790 10167 -10006 10201
rect -9132 10167 -8348 10201
rect -7474 10167 -6690 10201
rect -5816 10167 -5032 10201
rect -4158 10167 -3374 10201
rect -2500 10167 -1716 10201
rect -842 10167 -58 10201
rect 816 10167 1600 10201
rect 2474 10167 3258 10201
rect 4132 10167 4916 10201
rect 5790 10167 6574 10201
rect 7448 10167 8232 10201
rect 9106 10167 9890 10201
rect 10764 10167 11548 10201
rect 12422 10167 13206 10201
rect 14080 10167 14864 10201
rect 15738 10167 16522 10201
rect 17396 10167 18180 10201
rect 19054 10167 19838 10201
rect 20712 10167 21496 10201
rect 22370 10167 23154 10201
rect 24028 10167 24812 10201
rect 25686 10167 26470 10201
rect 27344 10167 28128 10201
rect 29002 10167 29786 10201
rect 30660 10167 31444 10201
rect 32318 10167 33102 10201
rect -32344 8639 -31560 8673
rect -30686 8639 -29902 8673
rect -29028 8639 -28244 8673
rect -27370 8639 -26586 8673
rect -25712 8639 -24928 8673
rect -24054 8639 -23270 8673
rect -22396 8639 -21612 8673
rect -20738 8639 -19954 8673
rect -19080 8639 -18296 8673
rect -17422 8639 -16638 8673
rect -15764 8639 -14980 8673
rect -14106 8639 -13322 8673
rect -12448 8639 -11664 8673
rect -10790 8639 -10006 8673
rect -9132 8639 -8348 8673
rect -7474 8639 -6690 8673
rect -5816 8639 -5032 8673
rect -4158 8639 -3374 8673
rect -2500 8639 -1716 8673
rect -842 8639 -58 8673
rect 816 8639 1600 8673
rect 2474 8639 3258 8673
rect 4132 8639 4916 8673
rect 5790 8639 6574 8673
rect 7448 8639 8232 8673
rect 9106 8639 9890 8673
rect 10764 8639 11548 8673
rect 12422 8639 13206 8673
rect 14080 8639 14864 8673
rect 15738 8639 16522 8673
rect 17396 8639 18180 8673
rect 19054 8639 19838 8673
rect 20712 8639 21496 8673
rect 22370 8639 23154 8673
rect 24028 8639 24812 8673
rect 25686 8639 26470 8673
rect 27344 8639 28128 8673
rect 29002 8639 29786 8673
rect 30660 8639 31444 8673
rect 32318 8639 33102 8673
rect -32344 8531 -31560 8565
rect -30686 8531 -29902 8565
rect -29028 8531 -28244 8565
rect -27370 8531 -26586 8565
rect -25712 8531 -24928 8565
rect -24054 8531 -23270 8565
rect -22396 8531 -21612 8565
rect -20738 8531 -19954 8565
rect -19080 8531 -18296 8565
rect -17422 8531 -16638 8565
rect -15764 8531 -14980 8565
rect -14106 8531 -13322 8565
rect -12448 8531 -11664 8565
rect -10790 8531 -10006 8565
rect -9132 8531 -8348 8565
rect -7474 8531 -6690 8565
rect -5816 8531 -5032 8565
rect -4158 8531 -3374 8565
rect -2500 8531 -1716 8565
rect -842 8531 -58 8565
rect 816 8531 1600 8565
rect 2474 8531 3258 8565
rect 4132 8531 4916 8565
rect 5790 8531 6574 8565
rect 7448 8531 8232 8565
rect 9106 8531 9890 8565
rect 10764 8531 11548 8565
rect 12422 8531 13206 8565
rect 14080 8531 14864 8565
rect 15738 8531 16522 8565
rect 17396 8531 18180 8565
rect 19054 8531 19838 8565
rect 20712 8531 21496 8565
rect 22370 8531 23154 8565
rect 24028 8531 24812 8565
rect 25686 8531 26470 8565
rect 27344 8531 28128 8565
rect 29002 8531 29786 8565
rect 30660 8531 31444 8565
rect 32318 8531 33102 8565
rect -32344 7003 -31560 7037
rect -30686 7003 -29902 7037
rect -29028 7003 -28244 7037
rect -27370 7003 -26586 7037
rect -25712 7003 -24928 7037
rect -24054 7003 -23270 7037
rect -22396 7003 -21612 7037
rect -20738 7003 -19954 7037
rect -19080 7003 -18296 7037
rect -17422 7003 -16638 7037
rect -15764 7003 -14980 7037
rect -14106 7003 -13322 7037
rect -12448 7003 -11664 7037
rect -10790 7003 -10006 7037
rect -9132 7003 -8348 7037
rect -7474 7003 -6690 7037
rect -5816 7003 -5032 7037
rect -4158 7003 -3374 7037
rect -2500 7003 -1716 7037
rect -842 7003 -58 7037
rect 816 7003 1600 7037
rect 2474 7003 3258 7037
rect 4132 7003 4916 7037
rect 5790 7003 6574 7037
rect 7448 7003 8232 7037
rect 9106 7003 9890 7037
rect 10764 7003 11548 7037
rect 12422 7003 13206 7037
rect 14080 7003 14864 7037
rect 15738 7003 16522 7037
rect 17396 7003 18180 7037
rect 19054 7003 19838 7037
rect 20712 7003 21496 7037
rect 22370 7003 23154 7037
rect 24028 7003 24812 7037
rect 25686 7003 26470 7037
rect 27344 7003 28128 7037
rect 29002 7003 29786 7037
rect 30660 7003 31444 7037
rect 32318 7003 33102 7037
rect -32344 6893 -31560 6927
rect -30686 6893 -29902 6927
rect -29028 6893 -28244 6927
rect -27370 6893 -26586 6927
rect -25712 6893 -24928 6927
rect -24054 6893 -23270 6927
rect -22396 6893 -21612 6927
rect -20738 6893 -19954 6927
rect -19080 6893 -18296 6927
rect -17422 6893 -16638 6927
rect -15764 6893 -14980 6927
rect -14106 6893 -13322 6927
rect -12448 6893 -11664 6927
rect -10790 6893 -10006 6927
rect -9132 6893 -8348 6927
rect -7474 6893 -6690 6927
rect -5816 6893 -5032 6927
rect -4158 6893 -3374 6927
rect -2500 6893 -1716 6927
rect -842 6893 -58 6927
rect 816 6893 1600 6927
rect 2474 6893 3258 6927
rect 4132 6893 4916 6927
rect 5790 6893 6574 6927
rect 7448 6893 8232 6927
rect 9106 6893 9890 6927
rect 10764 6893 11548 6927
rect 12422 6893 13206 6927
rect 14080 6893 14864 6927
rect 15738 6893 16522 6927
rect 17396 6893 18180 6927
rect 19054 6893 19838 6927
rect 20712 6893 21496 6927
rect 22370 6893 23154 6927
rect 24028 6893 24812 6927
rect 25686 6893 26470 6927
rect 27344 6893 28128 6927
rect 29002 6893 29786 6927
rect 30660 6893 31444 6927
rect 32318 6893 33102 6927
rect -32344 5365 -31560 5399
rect -30686 5365 -29902 5399
rect -29028 5365 -28244 5399
rect -27370 5365 -26586 5399
rect -25712 5365 -24928 5399
rect -24054 5365 -23270 5399
rect -22396 5365 -21612 5399
rect -20738 5365 -19954 5399
rect -19080 5365 -18296 5399
rect -17422 5365 -16638 5399
rect -15764 5365 -14980 5399
rect -14106 5365 -13322 5399
rect -12448 5365 -11664 5399
rect -10790 5365 -10006 5399
rect -9132 5365 -8348 5399
rect -7474 5365 -6690 5399
rect -5816 5365 -5032 5399
rect -4158 5365 -3374 5399
rect -2500 5365 -1716 5399
rect -842 5365 -58 5399
rect 816 5365 1600 5399
rect 2474 5365 3258 5399
rect 4132 5365 4916 5399
rect 5790 5365 6574 5399
rect 7448 5365 8232 5399
rect 9106 5365 9890 5399
rect 10764 5365 11548 5399
rect 12422 5365 13206 5399
rect 14080 5365 14864 5399
rect 15738 5365 16522 5399
rect 17396 5365 18180 5399
rect 19054 5365 19838 5399
rect 20712 5365 21496 5399
rect 22370 5365 23154 5399
rect 24028 5365 24812 5399
rect 25686 5365 26470 5399
rect 27344 5365 28128 5399
rect 29002 5365 29786 5399
rect 30660 5365 31444 5399
rect 32318 5365 33102 5399
rect -32344 5257 -31560 5291
rect -30686 5257 -29902 5291
rect -29028 5257 -28244 5291
rect -27370 5257 -26586 5291
rect -25712 5257 -24928 5291
rect -24054 5257 -23270 5291
rect -22396 5257 -21612 5291
rect -20738 5257 -19954 5291
rect -19080 5257 -18296 5291
rect -17422 5257 -16638 5291
rect -15764 5257 -14980 5291
rect -14106 5257 -13322 5291
rect -12448 5257 -11664 5291
rect -10790 5257 -10006 5291
rect -9132 5257 -8348 5291
rect -7474 5257 -6690 5291
rect -5816 5257 -5032 5291
rect -4158 5257 -3374 5291
rect -2500 5257 -1716 5291
rect -842 5257 -58 5291
rect 816 5257 1600 5291
rect 2474 5257 3258 5291
rect 4132 5257 4916 5291
rect 5790 5257 6574 5291
rect 7448 5257 8232 5291
rect 9106 5257 9890 5291
rect 10764 5257 11548 5291
rect 12422 5257 13206 5291
rect 14080 5257 14864 5291
rect 15738 5257 16522 5291
rect 17396 5257 18180 5291
rect 19054 5257 19838 5291
rect 20712 5257 21496 5291
rect 22370 5257 23154 5291
rect 24028 5257 24812 5291
rect 25686 5257 26470 5291
rect 27344 5257 28128 5291
rect 29002 5257 29786 5291
rect 30660 5257 31444 5291
rect 32318 5257 33102 5291
rect -32344 3729 -31560 3763
rect -30686 3729 -29902 3763
rect -29028 3729 -28244 3763
rect -27370 3729 -26586 3763
rect -25712 3729 -24928 3763
rect -24054 3729 -23270 3763
rect -22396 3729 -21612 3763
rect -20738 3729 -19954 3763
rect -19080 3729 -18296 3763
rect -17422 3729 -16638 3763
rect -15764 3729 -14980 3763
rect -14106 3729 -13322 3763
rect -12448 3729 -11664 3763
rect -10790 3729 -10006 3763
rect -9132 3729 -8348 3763
rect -7474 3729 -6690 3763
rect -5816 3729 -5032 3763
rect -4158 3729 -3374 3763
rect -2500 3729 -1716 3763
rect -842 3729 -58 3763
rect 816 3729 1600 3763
rect 2474 3729 3258 3763
rect 4132 3729 4916 3763
rect 5790 3729 6574 3763
rect 7448 3729 8232 3763
rect 9106 3729 9890 3763
rect 10764 3729 11548 3763
rect 12422 3729 13206 3763
rect 14080 3729 14864 3763
rect 15738 3729 16522 3763
rect 17396 3729 18180 3763
rect 19054 3729 19838 3763
rect 20712 3729 21496 3763
rect 22370 3729 23154 3763
rect 24028 3729 24812 3763
rect 25686 3729 26470 3763
rect 27344 3729 28128 3763
rect 29002 3729 29786 3763
rect 30660 3729 31444 3763
rect 32318 3729 33102 3763
rect -32344 3621 -31560 3655
rect -30686 3621 -29902 3655
rect -29028 3621 -28244 3655
rect -27370 3621 -26586 3655
rect -25712 3621 -24928 3655
rect -24054 3621 -23270 3655
rect -22396 3621 -21612 3655
rect -20738 3621 -19954 3655
rect -19080 3621 -18296 3655
rect -17422 3621 -16638 3655
rect -15764 3621 -14980 3655
rect -14106 3621 -13322 3655
rect -12448 3621 -11664 3655
rect -10790 3621 -10006 3655
rect -9132 3621 -8348 3655
rect -7474 3621 -6690 3655
rect -5816 3621 -5032 3655
rect -4158 3621 -3374 3655
rect -2500 3621 -1716 3655
rect -842 3621 -58 3655
rect 816 3621 1600 3655
rect 2474 3621 3258 3655
rect 4132 3621 4916 3655
rect 5790 3621 6574 3655
rect 7448 3621 8232 3655
rect 9106 3621 9890 3655
rect 10764 3621 11548 3655
rect 12422 3621 13206 3655
rect 14080 3621 14864 3655
rect 15738 3621 16522 3655
rect 17396 3621 18180 3655
rect 19054 3621 19838 3655
rect 20712 3621 21496 3655
rect 22370 3621 23154 3655
rect 24028 3621 24812 3655
rect 25686 3621 26470 3655
rect 27344 3621 28128 3655
rect 29002 3621 29786 3655
rect 30660 3621 31444 3655
rect 32318 3621 33102 3655
rect -32344 2093 -31560 2127
rect -30686 2093 -29902 2127
rect -29028 2093 -28244 2127
rect -27370 2093 -26586 2127
rect -25712 2093 -24928 2127
rect -24054 2093 -23270 2127
rect -22396 2093 -21612 2127
rect -20738 2093 -19954 2127
rect -19080 2093 -18296 2127
rect -17422 2093 -16638 2127
rect -15764 2093 -14980 2127
rect -14106 2093 -13322 2127
rect -12448 2093 -11664 2127
rect -10790 2093 -10006 2127
rect -9132 2093 -8348 2127
rect -7474 2093 -6690 2127
rect -5816 2093 -5032 2127
rect -4158 2093 -3374 2127
rect -2500 2093 -1716 2127
rect -842 2093 -58 2127
rect 816 2093 1600 2127
rect 2474 2093 3258 2127
rect 4132 2093 4916 2127
rect 5790 2093 6574 2127
rect 7448 2093 8232 2127
rect 9106 2093 9890 2127
rect 10764 2093 11548 2127
rect 12422 2093 13206 2127
rect 14080 2093 14864 2127
rect 15738 2093 16522 2127
rect 17396 2093 18180 2127
rect 19054 2093 19838 2127
rect 20712 2093 21496 2127
rect 22370 2093 23154 2127
rect 24028 2093 24812 2127
rect 25686 2093 26470 2127
rect 27344 2093 28128 2127
rect 29002 2093 29786 2127
rect 30660 2093 31444 2127
rect 32318 2093 33102 2127
rect -32344 1985 -31560 2019
rect -30686 1985 -29902 2019
rect -29028 1985 -28244 2019
rect -27370 1985 -26586 2019
rect -25712 1985 -24928 2019
rect -24054 1985 -23270 2019
rect -22396 1985 -21612 2019
rect -20738 1985 -19954 2019
rect -19080 1985 -18296 2019
rect -17422 1985 -16638 2019
rect -15764 1985 -14980 2019
rect -14106 1985 -13322 2019
rect -12448 1985 -11664 2019
rect -10790 1985 -10006 2019
rect -9132 1985 -8348 2019
rect -7474 1985 -6690 2019
rect -5816 1985 -5032 2019
rect -4158 1985 -3374 2019
rect -2500 1985 -1716 2019
rect -842 1985 -58 2019
rect 816 1985 1600 2019
rect 2474 1985 3258 2019
rect 4132 1985 4916 2019
rect 5790 1985 6574 2019
rect 7448 1985 8232 2019
rect 9106 1985 9890 2019
rect 10764 1985 11548 2019
rect 12422 1985 13206 2019
rect 14080 1985 14864 2019
rect 15738 1985 16522 2019
rect 17396 1985 18180 2019
rect 19054 1985 19838 2019
rect 20712 1985 21496 2019
rect 22370 1985 23154 2019
rect 24028 1985 24812 2019
rect 25686 1985 26470 2019
rect 27344 1985 28128 2019
rect 29002 1985 29786 2019
rect 30660 1985 31444 2019
rect 32318 1985 33102 2019
rect -32344 457 -31560 491
rect -30686 457 -29902 491
rect -29028 457 -28244 491
rect -27370 457 -26586 491
rect -25712 457 -24928 491
rect -24054 457 -23270 491
rect -22396 457 -21612 491
rect -20738 457 -19954 491
rect -19080 457 -18296 491
rect -17422 457 -16638 491
rect -15764 457 -14980 491
rect -14106 457 -13322 491
rect -12448 457 -11664 491
rect -10790 457 -10006 491
rect -9132 457 -8348 491
rect -7474 457 -6690 491
rect -5816 457 -5032 491
rect -4158 457 -3374 491
rect -2500 457 -1716 491
rect -842 457 -58 491
rect 816 457 1600 491
rect 2474 457 3258 491
rect 4132 457 4916 491
rect 5790 457 6574 491
rect 7448 457 8232 491
rect 9106 457 9890 491
rect 10764 457 11548 491
rect 12422 457 13206 491
rect 14080 457 14864 491
rect 15738 457 16522 491
rect 17396 457 18180 491
rect 19054 457 19838 491
rect 20712 457 21496 491
rect 22370 457 23154 491
rect 24028 457 24812 491
rect 25686 457 26470 491
rect 27344 457 28128 491
rect 29002 457 29786 491
rect 30660 457 31444 491
rect 32318 457 33102 491
rect 184 143 218 177
rect 376 143 410 177
rect 88 -385 122 -351
rect 280 -385 314 -351
rect 136 -510 170 -476
rect 328 -510 362 -476
rect 40 -820 74 -786
rect 232 -820 266 -786
<< locali >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -32416 16855 -31428 17046
rect -32416 16821 -32346 16855
rect -31562 16821 -31428 16855
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -32416 15327 -31428 16821
rect -30764 16855 -29776 17116
rect -30764 16821 -30688 16855
rect -29904 16821 -29776 16855
rect -32416 15293 -32346 15327
rect -31562 15293 -31428 15327
rect -32416 15219 -31428 15293
rect -32416 15185 -32346 15219
rect -31562 15185 -31428 15219
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -32416 13691 -31428 15185
rect -30764 15327 -29776 16821
rect -29158 16855 -28170 17046
rect -29158 16821 -29030 16855
rect -28246 16821 -28170 16855
rect -30764 15293 -30688 15327
rect -29904 15293 -29776 15327
rect -30764 15219 -29776 15293
rect -30764 15185 -30688 15219
rect -29904 15185 -29776 15219
rect -32416 13657 -32346 13691
rect -31562 13657 -31428 13691
rect -32416 13473 -31428 13657
rect -32416 13439 -32344 13473
rect -31560 13439 -31428 13473
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -32416 11945 -31428 13439
rect -30764 13691 -29776 15185
rect -29158 15327 -28170 16821
rect -27458 16855 -26470 17116
rect -27458 16821 -27372 16855
rect -26588 16821 -26470 16855
rect -29158 15293 -29030 15327
rect -28246 15293 -28170 15327
rect -29158 15219 -28170 15293
rect -29158 15185 -29030 15219
rect -28246 15185 -28170 15219
rect -30764 13657 -30688 13691
rect -29904 13657 -29776 13691
rect -30764 13473 -29776 13657
rect -30764 13439 -30686 13473
rect -29902 13439 -29776 13473
rect -32416 11911 -32344 11945
rect -31560 11911 -31428 11945
rect -32416 11837 -31428 11911
rect -32416 11803 -32344 11837
rect -31560 11803 -31428 11837
rect -34456 9946 -33510 11480
rect -32416 10309 -31428 11803
rect -30764 11945 -29776 13439
rect -29158 13691 -28170 15185
rect -27458 15327 -26470 16821
rect -25830 16855 -24842 17092
rect -25830 16821 -25714 16855
rect -24930 16821 -24842 16855
rect -27458 15293 -27372 15327
rect -26588 15293 -26470 15327
rect -27458 15219 -26470 15293
rect -27458 15185 -27372 15219
rect -26588 15185 -26470 15219
rect -29158 13657 -29030 13691
rect -28246 13657 -28170 13691
rect -29158 13473 -28170 13657
rect -29158 13439 -29028 13473
rect -28244 13439 -28170 13473
rect -30764 11911 -30686 11945
rect -29902 11911 -29776 11945
rect -30764 11837 -29776 11911
rect -30764 11803 -30686 11837
rect -29902 11803 -29776 11837
rect -32416 10275 -32344 10309
rect -31560 10275 -31428 10309
rect -32416 10201 -31428 10275
rect -32416 10167 -32344 10201
rect -31560 10167 -31428 10201
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -32416 8673 -31428 10167
rect -30764 10309 -29776 11803
rect -29158 11945 -28170 13439
rect -27458 13691 -26470 15185
rect -25830 15327 -24842 16821
rect -24154 16855 -23166 17116
rect -24154 16821 -24056 16855
rect -23272 16821 -23166 16855
rect -25830 15293 -25714 15327
rect -24930 15293 -24842 15327
rect -25830 15219 -24842 15293
rect -25830 15185 -25714 15219
rect -24930 15185 -24842 15219
rect -27458 13657 -27372 13691
rect -26588 13657 -26470 13691
rect -27458 13473 -26470 13657
rect -27458 13439 -27370 13473
rect -26586 13439 -26470 13473
rect -29158 11911 -29028 11945
rect -28244 11911 -28170 11945
rect -29158 11837 -28170 11911
rect -29158 11803 -29028 11837
rect -28244 11803 -28170 11837
rect -30764 10275 -30686 10309
rect -29902 10275 -29776 10309
rect -30764 10201 -29776 10275
rect -30764 10167 -30686 10201
rect -29902 10167 -29776 10201
rect -32416 8639 -32344 8673
rect -31560 8639 -31428 8673
rect -32416 8565 -31428 8639
rect -32416 8531 -32344 8565
rect -31560 8531 -31428 8565
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -32416 7037 -31428 8531
rect -30764 8673 -29776 10167
rect -29158 10309 -28170 11803
rect -27458 11945 -26470 13439
rect -25830 13691 -24842 15185
rect -24154 15327 -23166 16821
rect -22502 16855 -21514 17070
rect -22502 16821 -22398 16855
rect -21614 16821 -21514 16855
rect -24154 15293 -24056 15327
rect -23272 15293 -23166 15327
rect -24154 15219 -23166 15293
rect -24154 15185 -24056 15219
rect -23272 15185 -23166 15219
rect -25830 13657 -25714 13691
rect -24930 13657 -24842 13691
rect -25830 13473 -24842 13657
rect -25830 13439 -25712 13473
rect -24928 13439 -24842 13473
rect -27458 11911 -27370 11945
rect -26586 11911 -26470 11945
rect -27458 11837 -26470 11911
rect -27458 11803 -27370 11837
rect -26586 11803 -26470 11837
rect -29158 10275 -29028 10309
rect -28244 10275 -28170 10309
rect -29158 10201 -28170 10275
rect -29158 10167 -29028 10201
rect -28244 10167 -28170 10201
rect -30764 8639 -30686 8673
rect -29902 8639 -29776 8673
rect -30764 8565 -29776 8639
rect -30764 8531 -30686 8565
rect -29902 8531 -29776 8565
rect -32416 7003 -32344 7037
rect -31560 7003 -31428 7037
rect -32416 6927 -31428 7003
rect -32416 6893 -32344 6927
rect -31560 6893 -31428 6927
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -32416 5399 -31428 6893
rect -30764 7037 -29776 8531
rect -29158 8673 -28170 10167
rect -27458 10309 -26470 11803
rect -25830 11945 -24842 13439
rect -24154 13691 -23166 15185
rect -22502 15327 -21514 16821
rect -20872 16855 -19884 17092
rect -20872 16821 -20740 16855
rect -19956 16821 -19884 16855
rect -22502 15293 -22398 15327
rect -21614 15293 -21514 15327
rect -22502 15219 -21514 15293
rect -22502 15185 -22398 15219
rect -21614 15185 -21514 15219
rect -24154 13657 -24056 13691
rect -23272 13657 -23166 13691
rect -24154 13473 -23166 13657
rect -24154 13439 -24054 13473
rect -23270 13439 -23166 13473
rect -25830 11911 -25712 11945
rect -24928 11911 -24842 11945
rect -25830 11837 -24842 11911
rect -25830 11803 -25712 11837
rect -24928 11803 -24842 11837
rect -27458 10275 -27370 10309
rect -26586 10275 -26470 10309
rect -27458 10201 -26470 10275
rect -27458 10167 -27370 10201
rect -26586 10167 -26470 10201
rect -29158 8639 -29028 8673
rect -28244 8639 -28170 8673
rect -29158 8565 -28170 8639
rect -29158 8531 -29028 8565
rect -28244 8531 -28170 8565
rect -30764 7003 -30686 7037
rect -29902 7003 -29776 7037
rect -30764 6927 -29776 7003
rect -30764 6893 -30686 6927
rect -29902 6893 -29776 6927
rect -32416 5365 -32344 5399
rect -31560 5365 -31428 5399
rect -32416 5291 -31428 5365
rect -32416 5257 -32344 5291
rect -31560 5257 -31428 5291
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -32416 3763 -31428 5257
rect -30764 5399 -29776 6893
rect -29158 7037 -28170 8531
rect -27458 8673 -26470 10167
rect -25830 10309 -24842 11803
rect -24154 11945 -23166 13439
rect -22502 13691 -21514 15185
rect -20872 15327 -19884 16821
rect -19220 16855 -18232 17070
rect -19220 16821 -19082 16855
rect -18298 16821 -18232 16855
rect -20872 15293 -20740 15327
rect -19956 15293 -19884 15327
rect -20872 15219 -19884 15293
rect -20872 15185 -20740 15219
rect -19956 15185 -19884 15219
rect -22502 13657 -22398 13691
rect -21614 13657 -21514 13691
rect -22502 13473 -21514 13657
rect -22502 13439 -22396 13473
rect -21612 13439 -21514 13473
rect -24154 11911 -24054 11945
rect -23270 11911 -23166 11945
rect -24154 11837 -23166 11911
rect -24154 11803 -24054 11837
rect -23270 11803 -23166 11837
rect -25830 10275 -25712 10309
rect -24928 10275 -24842 10309
rect -25830 10201 -24842 10275
rect -25830 10167 -25712 10201
rect -24928 10167 -24842 10201
rect -27458 8639 -27370 8673
rect -26586 8639 -26470 8673
rect -27458 8565 -26470 8639
rect -27458 8531 -27370 8565
rect -26586 8531 -26470 8565
rect -29158 7003 -29028 7037
rect -28244 7003 -28170 7037
rect -29158 6927 -28170 7003
rect -29158 6893 -29028 6927
rect -28244 6893 -28170 6927
rect -30764 5365 -30686 5399
rect -29902 5365 -29776 5399
rect -30764 5291 -29776 5365
rect -30764 5257 -30686 5291
rect -29902 5257 -29776 5291
rect -32416 3729 -32344 3763
rect -31560 3729 -31428 3763
rect -32416 3655 -31428 3729
rect -32416 3621 -32344 3655
rect -31560 3621 -31428 3655
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -32416 2127 -31428 3621
rect -30764 3763 -29776 5257
rect -29158 5399 -28170 6893
rect -27458 7037 -26470 8531
rect -25830 8673 -24842 10167
rect -24154 10309 -23166 11803
rect -22502 11945 -21514 13439
rect -20872 13691 -19884 15185
rect -19220 15327 -18232 16821
rect -17520 16855 -16532 17092
rect -17520 16821 -17424 16855
rect -16640 16821 -16532 16855
rect -19220 15293 -19082 15327
rect -18298 15293 -18232 15327
rect -19220 15219 -18232 15293
rect -19220 15185 -19082 15219
rect -18298 15185 -18232 15219
rect -20872 13657 -20740 13691
rect -19956 13657 -19884 13691
rect -20872 13473 -19884 13657
rect -20872 13439 -20738 13473
rect -19954 13439 -19884 13473
rect -22502 11911 -22396 11945
rect -21612 11911 -21514 11945
rect -22502 11837 -21514 11911
rect -22502 11803 -22396 11837
rect -21612 11803 -21514 11837
rect -24154 10275 -24054 10309
rect -23270 10275 -23166 10309
rect -24154 10201 -23166 10275
rect -24154 10167 -24054 10201
rect -23270 10167 -23166 10201
rect -25830 8639 -25712 8673
rect -24928 8639 -24842 8673
rect -25830 8565 -24842 8639
rect -25830 8531 -25712 8565
rect -24928 8531 -24842 8565
rect -27458 7003 -27370 7037
rect -26586 7003 -26470 7037
rect -27458 6927 -26470 7003
rect -27458 6893 -27370 6927
rect -26586 6893 -26470 6927
rect -29158 5365 -29028 5399
rect -28244 5365 -28170 5399
rect -29158 5291 -28170 5365
rect -29158 5257 -29028 5291
rect -28244 5257 -28170 5291
rect -30764 3729 -30686 3763
rect -29902 3729 -29776 3763
rect -30764 3655 -29776 3729
rect -30764 3621 -30686 3655
rect -29902 3621 -29776 3655
rect -32416 2093 -32344 2127
rect -31560 2093 -31428 2127
rect -32416 2019 -31428 2093
rect -32416 1985 -32344 2019
rect -31560 1985 -31428 2019
rect -34456 388 -33510 1480
rect -32416 491 -31428 1985
rect -30764 2127 -29776 3621
rect -29158 3763 -28170 5257
rect -27458 5399 -26470 6893
rect -25830 7037 -24842 8531
rect -24154 8673 -23166 10167
rect -22502 10309 -21514 11803
rect -20872 11945 -19884 13439
rect -19220 13691 -18232 15185
rect -17520 15327 -16532 16821
rect -15962 16855 -14974 17092
rect -14214 16855 -13226 17116
rect -15962 16821 -15766 16855
rect -14982 16821 -14966 16855
rect -14214 16821 -14108 16855
rect -13324 16821 -13226 16855
rect -17520 15293 -17424 15327
rect -16640 15293 -16532 15327
rect -17520 15219 -16532 15293
rect -17520 15185 -17424 15219
rect -16640 15185 -16532 15219
rect -19220 13657 -19082 13691
rect -18298 13657 -18232 13691
rect -19220 13473 -18232 13657
rect -19220 13439 -19080 13473
rect -18296 13439 -18232 13473
rect -20872 11911 -20738 11945
rect -19954 11911 -19884 11945
rect -20872 11837 -19884 11911
rect -20872 11803 -20738 11837
rect -19954 11803 -19884 11837
rect -22502 10275 -22396 10309
rect -21612 10275 -21514 10309
rect -22502 10201 -21514 10275
rect -22502 10167 -22396 10201
rect -21612 10167 -21514 10201
rect -24154 8639 -24054 8673
rect -23270 8639 -23166 8673
rect -24154 8565 -23166 8639
rect -24154 8531 -24054 8565
rect -23270 8531 -23166 8565
rect -25830 7003 -25712 7037
rect -24928 7003 -24842 7037
rect -25830 6927 -24842 7003
rect -25830 6893 -25712 6927
rect -24928 6893 -24842 6927
rect -27458 5365 -27370 5399
rect -26586 5365 -26470 5399
rect -27458 5291 -26470 5365
rect -27458 5257 -27370 5291
rect -26586 5257 -26470 5291
rect -29158 3729 -29028 3763
rect -28244 3729 -28170 3763
rect -29158 3655 -28170 3729
rect -29158 3621 -29028 3655
rect -28244 3621 -28170 3655
rect -30764 2093 -30686 2127
rect -29902 2093 -29776 2127
rect -30764 2019 -29776 2093
rect -30764 1985 -30686 2019
rect -29902 1985 -29776 2019
rect -32416 457 -32344 491
rect -31560 457 -31428 491
rect -32416 426 -31428 457
rect -30764 491 -29776 1985
rect -29158 2127 -28170 3621
rect -27458 3763 -26470 5257
rect -25830 5399 -24842 6893
rect -24154 7037 -23166 8531
rect -22502 8673 -21514 10167
rect -20872 10309 -19884 11803
rect -19220 11945 -18232 13439
rect -17520 13691 -16532 15185
rect -15962 15327 -14974 16821
rect -14214 15327 -13226 16821
rect -12562 16855 -11574 17116
rect -12562 16821 -12450 16855
rect -11666 16821 -11574 16855
rect -15962 15293 -15766 15327
rect -14982 15293 -14966 15327
rect -14214 15293 -14108 15327
rect -13324 15293 -13226 15327
rect -15962 15219 -14974 15293
rect -14214 15219 -13226 15293
rect -15962 15185 -15766 15219
rect -14982 15185 -14966 15219
rect -14214 15185 -14108 15219
rect -13324 15185 -13226 15219
rect -17520 13657 -17424 13691
rect -16640 13657 -16532 13691
rect -17520 13473 -16532 13657
rect -17520 13439 -17422 13473
rect -16638 13439 -16532 13473
rect -19220 11911 -19080 11945
rect -18296 11911 -18232 11945
rect -19220 11837 -18232 11911
rect -19220 11803 -19080 11837
rect -18296 11803 -18232 11837
rect -20872 10275 -20738 10309
rect -19954 10275 -19884 10309
rect -20872 10201 -19884 10275
rect -20872 10167 -20738 10201
rect -19954 10167 -19884 10201
rect -22502 8639 -22396 8673
rect -21612 8639 -21514 8673
rect -22502 8565 -21514 8639
rect -22502 8531 -22396 8565
rect -21612 8531 -21514 8565
rect -24154 7003 -24054 7037
rect -23270 7003 -23166 7037
rect -24154 6927 -23166 7003
rect -24154 6893 -24054 6927
rect -23270 6893 -23166 6927
rect -25830 5365 -25712 5399
rect -24928 5365 -24842 5399
rect -25830 5291 -24842 5365
rect -25830 5257 -25712 5291
rect -24928 5257 -24842 5291
rect -27458 3729 -27370 3763
rect -26586 3729 -26470 3763
rect -27458 3655 -26470 3729
rect -27458 3621 -27370 3655
rect -26586 3621 -26470 3655
rect -29158 2093 -29028 2127
rect -28244 2093 -28170 2127
rect -29158 2019 -28170 2093
rect -29158 1985 -29028 2019
rect -28244 1985 -28170 2019
rect -30764 457 -30686 491
rect -29902 457 -29776 491
rect -30764 426 -29776 457
rect -29158 491 -28170 1985
rect -27458 2127 -26470 3621
rect -25830 3763 -24842 5257
rect -24154 5399 -23166 6893
rect -22502 7037 -21514 8531
rect -20872 8673 -19884 10167
rect -19220 10309 -18232 11803
rect -17520 11945 -16532 13439
rect -15962 13691 -14974 15185
rect -14214 13691 -13226 15185
rect -12562 15327 -11574 16821
rect -10932 16855 -9944 17116
rect -10932 16821 -10792 16855
rect -10008 16821 -9944 16855
rect -12562 15293 -12450 15327
rect -11666 15293 -11574 15327
rect -12562 15219 -11574 15293
rect -12562 15185 -12450 15219
rect -11666 15185 -11574 15219
rect -15962 13657 -15766 13691
rect -14982 13657 -14966 13691
rect -14214 13657 -14108 13691
rect -13324 13657 -13226 13691
rect -15962 13473 -14974 13657
rect -14214 13473 -13226 13657
rect -15962 13439 -15764 13473
rect -14980 13439 -14964 13473
rect -14214 13439 -14106 13473
rect -13322 13439 -13226 13473
rect -17520 11911 -17422 11945
rect -16638 11911 -16532 11945
rect -17520 11837 -16532 11911
rect -17520 11803 -17422 11837
rect -16638 11803 -16532 11837
rect -19220 10275 -19080 10309
rect -18296 10275 -18232 10309
rect -19220 10201 -18232 10275
rect -19220 10167 -19080 10201
rect -18296 10167 -18232 10201
rect -20872 8639 -20738 8673
rect -19954 8639 -19884 8673
rect -20872 8565 -19884 8639
rect -20872 8531 -20738 8565
rect -19954 8531 -19884 8565
rect -22502 7003 -22396 7037
rect -21612 7003 -21514 7037
rect -22502 6927 -21514 7003
rect -22502 6893 -22396 6927
rect -21612 6893 -21514 6927
rect -24154 5365 -24054 5399
rect -23270 5365 -23166 5399
rect -24154 5291 -23166 5365
rect -24154 5257 -24054 5291
rect -23270 5257 -23166 5291
rect -25830 3729 -25712 3763
rect -24928 3729 -24842 3763
rect -25830 3655 -24842 3729
rect -25830 3621 -25712 3655
rect -24928 3621 -24842 3655
rect -27458 2093 -27370 2127
rect -26586 2093 -26470 2127
rect -27458 2019 -26470 2093
rect -27458 1985 -27370 2019
rect -26586 1985 -26470 2019
rect -29158 457 -29028 491
rect -28244 457 -28170 491
rect -29158 426 -28170 457
rect -27458 491 -26470 1985
rect -25830 2127 -24842 3621
rect -24154 3763 -23166 5257
rect -22502 5399 -21514 6893
rect -20872 7037 -19884 8531
rect -19220 8673 -18232 10167
rect -17520 10309 -16532 11803
rect -15962 11945 -14974 13439
rect -14214 11945 -13226 13439
rect -12562 13691 -11574 15185
rect -10932 15327 -9944 16821
rect -9254 16855 -8266 17116
rect -9254 16821 -9134 16855
rect -8350 16821 -8266 16855
rect -10932 15293 -10792 15327
rect -10008 15293 -9944 15327
rect -10932 15219 -9944 15293
rect -10932 15185 -10792 15219
rect -10008 15185 -9944 15219
rect -12562 13657 -12450 13691
rect -11666 13657 -11574 13691
rect -12562 13473 -11574 13657
rect -12562 13439 -12448 13473
rect -11664 13439 -11574 13473
rect -15962 11911 -15764 11945
rect -14980 11911 -14964 11945
rect -14214 11911 -14106 11945
rect -13322 11911 -13226 11945
rect -15962 11837 -14974 11911
rect -14214 11837 -13226 11911
rect -15962 11803 -15764 11837
rect -14980 11803 -14964 11837
rect -14214 11803 -14106 11837
rect -13322 11803 -13226 11837
rect -17520 10275 -17422 10309
rect -16638 10275 -16532 10309
rect -17520 10201 -16532 10275
rect -17520 10167 -17422 10201
rect -16638 10167 -16532 10201
rect -19220 8639 -19080 8673
rect -18296 8639 -18232 8673
rect -19220 8565 -18232 8639
rect -19220 8531 -19080 8565
rect -18296 8531 -18232 8565
rect -20872 7003 -20738 7037
rect -19954 7003 -19884 7037
rect -20872 6927 -19884 7003
rect -20872 6893 -20738 6927
rect -19954 6893 -19884 6927
rect -22502 5365 -22396 5399
rect -21612 5365 -21514 5399
rect -22502 5291 -21514 5365
rect -22502 5257 -22396 5291
rect -21612 5257 -21514 5291
rect -24154 3729 -24054 3763
rect -23270 3729 -23166 3763
rect -24154 3655 -23166 3729
rect -24154 3621 -24054 3655
rect -23270 3621 -23166 3655
rect -25830 2093 -25712 2127
rect -24928 2093 -24842 2127
rect -25830 2019 -24842 2093
rect -25830 1985 -25712 2019
rect -24928 1985 -24842 2019
rect -27458 457 -27370 491
rect -26586 457 -26470 491
rect -27458 426 -26470 457
rect -25830 491 -24842 1985
rect -24154 2127 -23166 3621
rect -22502 3763 -21514 5257
rect -20872 5399 -19884 6893
rect -19220 7037 -18232 8531
rect -17520 8673 -16532 10167
rect -15962 10309 -14974 11803
rect -14214 10309 -13226 11803
rect -12562 11945 -11574 13439
rect -10932 13691 -9944 15185
rect -9254 15327 -8266 16821
rect -7556 16855 -6568 17092
rect -7556 16821 -7476 16855
rect -6692 16821 -6568 16855
rect -9254 15293 -9134 15327
rect -8350 15293 -8266 15327
rect -9254 15219 -8266 15293
rect -9254 15185 -9134 15219
rect -8350 15185 -8266 15219
rect -10932 13657 -10792 13691
rect -10008 13657 -9944 13691
rect -10932 13473 -9944 13657
rect -10932 13439 -10790 13473
rect -10006 13439 -9944 13473
rect -12562 11911 -12448 11945
rect -11664 11911 -11574 11945
rect -12562 11837 -11574 11911
rect -12562 11803 -12448 11837
rect -11664 11803 -11574 11837
rect -15962 10275 -15764 10309
rect -14980 10275 -14964 10309
rect -14214 10275 -14106 10309
rect -13322 10275 -13226 10309
rect -15962 10201 -14974 10275
rect -14214 10201 -13226 10275
rect -15962 10167 -15764 10201
rect -14980 10167 -14964 10201
rect -14214 10167 -14106 10201
rect -13322 10167 -13226 10201
rect -17520 8639 -17422 8673
rect -16638 8639 -16532 8673
rect -17520 8565 -16532 8639
rect -17520 8531 -17422 8565
rect -16638 8531 -16532 8565
rect -19220 7003 -19080 7037
rect -18296 7003 -18232 7037
rect -19220 6927 -18232 7003
rect -19220 6893 -19080 6927
rect -18296 6893 -18232 6927
rect -20872 5365 -20738 5399
rect -19954 5365 -19884 5399
rect -20872 5291 -19884 5365
rect -20872 5257 -20738 5291
rect -19954 5257 -19884 5291
rect -22502 3729 -22396 3763
rect -21612 3729 -21514 3763
rect -22502 3655 -21514 3729
rect -22502 3621 -22396 3655
rect -21612 3621 -21514 3655
rect -24154 2093 -24054 2127
rect -23270 2093 -23166 2127
rect -24154 2019 -23166 2093
rect -24154 1985 -24054 2019
rect -23270 1985 -23166 2019
rect -25830 457 -25712 491
rect -24928 457 -24842 491
rect -25830 426 -24842 457
rect -24154 491 -23166 1985
rect -22502 2127 -21514 3621
rect -20872 3763 -19884 5257
rect -19220 5399 -18232 6893
rect -17520 7037 -16532 8531
rect -15962 8673 -14974 10167
rect -14214 8673 -13226 10167
rect -12562 10309 -11574 11803
rect -10932 11945 -9944 13439
rect -9254 13691 -8266 15185
rect -7556 15327 -6568 16821
rect -5926 16855 -4938 17140
rect -5926 16821 -5818 16855
rect -5034 16821 -4938 16855
rect -7556 15293 -7476 15327
rect -6692 15293 -6568 15327
rect -7556 15219 -6568 15293
rect -7556 15185 -7476 15219
rect -6692 15185 -6568 15219
rect -9254 13657 -9134 13691
rect -8350 13657 -8266 13691
rect -9254 13473 -8266 13657
rect -9254 13439 -9132 13473
rect -8348 13439 -8266 13473
rect -10932 11911 -10790 11945
rect -10006 11911 -9944 11945
rect -10932 11837 -9944 11911
rect -10932 11803 -10790 11837
rect -10006 11803 -9944 11837
rect -12562 10275 -12448 10309
rect -11664 10275 -11574 10309
rect -12562 10201 -11574 10275
rect -12562 10167 -12448 10201
rect -11664 10167 -11574 10201
rect -15962 8639 -15764 8673
rect -14980 8639 -14964 8673
rect -14214 8639 -14106 8673
rect -13322 8639 -13226 8673
rect -15962 8565 -14974 8639
rect -14214 8565 -13226 8639
rect -15962 8531 -15764 8565
rect -14980 8531 -14964 8565
rect -14214 8531 -14106 8565
rect -13322 8531 -13226 8565
rect -17520 7003 -17422 7037
rect -16638 7003 -16532 7037
rect -17520 6927 -16532 7003
rect -17520 6893 -17422 6927
rect -16638 6893 -16532 6927
rect -19220 5365 -19080 5399
rect -18296 5365 -18232 5399
rect -19220 5291 -18232 5365
rect -19220 5257 -19080 5291
rect -18296 5257 -18232 5291
rect -20872 3729 -20738 3763
rect -19954 3729 -19884 3763
rect -20872 3655 -19884 3729
rect -20872 3621 -20738 3655
rect -19954 3621 -19884 3655
rect -22502 2093 -22396 2127
rect -21612 2093 -21514 2127
rect -22502 2019 -21514 2093
rect -22502 1985 -22396 2019
rect -21612 1985 -21514 2019
rect -24154 457 -24054 491
rect -23270 457 -23166 491
rect -24154 426 -23166 457
rect -22502 491 -21514 1985
rect -20872 2127 -19884 3621
rect -19220 3763 -18232 5257
rect -17520 5399 -16532 6893
rect -15962 7037 -14974 8531
rect -14214 7037 -13226 8531
rect -12562 8673 -11574 10167
rect -10932 10309 -9944 11803
rect -9254 11945 -8266 13439
rect -7556 13691 -6568 15185
rect -5926 15327 -4938 16821
rect -4250 16855 -3262 17116
rect -4250 16821 -4160 16855
rect -3376 16821 -3262 16855
rect -5926 15293 -5818 15327
rect -5034 15293 -4938 15327
rect -5926 15219 -4938 15293
rect -5926 15185 -5818 15219
rect -5034 15185 -4938 15219
rect -7556 13657 -7476 13691
rect -6692 13657 -6568 13691
rect -7556 13473 -6568 13657
rect -7556 13439 -7474 13473
rect -6690 13439 -6568 13473
rect -9254 11911 -9132 11945
rect -8348 11911 -8266 11945
rect -9254 11837 -8266 11911
rect -9254 11803 -9132 11837
rect -8348 11803 -8266 11837
rect -10932 10275 -10790 10309
rect -10006 10275 -9944 10309
rect -10932 10201 -9944 10275
rect -10932 10167 -10790 10201
rect -10006 10167 -9944 10201
rect -12562 8639 -12448 8673
rect -11664 8639 -11574 8673
rect -12562 8565 -11574 8639
rect -12562 8531 -12448 8565
rect -11664 8531 -11574 8565
rect -15962 7003 -15764 7037
rect -14980 7003 -14964 7037
rect -14214 7003 -14106 7037
rect -13322 7003 -13226 7037
rect -15962 6927 -14974 7003
rect -14214 6927 -13226 7003
rect -15962 6893 -15764 6927
rect -14980 6893 -14964 6927
rect -14214 6893 -14106 6927
rect -13322 6893 -13226 6927
rect -17520 5365 -17422 5399
rect -16638 5365 -16532 5399
rect -17520 5291 -16532 5365
rect -17520 5257 -17422 5291
rect -16638 5257 -16532 5291
rect -19220 3729 -19080 3763
rect -18296 3729 -18232 3763
rect -19220 3655 -18232 3729
rect -19220 3621 -19080 3655
rect -18296 3621 -18232 3655
rect -20872 2093 -20738 2127
rect -19954 2093 -19884 2127
rect -20872 2019 -19884 2093
rect -20872 1985 -20738 2019
rect -19954 1985 -19884 2019
rect -22502 457 -22396 491
rect -21612 457 -21514 491
rect -22502 426 -21514 457
rect -20872 491 -19884 1985
rect -19220 2127 -18232 3621
rect -17520 3763 -16532 5257
rect -15962 5399 -14974 6893
rect -14214 5399 -13226 6893
rect -12562 7037 -11574 8531
rect -10932 8673 -9944 10167
rect -9254 10309 -8266 11803
rect -7556 11945 -6568 13439
rect -5926 13691 -4938 15185
rect -4250 15327 -3262 16821
rect -2598 16855 -1610 17140
rect -2598 16821 -2502 16855
rect -1718 16821 -1610 16855
rect -4250 15293 -4160 15327
rect -3376 15293 -3262 15327
rect -4250 15219 -3262 15293
rect -4250 15185 -4160 15219
rect -3376 15185 -3262 15219
rect -5926 13657 -5818 13691
rect -5034 13657 -4938 13691
rect -5926 13473 -4938 13657
rect -5926 13439 -5816 13473
rect -5032 13439 -4938 13473
rect -7556 11911 -7474 11945
rect -6690 11911 -6568 11945
rect -7556 11837 -6568 11911
rect -7556 11803 -7474 11837
rect -6690 11803 -6568 11837
rect -9254 10275 -9132 10309
rect -8348 10275 -8266 10309
rect -9254 10201 -8266 10275
rect -9254 10167 -9132 10201
rect -8348 10167 -8266 10201
rect -10932 8639 -10790 8673
rect -10006 8639 -9944 8673
rect -10932 8565 -9944 8639
rect -10932 8531 -10790 8565
rect -10006 8531 -9944 8565
rect -12562 7003 -12448 7037
rect -11664 7003 -11574 7037
rect -12562 6927 -11574 7003
rect -12562 6893 -12448 6927
rect -11664 6893 -11574 6927
rect -15962 5365 -15764 5399
rect -14980 5365 -14964 5399
rect -14214 5365 -14106 5399
rect -13322 5365 -13226 5399
rect -15962 5291 -14974 5365
rect -14214 5291 -13226 5365
rect -15962 5257 -15764 5291
rect -14980 5257 -14964 5291
rect -14214 5257 -14106 5291
rect -13322 5257 -13226 5291
rect -17520 3729 -17422 3763
rect -16638 3729 -16532 3763
rect -17520 3655 -16532 3729
rect -17520 3621 -17422 3655
rect -16638 3621 -16532 3655
rect -19220 2093 -19080 2127
rect -18296 2093 -18232 2127
rect -19220 2019 -18232 2093
rect -19220 1985 -19080 2019
rect -18296 1985 -18232 2019
rect -20872 457 -20738 491
rect -19954 457 -19884 491
rect -20872 426 -19884 457
rect -19220 491 -18232 1985
rect -17520 2127 -16532 3621
rect -15962 3763 -14974 5257
rect -14214 3763 -13226 5257
rect -12562 5399 -11574 6893
rect -10932 7037 -9944 8531
rect -9254 8673 -8266 10167
rect -7556 10309 -6568 11803
rect -5926 11945 -4938 13439
rect -4250 13691 -3262 15185
rect -2598 15327 -1610 16821
rect -968 16855 20 17116
rect -968 16821 -844 16855
rect -60 16821 20 16855
rect -2598 15293 -2502 15327
rect -1718 15293 -1610 15327
rect -2598 15219 -1610 15293
rect -2598 15185 -2502 15219
rect -1718 15185 -1610 15219
rect -4250 13657 -4160 13691
rect -3376 13657 -3262 13691
rect -4250 13473 -3262 13657
rect -4250 13439 -4158 13473
rect -3374 13439 -3262 13473
rect -5926 11911 -5816 11945
rect -5032 11911 -4938 11945
rect -5926 11837 -4938 11911
rect -5926 11803 -5816 11837
rect -5032 11803 -4938 11837
rect -7556 10275 -7474 10309
rect -6690 10275 -6568 10309
rect -7556 10201 -6568 10275
rect -7556 10167 -7474 10201
rect -6690 10167 -6568 10201
rect -9254 8639 -9132 8673
rect -8348 8639 -8266 8673
rect -9254 8565 -8266 8639
rect -9254 8531 -9132 8565
rect -8348 8531 -8266 8565
rect -10932 7003 -10790 7037
rect -10006 7003 -9944 7037
rect -10932 6927 -9944 7003
rect -10932 6893 -10790 6927
rect -10006 6893 -9944 6927
rect -12562 5365 -12448 5399
rect -11664 5365 -11574 5399
rect -12562 5291 -11574 5365
rect -12562 5257 -12448 5291
rect -11664 5257 -11574 5291
rect -15962 3729 -15764 3763
rect -14980 3729 -14964 3763
rect -14214 3729 -14106 3763
rect -13322 3729 -13226 3763
rect -15962 3655 -14974 3729
rect -14214 3655 -13226 3729
rect -15962 3621 -15764 3655
rect -14980 3621 -14964 3655
rect -14214 3621 -14106 3655
rect -13322 3621 -13226 3655
rect -17520 2093 -17422 2127
rect -16638 2093 -16532 2127
rect -17520 2019 -16532 2093
rect -17520 1985 -17422 2019
rect -16638 1985 -16532 2019
rect -19220 457 -19080 491
rect -18296 457 -18232 491
rect -19220 426 -18232 457
rect -17520 491 -16532 1985
rect -15962 2127 -14974 3621
rect -14214 2127 -13226 3621
rect -12562 3763 -11574 5257
rect -10932 5399 -9944 6893
rect -9254 7037 -8266 8531
rect -7556 8673 -6568 10167
rect -5926 10309 -4938 11803
rect -4250 11945 -3262 13439
rect -2598 13691 -1610 15185
rect -968 15327 20 16821
rect 754 16855 1742 17116
rect 754 16821 814 16855
rect 1598 16821 1742 16855
rect -968 15293 -844 15327
rect -60 15293 20 15327
rect -968 15219 20 15293
rect -968 15185 -844 15219
rect -60 15185 20 15219
rect -2598 13657 -2502 13691
rect -1718 13657 -1610 13691
rect -2598 13473 -1610 13657
rect -2598 13439 -2500 13473
rect -1716 13439 -1610 13473
rect -4250 11911 -4158 11945
rect -3374 11911 -3262 11945
rect -4250 11837 -3262 11911
rect -4250 11803 -4158 11837
rect -3374 11803 -3262 11837
rect -5926 10275 -5816 10309
rect -5032 10275 -4938 10309
rect -5926 10201 -4938 10275
rect -5926 10167 -5816 10201
rect -5032 10167 -4938 10201
rect -7556 8639 -7474 8673
rect -6690 8639 -6568 8673
rect -7556 8565 -6568 8639
rect -7556 8531 -7474 8565
rect -6690 8531 -6568 8565
rect -9254 7003 -9132 7037
rect -8348 7003 -8266 7037
rect -9254 6927 -8266 7003
rect -9254 6893 -9132 6927
rect -8348 6893 -8266 6927
rect -10932 5365 -10790 5399
rect -10006 5365 -9944 5399
rect -10932 5291 -9944 5365
rect -10932 5257 -10790 5291
rect -10006 5257 -9944 5291
rect -12562 3729 -12448 3763
rect -11664 3729 -11574 3763
rect -12562 3655 -11574 3729
rect -12562 3621 -12448 3655
rect -11664 3621 -11574 3655
rect -15962 2093 -15764 2127
rect -14980 2093 -14964 2127
rect -14214 2093 -14106 2127
rect -13322 2093 -13226 2127
rect -15962 2019 -14974 2093
rect -14214 2019 -13226 2093
rect -15962 1985 -15764 2019
rect -14980 1985 -14964 2019
rect -14214 1985 -14106 2019
rect -13322 1985 -13226 2019
rect -17520 457 -17422 491
rect -16638 457 -16532 491
rect -17520 426 -16532 457
rect -15962 491 -14974 1985
rect -14214 491 -13226 1985
rect -12562 2127 -11574 3621
rect -10932 3763 -9944 5257
rect -9254 5399 -8266 6893
rect -7556 7037 -6568 8531
rect -5926 8673 -4938 10167
rect -4250 10309 -3262 11803
rect -2598 11945 -1610 13439
rect -968 13691 20 15185
rect 754 15327 1742 16821
rect 2360 16855 3348 17116
rect 2360 16821 2472 16855
rect 3256 16821 3348 16855
rect 754 15293 814 15327
rect 1598 15293 1742 15327
rect 754 15219 1742 15293
rect 754 15185 814 15219
rect 1598 15185 1742 15219
rect -968 13657 -844 13691
rect -60 13657 20 13691
rect -968 13473 20 13657
rect -968 13439 -842 13473
rect -58 13439 20 13473
rect -2598 11911 -2500 11945
rect -1716 11911 -1610 11945
rect -2598 11837 -1610 11911
rect -2598 11803 -2500 11837
rect -1716 11803 -1610 11837
rect -4250 10275 -4158 10309
rect -3374 10275 -3262 10309
rect -4250 10201 -3262 10275
rect -4250 10167 -4158 10201
rect -3374 10167 -3262 10201
rect -5926 8639 -5816 8673
rect -5032 8639 -4938 8673
rect -5926 8565 -4938 8639
rect -5926 8531 -5816 8565
rect -5032 8531 -4938 8565
rect -7556 7003 -7474 7037
rect -6690 7003 -6568 7037
rect -7556 6927 -6568 7003
rect -7556 6893 -7474 6927
rect -6690 6893 -6568 6927
rect -9254 5365 -9132 5399
rect -8348 5365 -8266 5399
rect -9254 5291 -8266 5365
rect -9254 5257 -9132 5291
rect -8348 5257 -8266 5291
rect -10932 3729 -10790 3763
rect -10006 3729 -9944 3763
rect -10932 3655 -9944 3729
rect -10932 3621 -10790 3655
rect -10006 3621 -9944 3655
rect -12562 2093 -12448 2127
rect -11664 2093 -11574 2127
rect -12562 2019 -11574 2093
rect -12562 1985 -12448 2019
rect -11664 1985 -11574 2019
rect -15962 457 -15764 491
rect -14980 457 -14964 491
rect -15962 426 -14964 457
rect -14214 457 -14106 491
rect -13322 457 -13226 491
rect -14214 426 -13226 457
rect -12562 491 -11574 1985
rect -10932 2127 -9944 3621
rect -9254 3763 -8266 5257
rect -7556 5399 -6568 6893
rect -5926 7037 -4938 8531
rect -4250 8673 -3262 10167
rect -2598 10309 -1610 11803
rect -968 11945 20 13439
rect 754 13691 1742 15185
rect 2360 15327 3348 16821
rect 4060 16855 5048 17116
rect 4060 16821 4130 16855
rect 4914 16821 5048 16855
rect 2360 15293 2472 15327
rect 3256 15293 3348 15327
rect 2360 15219 3348 15293
rect 2360 15185 2472 15219
rect 3256 15185 3348 15219
rect 754 13657 814 13691
rect 1598 13657 1742 13691
rect 754 13473 1742 13657
rect 754 13439 816 13473
rect 1600 13439 1742 13473
rect -968 11911 -842 11945
rect -58 11911 20 11945
rect -968 11837 20 11911
rect -968 11803 -842 11837
rect -58 11803 20 11837
rect -2598 10275 -2500 10309
rect -1716 10275 -1610 10309
rect -2598 10201 -1610 10275
rect -2598 10167 -2500 10201
rect -1716 10167 -1610 10201
rect -4250 8639 -4158 8673
rect -3374 8639 -3262 8673
rect -4250 8565 -3262 8639
rect -4250 8531 -4158 8565
rect -3374 8531 -3262 8565
rect -5926 7003 -5816 7037
rect -5032 7003 -4938 7037
rect -5926 6927 -4938 7003
rect -5926 6893 -5816 6927
rect -5032 6893 -4938 6927
rect -7556 5365 -7474 5399
rect -6690 5365 -6568 5399
rect -7556 5291 -6568 5365
rect -7556 5257 -7474 5291
rect -6690 5257 -6568 5291
rect -9254 3729 -9132 3763
rect -8348 3729 -8266 3763
rect -9254 3655 -8266 3729
rect -9254 3621 -9132 3655
rect -8348 3621 -8266 3655
rect -10932 2093 -10790 2127
rect -10006 2093 -9944 2127
rect -10932 2019 -9944 2093
rect -10932 1985 -10790 2019
rect -10006 1985 -9944 2019
rect -12562 457 -12448 491
rect -11664 457 -11574 491
rect -12562 426 -11574 457
rect -10932 491 -9944 1985
rect -9254 2127 -8266 3621
rect -7556 3763 -6568 5257
rect -5926 5399 -4938 6893
rect -4250 7037 -3262 8531
rect -2598 8673 -1610 10167
rect -968 10309 20 11803
rect 754 11945 1742 13439
rect 2360 13691 3348 15185
rect 4060 15327 5048 16821
rect 5736 16855 6724 17116
rect 5736 16821 5788 16855
rect 6572 16821 6724 16855
rect 4060 15293 4130 15327
rect 4914 15293 5048 15327
rect 4060 15219 5048 15293
rect 4060 15185 4130 15219
rect 4914 15185 5048 15219
rect 2360 13657 2472 13691
rect 3256 13657 3348 13691
rect 2360 13473 3348 13657
rect 2360 13439 2474 13473
rect 3258 13439 3348 13473
rect 754 11911 816 11945
rect 1600 11911 1742 11945
rect 754 11837 1742 11911
rect 754 11803 816 11837
rect 1600 11803 1742 11837
rect -968 10275 -842 10309
rect -58 10275 20 10309
rect -968 10201 20 10275
rect -968 10167 -842 10201
rect -58 10167 20 10201
rect -2598 8639 -2500 8673
rect -1716 8639 -1610 8673
rect -2598 8565 -1610 8639
rect -2598 8531 -2500 8565
rect -1716 8531 -1610 8565
rect -4250 7003 -4158 7037
rect -3374 7003 -3262 7037
rect -4250 6927 -3262 7003
rect -4250 6893 -4158 6927
rect -3374 6893 -3262 6927
rect -5926 5365 -5816 5399
rect -5032 5365 -4938 5399
rect -5926 5291 -4938 5365
rect -5926 5257 -5816 5291
rect -5032 5257 -4938 5291
rect -7556 3729 -7474 3763
rect -6690 3729 -6568 3763
rect -7556 3655 -6568 3729
rect -7556 3621 -7474 3655
rect -6690 3621 -6568 3655
rect -9254 2093 -9132 2127
rect -8348 2093 -8266 2127
rect -9254 2019 -8266 2093
rect -9254 1985 -9132 2019
rect -8348 1985 -8266 2019
rect -10932 457 -10790 491
rect -10006 457 -9944 491
rect -10932 426 -9944 457
rect -9254 491 -8266 1985
rect -7556 2127 -6568 3621
rect -5926 3763 -4938 5257
rect -4250 5399 -3262 6893
rect -2598 7037 -1610 8531
rect -968 8673 20 10167
rect 754 10309 1742 11803
rect 2360 11945 3348 13439
rect 4060 13691 5048 15185
rect 5736 15327 6724 16821
rect 7366 16855 8354 17092
rect 7366 16821 7446 16855
rect 8230 16821 8354 16855
rect 5736 15293 5788 15327
rect 6572 15293 6724 15327
rect 5736 15219 6724 15293
rect 5736 15185 5788 15219
rect 6572 15185 6724 15219
rect 4060 13657 4130 13691
rect 4914 13657 5048 13691
rect 4060 13473 5048 13657
rect 4060 13439 4132 13473
rect 4916 13439 5048 13473
rect 2360 11911 2474 11945
rect 3258 11911 3348 11945
rect 2360 11837 3348 11911
rect 2360 11803 2474 11837
rect 3258 11803 3348 11837
rect 754 10275 816 10309
rect 1600 10275 1742 10309
rect 754 10201 1742 10275
rect 754 10167 816 10201
rect 1600 10167 1742 10201
rect -968 8639 -842 8673
rect -58 8639 20 8673
rect -968 8565 20 8639
rect -968 8531 -842 8565
rect -58 8531 20 8565
rect -2598 7003 -2500 7037
rect -1716 7003 -1610 7037
rect -2598 6927 -1610 7003
rect -2598 6893 -2500 6927
rect -1716 6893 -1610 6927
rect -4250 5365 -4158 5399
rect -3374 5365 -3262 5399
rect -4250 5291 -3262 5365
rect -4250 5257 -4158 5291
rect -3374 5257 -3262 5291
rect -5926 3729 -5816 3763
rect -5032 3729 -4938 3763
rect -5926 3655 -4938 3729
rect -5926 3621 -5816 3655
rect -5032 3621 -4938 3655
rect -7556 2093 -7474 2127
rect -6690 2093 -6568 2127
rect -7556 2019 -6568 2093
rect -7556 1985 -7474 2019
rect -6690 1985 -6568 2019
rect -9254 457 -9132 491
rect -8348 457 -8266 491
rect -9254 426 -8266 457
rect -7556 491 -6568 1985
rect -5926 2127 -4938 3621
rect -4250 3763 -3262 5257
rect -2598 5399 -1610 6893
rect -968 7037 20 8531
rect 754 8673 1742 10167
rect 2360 10309 3348 11803
rect 4060 11945 5048 13439
rect 5736 13691 6724 15185
rect 7366 15327 8354 16821
rect 8994 16855 9982 17116
rect 8994 16821 9104 16855
rect 9888 16821 9982 16855
rect 7366 15293 7446 15327
rect 8230 15293 8354 15327
rect 7366 15219 8354 15293
rect 7366 15185 7446 15219
rect 8230 15185 8354 15219
rect 5736 13657 5788 13691
rect 6572 13657 6724 13691
rect 5736 13473 6724 13657
rect 5736 13439 5790 13473
rect 6574 13439 6724 13473
rect 4060 11911 4132 11945
rect 4916 11911 5048 11945
rect 4060 11837 5048 11911
rect 4060 11803 4132 11837
rect 4916 11803 5048 11837
rect 2360 10275 2474 10309
rect 3258 10275 3348 10309
rect 2360 10201 3348 10275
rect 2360 10167 2474 10201
rect 3258 10167 3348 10201
rect 754 8639 816 8673
rect 1600 8639 1742 8673
rect 754 8565 1742 8639
rect 754 8531 816 8565
rect 1600 8531 1742 8565
rect -968 7003 -842 7037
rect -58 7003 20 7037
rect -968 6927 20 7003
rect -968 6893 -842 6927
rect -58 6893 20 6927
rect -2598 5365 -2500 5399
rect -1716 5365 -1610 5399
rect -2598 5291 -1610 5365
rect -2598 5257 -2500 5291
rect -1716 5257 -1610 5291
rect -4250 3729 -4158 3763
rect -3374 3729 -3262 3763
rect -4250 3655 -3262 3729
rect -4250 3621 -4158 3655
rect -3374 3621 -3262 3655
rect -5926 2093 -5816 2127
rect -5032 2093 -4938 2127
rect -5926 2019 -4938 2093
rect -5926 1985 -5816 2019
rect -5032 1985 -4938 2019
rect -7556 457 -7474 491
rect -6690 457 -6568 491
rect -7556 426 -6568 457
rect -5926 491 -4938 1985
rect -4250 2127 -3262 3621
rect -2598 3763 -1610 5257
rect -968 5399 20 6893
rect 754 7037 1742 8531
rect 2360 8673 3348 10167
rect 4060 10309 5048 11803
rect 5736 11945 6724 13439
rect 7366 13691 8354 15185
rect 8994 15327 9982 16821
rect 10678 16855 11666 17070
rect 10678 16821 10762 16855
rect 11546 16821 11666 16855
rect 8994 15293 9104 15327
rect 9888 15293 9982 15327
rect 8994 15219 9982 15293
rect 8994 15185 9104 15219
rect 9888 15185 9982 15219
rect 7366 13657 7446 13691
rect 8230 13657 8354 13691
rect 7366 13473 8354 13657
rect 7366 13439 7448 13473
rect 8232 13439 8354 13473
rect 5736 11911 5790 11945
rect 6574 11911 6724 11945
rect 5736 11837 6724 11911
rect 5736 11803 5790 11837
rect 6574 11803 6724 11837
rect 4060 10275 4132 10309
rect 4916 10275 5048 10309
rect 4060 10201 5048 10275
rect 4060 10167 4132 10201
rect 4916 10167 5048 10201
rect 2360 8639 2474 8673
rect 3258 8639 3348 8673
rect 2360 8565 3348 8639
rect 2360 8531 2474 8565
rect 3258 8531 3348 8565
rect 754 7003 816 7037
rect 1600 7003 1742 7037
rect 754 6927 1742 7003
rect 754 6893 816 6927
rect 1600 6893 1742 6927
rect -968 5365 -842 5399
rect -58 5365 20 5399
rect -968 5291 20 5365
rect -968 5257 -842 5291
rect -58 5257 20 5291
rect -2598 3729 -2500 3763
rect -1716 3729 -1610 3763
rect -2598 3655 -1610 3729
rect -2598 3621 -2500 3655
rect -1716 3621 -1610 3655
rect -4250 2093 -4158 2127
rect -3374 2093 -3262 2127
rect -4250 2019 -3262 2093
rect -4250 1985 -4158 2019
rect -3374 1985 -3262 2019
rect -5926 457 -5816 491
rect -5032 457 -4938 491
rect -5926 426 -4938 457
rect -4250 491 -3262 1985
rect -2598 2127 -1610 3621
rect -968 3763 20 5257
rect 754 5399 1742 6893
rect 2360 7037 3348 8531
rect 4060 8673 5048 10167
rect 5736 10309 6724 11803
rect 7366 11945 8354 13439
rect 8994 13691 9982 15185
rect 10678 15327 11666 16821
rect 12352 16855 13340 17086
rect 12352 16821 12420 16855
rect 13204 16821 13340 16855
rect 10678 15293 10762 15327
rect 11546 15293 11666 15327
rect 10678 15219 11666 15293
rect 10678 15185 10762 15219
rect 11546 15185 11666 15219
rect 8994 13657 9104 13691
rect 9888 13657 9982 13691
rect 8994 13473 9982 13657
rect 8994 13439 9106 13473
rect 9890 13439 9982 13473
rect 7366 11911 7448 11945
rect 8232 11911 8354 11945
rect 7366 11837 8354 11911
rect 7366 11803 7448 11837
rect 8232 11803 8354 11837
rect 5736 10275 5790 10309
rect 6574 10275 6724 10309
rect 5736 10201 6724 10275
rect 5736 10167 5790 10201
rect 6574 10167 6724 10201
rect 4060 8639 4132 8673
rect 4916 8639 5048 8673
rect 4060 8565 5048 8639
rect 4060 8531 4132 8565
rect 4916 8531 5048 8565
rect 2360 7003 2474 7037
rect 3258 7003 3348 7037
rect 2360 6927 3348 7003
rect 2360 6893 2474 6927
rect 3258 6893 3348 6927
rect 754 5365 816 5399
rect 1600 5365 1742 5399
rect 754 5291 1742 5365
rect 754 5257 816 5291
rect 1600 5257 1742 5291
rect -968 3729 -842 3763
rect -58 3729 20 3763
rect -968 3655 20 3729
rect -968 3621 -842 3655
rect -58 3621 20 3655
rect -2598 2093 -2500 2127
rect -1716 2093 -1610 2127
rect -2598 2019 -1610 2093
rect -2598 1985 -2500 2019
rect -1716 1985 -1610 2019
rect -4250 457 -4158 491
rect -3374 457 -3262 491
rect -4250 426 -3262 457
rect -2598 491 -1610 1985
rect -968 2127 20 3621
rect 754 3763 1742 5257
rect 2360 5399 3348 6893
rect 4060 7037 5048 8531
rect 5736 8673 6724 10167
rect 7366 10309 8354 11803
rect 8994 11945 9982 13439
rect 10678 13691 11666 15185
rect 12352 15327 13340 16821
rect 14002 16855 14990 17110
rect 14002 16821 14078 16855
rect 14862 16821 14990 16855
rect 12352 15293 12420 15327
rect 13204 15293 13340 15327
rect 12352 15219 13340 15293
rect 12352 15185 12420 15219
rect 13204 15185 13340 15219
rect 10678 13657 10762 13691
rect 11546 13657 11666 13691
rect 10678 13473 11666 13657
rect 10678 13439 10764 13473
rect 11548 13439 11666 13473
rect 8994 11911 9106 11945
rect 9890 11911 9982 11945
rect 8994 11837 9982 11911
rect 8994 11803 9106 11837
rect 9890 11803 9982 11837
rect 7366 10275 7448 10309
rect 8232 10275 8354 10309
rect 7366 10201 8354 10275
rect 7366 10167 7448 10201
rect 8232 10167 8354 10201
rect 5736 8639 5790 8673
rect 6574 8639 6724 8673
rect 5736 8565 6724 8639
rect 5736 8531 5790 8565
rect 6574 8531 6724 8565
rect 4060 7003 4132 7037
rect 4916 7003 5048 7037
rect 4060 6927 5048 7003
rect 4060 6893 4132 6927
rect 4916 6893 5048 6927
rect 2360 5365 2474 5399
rect 3258 5365 3348 5399
rect 2360 5291 3348 5365
rect 2360 5257 2474 5291
rect 3258 5257 3348 5291
rect 754 3729 816 3763
rect 1600 3729 1742 3763
rect 754 3655 1742 3729
rect 754 3621 816 3655
rect 1600 3621 1742 3655
rect -968 2093 -842 2127
rect -58 2093 20 2127
rect -968 2019 20 2093
rect -968 1985 -842 2019
rect -58 1985 20 2019
rect -2598 457 -2500 491
rect -1716 457 -1610 491
rect -2598 426 -1610 457
rect -968 491 20 1985
rect 754 2127 1742 3621
rect 2360 3763 3348 5257
rect 4060 5399 5048 6893
rect 5736 7037 6724 8531
rect 7366 8673 8354 10167
rect 8994 10309 9982 11803
rect 10678 11945 11666 13439
rect 12352 13691 13340 15185
rect 14002 15327 14990 16821
rect 15608 16855 16596 17086
rect 15608 16821 15736 16855
rect 16520 16821 16596 16855
rect 14002 15293 14078 15327
rect 14862 15293 14990 15327
rect 14002 15219 14990 15293
rect 14002 15185 14078 15219
rect 14862 15185 14990 15219
rect 12352 13657 12420 13691
rect 13204 13657 13340 13691
rect 12352 13473 13340 13657
rect 12352 13439 12422 13473
rect 13206 13439 13340 13473
rect 10678 11911 10764 11945
rect 11548 11911 11666 11945
rect 10678 11837 11666 11911
rect 10678 11803 10764 11837
rect 11548 11803 11666 11837
rect 8994 10275 9106 10309
rect 9890 10275 9982 10309
rect 8994 10201 9982 10275
rect 8994 10167 9106 10201
rect 9890 10167 9982 10201
rect 7366 8639 7448 8673
rect 8232 8639 8354 8673
rect 7366 8565 8354 8639
rect 7366 8531 7448 8565
rect 8232 8531 8354 8565
rect 5736 7003 5790 7037
rect 6574 7003 6724 7037
rect 5736 6927 6724 7003
rect 5736 6893 5790 6927
rect 6574 6893 6724 6927
rect 4060 5365 4132 5399
rect 4916 5365 5048 5399
rect 4060 5291 5048 5365
rect 4060 5257 4132 5291
rect 4916 5257 5048 5291
rect 2360 3729 2474 3763
rect 3258 3729 3348 3763
rect 2360 3655 3348 3729
rect 2360 3621 2474 3655
rect 3258 3621 3348 3655
rect 754 2093 816 2127
rect 1600 2093 1742 2127
rect 754 2019 1742 2093
rect 754 1985 816 2019
rect 1600 1985 1742 2019
rect 754 512 1742 1985
rect 2360 2127 3348 3621
rect 4060 3763 5048 5257
rect 5736 5399 6724 6893
rect 7366 7037 8354 8531
rect 8994 8673 9982 10167
rect 10678 10309 11666 11803
rect 12352 11945 13340 13439
rect 14002 13691 14990 15185
rect 15608 15327 16596 16821
rect 17306 16855 18294 17110
rect 17306 16821 17394 16855
rect 18178 16821 18294 16855
rect 15608 15293 15736 15327
rect 16520 15293 16596 15327
rect 15608 15219 16596 15293
rect 15608 15185 15736 15219
rect 16520 15185 16596 15219
rect 14002 13657 14078 13691
rect 14862 13657 14990 13691
rect 14002 13473 14990 13657
rect 14002 13439 14080 13473
rect 14864 13439 14990 13473
rect 12352 11911 12422 11945
rect 13206 11911 13340 11945
rect 12352 11837 13340 11911
rect 12352 11803 12422 11837
rect 13206 11803 13340 11837
rect 10678 10275 10764 10309
rect 11548 10275 11666 10309
rect 10678 10201 11666 10275
rect 10678 10167 10764 10201
rect 11548 10167 11666 10201
rect 8994 8639 9106 8673
rect 9890 8639 9982 8673
rect 8994 8565 9982 8639
rect 8994 8531 9106 8565
rect 9890 8531 9982 8565
rect 7366 7003 7448 7037
rect 8232 7003 8354 7037
rect 7366 6927 8354 7003
rect 7366 6893 7448 6927
rect 8232 6893 8354 6927
rect 5736 5365 5790 5399
rect 6574 5365 6724 5399
rect 5736 5291 6724 5365
rect 5736 5257 5790 5291
rect 6574 5257 6724 5291
rect 4060 3729 4132 3763
rect 4916 3729 5048 3763
rect 4060 3655 5048 3729
rect 4060 3621 4132 3655
rect 4916 3621 5048 3655
rect 2360 2093 2474 2127
rect 3258 2093 3348 2127
rect 2360 2019 3348 2093
rect 2360 1985 2474 2019
rect 3258 1985 3348 2019
rect -968 457 -842 491
rect -58 457 20 491
rect -968 426 20 457
rect -32422 388 20 426
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -732 292 20 388
rect 760 491 1742 512
rect 760 470 816 491
rect 760 436 802 470
rect 1600 457 1742 491
rect 836 442 1742 457
rect 2360 491 3348 1985
rect 4060 2127 5048 3621
rect 5736 3763 6724 5257
rect 7366 5399 8354 6893
rect 8994 7037 9982 8531
rect 10678 8673 11666 10167
rect 12352 10309 13340 11803
rect 14002 11945 14990 13439
rect 15608 13691 16596 15185
rect 17306 15327 18294 16821
rect 18958 16855 19946 17086
rect 18958 16821 19052 16855
rect 19836 16821 19946 16855
rect 17306 15293 17394 15327
rect 18178 15293 18294 15327
rect 17306 15219 18294 15293
rect 17306 15185 17394 15219
rect 18178 15185 18294 15219
rect 15608 13657 15736 13691
rect 16520 13657 16596 13691
rect 15608 13473 16596 13657
rect 15608 13439 15738 13473
rect 16522 13439 16596 13473
rect 14002 11911 14080 11945
rect 14864 11911 14990 11945
rect 14002 11837 14990 11911
rect 14002 11803 14080 11837
rect 14864 11803 14990 11837
rect 12352 10275 12422 10309
rect 13206 10275 13340 10309
rect 12352 10201 13340 10275
rect 12352 10167 12422 10201
rect 13206 10167 13340 10201
rect 10678 8639 10764 8673
rect 11548 8639 11666 8673
rect 10678 8565 11666 8639
rect 10678 8531 10764 8565
rect 11548 8531 11666 8565
rect 8994 7003 9106 7037
rect 9890 7003 9982 7037
rect 8994 6927 9982 7003
rect 8994 6893 9106 6927
rect 9890 6893 9982 6927
rect 7366 5365 7448 5399
rect 8232 5365 8354 5399
rect 7366 5291 8354 5365
rect 7366 5257 7448 5291
rect 8232 5257 8354 5291
rect 5736 3729 5790 3763
rect 6574 3729 6724 3763
rect 5736 3655 6724 3729
rect 5736 3621 5790 3655
rect 6574 3621 6724 3655
rect 4060 2093 4132 2127
rect 4916 2093 5048 2127
rect 4060 2019 5048 2093
rect 4060 1985 4132 2019
rect 4916 1985 5048 2019
rect 2360 457 2474 491
rect 3258 457 3348 491
rect 2360 442 3348 457
rect 4060 491 5048 1985
rect 5736 2127 6724 3621
rect 7366 3763 8354 5257
rect 8994 5399 9982 6893
rect 10678 7037 11666 8531
rect 12352 8673 13340 10167
rect 14002 10309 14990 11803
rect 15608 11945 16596 13439
rect 17306 13691 18294 15185
rect 18958 15327 19946 16821
rect 20608 16855 21596 17110
rect 20608 16821 20710 16855
rect 21494 16821 21596 16855
rect 18958 15293 19052 15327
rect 19836 15293 19946 15327
rect 18958 15219 19946 15293
rect 18958 15185 19052 15219
rect 19836 15185 19946 15219
rect 17306 13657 17394 13691
rect 18178 13657 18294 13691
rect 17306 13473 18294 13657
rect 17306 13439 17396 13473
rect 18180 13439 18294 13473
rect 15608 11911 15738 11945
rect 16522 11911 16596 11945
rect 15608 11837 16596 11911
rect 15608 11803 15738 11837
rect 16522 11803 16596 11837
rect 14002 10275 14080 10309
rect 14864 10275 14990 10309
rect 14002 10201 14990 10275
rect 14002 10167 14080 10201
rect 14864 10167 14990 10201
rect 12352 8639 12422 8673
rect 13206 8639 13340 8673
rect 12352 8565 13340 8639
rect 12352 8531 12422 8565
rect 13206 8531 13340 8565
rect 10678 7003 10764 7037
rect 11548 7003 11666 7037
rect 10678 6927 11666 7003
rect 10678 6893 10764 6927
rect 11548 6893 11666 6927
rect 8994 5365 9106 5399
rect 9890 5365 9982 5399
rect 8994 5291 9982 5365
rect 8994 5257 9106 5291
rect 9890 5257 9982 5291
rect 7366 3729 7448 3763
rect 8232 3729 8354 3763
rect 7366 3655 8354 3729
rect 7366 3621 7448 3655
rect 8232 3621 8354 3655
rect 5736 2093 5790 2127
rect 6574 2093 6724 2127
rect 5736 2019 6724 2093
rect 5736 1985 5790 2019
rect 6574 1985 6724 2019
rect 4060 457 4132 491
rect 4916 457 5048 491
rect 4060 442 5048 457
rect 5736 491 6724 1985
rect 7366 2127 8354 3621
rect 8994 3763 9982 5257
rect 10678 5399 11666 6893
rect 12352 7037 13340 8531
rect 14002 8673 14990 10167
rect 15608 10309 16596 11803
rect 17306 11945 18294 13439
rect 18958 13691 19946 15185
rect 20608 15327 21596 16821
rect 22260 16855 23248 17086
rect 22260 16821 22368 16855
rect 23152 16821 23248 16855
rect 20608 15293 20710 15327
rect 21494 15293 21596 15327
rect 20608 15219 21596 15293
rect 20608 15185 20710 15219
rect 21494 15185 21596 15219
rect 18958 13657 19052 13691
rect 19836 13657 19946 13691
rect 18958 13473 19946 13657
rect 18958 13439 19054 13473
rect 19838 13439 19946 13473
rect 17306 11911 17396 11945
rect 18180 11911 18294 11945
rect 17306 11837 18294 11911
rect 17306 11803 17396 11837
rect 18180 11803 18294 11837
rect 15608 10275 15738 10309
rect 16522 10275 16596 10309
rect 15608 10201 16596 10275
rect 15608 10167 15738 10201
rect 16522 10167 16596 10201
rect 14002 8639 14080 8673
rect 14864 8639 14990 8673
rect 14002 8565 14990 8639
rect 14002 8531 14080 8565
rect 14864 8531 14990 8565
rect 12352 7003 12422 7037
rect 13206 7003 13340 7037
rect 12352 6927 13340 7003
rect 12352 6893 12422 6927
rect 13206 6893 13340 6927
rect 10678 5365 10764 5399
rect 11548 5365 11666 5399
rect 10678 5291 11666 5365
rect 10678 5257 10764 5291
rect 11548 5257 11666 5291
rect 8994 3729 9106 3763
rect 9890 3729 9982 3763
rect 8994 3655 9982 3729
rect 8994 3621 9106 3655
rect 9890 3621 9982 3655
rect 7366 2093 7448 2127
rect 8232 2093 8354 2127
rect 7366 2019 8354 2093
rect 7366 1985 7448 2019
rect 8232 1985 8354 2019
rect 5736 457 5790 491
rect 6574 457 6724 491
rect 5736 442 6724 457
rect 7366 491 8354 1985
rect 8994 2127 9982 3621
rect 10678 3763 11666 5257
rect 12352 5399 13340 6893
rect 14002 7037 14990 8531
rect 15608 8673 16596 10167
rect 17306 10309 18294 11803
rect 18958 11945 19946 13439
rect 20608 13691 21596 15185
rect 22260 15327 23248 16821
rect 23918 16855 24906 17088
rect 23918 16821 24026 16855
rect 24810 16821 24906 16855
rect 22260 15293 22368 15327
rect 23152 15293 23248 15327
rect 22260 15219 23248 15293
rect 22260 15185 22368 15219
rect 23152 15185 23248 15219
rect 20608 13657 20710 13691
rect 21494 13657 21596 13691
rect 20608 13473 21596 13657
rect 20608 13439 20712 13473
rect 21496 13439 21596 13473
rect 18958 11911 19054 11945
rect 19838 11911 19946 11945
rect 18958 11837 19946 11911
rect 18958 11803 19054 11837
rect 19838 11803 19946 11837
rect 17306 10275 17396 10309
rect 18180 10275 18294 10309
rect 17306 10201 18294 10275
rect 17306 10167 17396 10201
rect 18180 10167 18294 10201
rect 15608 8639 15738 8673
rect 16522 8639 16596 8673
rect 15608 8565 16596 8639
rect 15608 8531 15738 8565
rect 16522 8531 16596 8565
rect 14002 7003 14080 7037
rect 14864 7003 14990 7037
rect 14002 6927 14990 7003
rect 14002 6893 14080 6927
rect 14864 6893 14990 6927
rect 12352 5365 12422 5399
rect 13206 5365 13340 5399
rect 12352 5291 13340 5365
rect 12352 5257 12422 5291
rect 13206 5257 13340 5291
rect 10678 3729 10764 3763
rect 11548 3729 11666 3763
rect 10678 3655 11666 3729
rect 10678 3621 10764 3655
rect 11548 3621 11666 3655
rect 8994 2093 9106 2127
rect 9890 2093 9982 2127
rect 8994 2019 9982 2093
rect 8994 1985 9106 2019
rect 9890 1985 9982 2019
rect 7366 457 7448 491
rect 8232 457 8354 491
rect 7366 442 8354 457
rect 8994 491 9982 1985
rect 10678 2127 11666 3621
rect 12352 3763 13340 5257
rect 14002 5399 14990 6893
rect 15608 7037 16596 8531
rect 17306 8673 18294 10167
rect 18958 10309 19946 11803
rect 20608 11945 21596 13439
rect 22260 13691 23248 15185
rect 23918 15327 24906 16821
rect 25566 16855 26554 17088
rect 25566 16821 25684 16855
rect 26468 16821 26554 16855
rect 23918 15293 24026 15327
rect 24810 15293 24906 15327
rect 23918 15219 24906 15293
rect 23918 15185 24026 15219
rect 24810 15185 24906 15219
rect 22260 13657 22368 13691
rect 23152 13657 23248 13691
rect 22260 13473 23248 13657
rect 22260 13439 22370 13473
rect 23154 13439 23248 13473
rect 20608 11911 20712 11945
rect 21496 11911 21596 11945
rect 20608 11837 21596 11911
rect 20608 11803 20712 11837
rect 21496 11803 21596 11837
rect 18958 10275 19054 10309
rect 19838 10275 19946 10309
rect 18958 10201 19946 10275
rect 18958 10167 19054 10201
rect 19838 10167 19946 10201
rect 17306 8639 17396 8673
rect 18180 8639 18294 8673
rect 17306 8565 18294 8639
rect 17306 8531 17396 8565
rect 18180 8531 18294 8565
rect 15608 7003 15738 7037
rect 16522 7003 16596 7037
rect 15608 6927 16596 7003
rect 15608 6893 15738 6927
rect 16522 6893 16596 6927
rect 14002 5365 14080 5399
rect 14864 5365 14990 5399
rect 14002 5291 14990 5365
rect 14002 5257 14080 5291
rect 14864 5257 14990 5291
rect 12352 3729 12422 3763
rect 13206 3729 13340 3763
rect 12352 3655 13340 3729
rect 12352 3621 12422 3655
rect 13206 3621 13340 3655
rect 10678 2093 10764 2127
rect 11548 2093 11666 2127
rect 10678 2019 11666 2093
rect 10678 1985 10764 2019
rect 11548 1985 11666 2019
rect 8994 457 9106 491
rect 9890 457 9982 491
rect 8994 442 9982 457
rect 10678 491 11666 1985
rect 12352 2127 13340 3621
rect 14002 3763 14990 5257
rect 15608 5399 16596 6893
rect 17306 7037 18294 8531
rect 18958 8673 19946 10167
rect 20608 10309 21596 11803
rect 22260 11945 23248 13439
rect 23918 13691 24906 15185
rect 25566 15327 26554 16821
rect 27260 16855 28248 17088
rect 27260 16821 27342 16855
rect 28126 16821 28248 16855
rect 25566 15293 25684 15327
rect 26468 15293 26554 15327
rect 25566 15219 26554 15293
rect 25566 15185 25684 15219
rect 26468 15185 26554 15219
rect 23918 13657 24026 13691
rect 24810 13657 24906 13691
rect 23918 13473 24906 13657
rect 23918 13439 24028 13473
rect 24812 13439 24906 13473
rect 22260 11911 22370 11945
rect 23154 11911 23248 11945
rect 22260 11837 23248 11911
rect 22260 11803 22370 11837
rect 23154 11803 23248 11837
rect 20608 10275 20712 10309
rect 21496 10275 21596 10309
rect 20608 10201 21596 10275
rect 20608 10167 20712 10201
rect 21496 10167 21596 10201
rect 18958 8639 19054 8673
rect 19838 8639 19946 8673
rect 18958 8565 19946 8639
rect 18958 8531 19054 8565
rect 19838 8531 19946 8565
rect 17306 7003 17396 7037
rect 18180 7003 18294 7037
rect 17306 6927 18294 7003
rect 17306 6893 17396 6927
rect 18180 6893 18294 6927
rect 15608 5365 15738 5399
rect 16522 5365 16596 5399
rect 15608 5291 16596 5365
rect 15608 5257 15738 5291
rect 16522 5257 16596 5291
rect 14002 3729 14080 3763
rect 14864 3729 14990 3763
rect 14002 3655 14990 3729
rect 14002 3621 14080 3655
rect 14864 3621 14990 3655
rect 12352 2093 12422 2127
rect 13206 2093 13340 2127
rect 12352 2019 13340 2093
rect 12352 1985 12422 2019
rect 13206 1985 13340 2019
rect 10678 457 10764 491
rect 11548 457 11666 491
rect 10678 442 11666 457
rect 12352 491 13340 1985
rect 14002 2127 14990 3621
rect 15608 3763 16596 5257
rect 17306 5399 18294 6893
rect 18958 7037 19946 8531
rect 20608 8673 21596 10167
rect 22260 10309 23248 11803
rect 23918 11945 24906 13439
rect 25566 13691 26554 15185
rect 27260 15327 28248 16821
rect 28908 16855 29896 17136
rect 28908 16821 29000 16855
rect 29784 16821 29896 16855
rect 27260 15293 27342 15327
rect 28126 15293 28248 15327
rect 27260 15219 28248 15293
rect 27260 15185 27342 15219
rect 28126 15185 28248 15219
rect 25566 13657 25684 13691
rect 26468 13657 26554 13691
rect 25566 13473 26554 13657
rect 25566 13439 25686 13473
rect 26470 13439 26554 13473
rect 23918 11911 24028 11945
rect 24812 11911 24906 11945
rect 23918 11837 24906 11911
rect 23918 11803 24028 11837
rect 24812 11803 24906 11837
rect 22260 10275 22370 10309
rect 23154 10275 23248 10309
rect 22260 10201 23248 10275
rect 22260 10167 22370 10201
rect 23154 10167 23248 10201
rect 20608 8639 20712 8673
rect 21496 8639 21596 8673
rect 20608 8565 21596 8639
rect 20608 8531 20712 8565
rect 21496 8531 21596 8565
rect 18958 7003 19054 7037
rect 19838 7003 19946 7037
rect 18958 6927 19946 7003
rect 18958 6893 19054 6927
rect 19838 6893 19946 6927
rect 17306 5365 17396 5399
rect 18180 5365 18294 5399
rect 17306 5291 18294 5365
rect 17306 5257 17396 5291
rect 18180 5257 18294 5291
rect 15608 3729 15738 3763
rect 16522 3729 16596 3763
rect 15608 3655 16596 3729
rect 15608 3621 15738 3655
rect 16522 3621 16596 3655
rect 14002 2093 14080 2127
rect 14864 2093 14990 2127
rect 14002 2019 14990 2093
rect 14002 1985 14080 2019
rect 14864 1985 14990 2019
rect 12352 457 12422 491
rect 13206 457 13340 491
rect 12352 442 13340 457
rect 14002 491 14990 1985
rect 15608 2127 16596 3621
rect 17306 3763 18294 5257
rect 18958 5399 19946 6893
rect 20608 7037 21596 8531
rect 22260 8673 23248 10167
rect 23918 10309 24906 11803
rect 25566 11945 26554 13439
rect 27260 13691 28248 15185
rect 28908 15327 29896 16821
rect 30556 16855 31544 17112
rect 30556 16821 30658 16855
rect 31442 16821 31544 16855
rect 28908 15293 29000 15327
rect 29784 15293 29896 15327
rect 28908 15219 29896 15293
rect 28908 15185 29000 15219
rect 29784 15185 29896 15219
rect 27260 13657 27342 13691
rect 28126 13657 28248 13691
rect 27260 13473 28248 13657
rect 27260 13439 27344 13473
rect 28128 13439 28248 13473
rect 25566 11911 25686 11945
rect 26470 11911 26554 11945
rect 25566 11837 26554 11911
rect 25566 11803 25686 11837
rect 26470 11803 26554 11837
rect 23918 10275 24028 10309
rect 24812 10275 24906 10309
rect 23918 10201 24906 10275
rect 23918 10167 24028 10201
rect 24812 10167 24906 10201
rect 22260 8639 22370 8673
rect 23154 8639 23248 8673
rect 22260 8565 23248 8639
rect 22260 8531 22370 8565
rect 23154 8531 23248 8565
rect 20608 7003 20712 7037
rect 21496 7003 21596 7037
rect 20608 6927 21596 7003
rect 20608 6893 20712 6927
rect 21496 6893 21596 6927
rect 18958 5365 19054 5399
rect 19838 5365 19946 5399
rect 18958 5291 19946 5365
rect 18958 5257 19054 5291
rect 19838 5257 19946 5291
rect 17306 3729 17396 3763
rect 18180 3729 18294 3763
rect 17306 3655 18294 3729
rect 17306 3621 17396 3655
rect 18180 3621 18294 3655
rect 15608 2093 15738 2127
rect 16522 2093 16596 2127
rect 15608 2019 16596 2093
rect 15608 1985 15738 2019
rect 16522 1985 16596 2019
rect 14002 457 14080 491
rect 14864 457 14990 491
rect 14002 442 14990 457
rect 15608 491 16596 1985
rect 17306 2127 18294 3621
rect 18958 3763 19946 5257
rect 20608 5399 21596 6893
rect 22260 7037 23248 8531
rect 23918 8673 24906 10167
rect 25566 10309 26554 11803
rect 27260 11945 28248 13439
rect 28908 13691 29896 15185
rect 30556 15327 31544 16821
rect 32204 16855 33192 17064
rect 32204 16821 32316 16855
rect 33100 16821 33192 16855
rect 30556 15293 30658 15327
rect 31442 15293 31544 15327
rect 30556 15219 31544 15293
rect 30556 15185 30658 15219
rect 31442 15185 31544 15219
rect 28908 13657 29000 13691
rect 29784 13657 29896 13691
rect 28908 13473 29896 13657
rect 28908 13439 29002 13473
rect 29786 13439 29896 13473
rect 27260 11911 27344 11945
rect 28128 11911 28248 11945
rect 27260 11837 28248 11911
rect 27260 11803 27344 11837
rect 28128 11803 28248 11837
rect 25566 10275 25686 10309
rect 26470 10275 26554 10309
rect 25566 10201 26554 10275
rect 25566 10167 25686 10201
rect 26470 10167 26554 10201
rect 23918 8639 24028 8673
rect 24812 8639 24906 8673
rect 23918 8565 24906 8639
rect 23918 8531 24028 8565
rect 24812 8531 24906 8565
rect 22260 7003 22370 7037
rect 23154 7003 23248 7037
rect 22260 6927 23248 7003
rect 22260 6893 22370 6927
rect 23154 6893 23248 6927
rect 20608 5365 20712 5399
rect 21496 5365 21596 5399
rect 20608 5291 21596 5365
rect 20608 5257 20712 5291
rect 21496 5257 21596 5291
rect 18958 3729 19054 3763
rect 19838 3729 19946 3763
rect 18958 3655 19946 3729
rect 18958 3621 19054 3655
rect 19838 3621 19946 3655
rect 17306 2093 17396 2127
rect 18180 2093 18294 2127
rect 17306 2019 18294 2093
rect 17306 1985 17396 2019
rect 18180 1985 18294 2019
rect 15608 457 15738 491
rect 16522 457 16596 491
rect 15608 442 16596 457
rect 17306 491 18294 1985
rect 18958 2127 19946 3621
rect 20608 3763 21596 5257
rect 22260 5399 23248 6893
rect 23918 7037 24906 8531
rect 25566 8673 26554 10167
rect 27260 10309 28248 11803
rect 28908 11945 29896 13439
rect 30556 13691 31544 15185
rect 32204 15327 33192 16821
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 32204 15293 32316 15327
rect 33100 15293 33192 15327
rect 32204 15219 33192 15293
rect 32204 15185 32316 15219
rect 33100 15185 33192 15219
rect 30556 13657 30658 13691
rect 31442 13657 31544 13691
rect 30556 13473 31544 13657
rect 30556 13439 30660 13473
rect 31444 13439 31544 13473
rect 28908 11911 29002 11945
rect 29786 11911 29896 11945
rect 28908 11837 29896 11911
rect 28908 11803 29002 11837
rect 29786 11803 29896 11837
rect 27260 10275 27344 10309
rect 28128 10275 28248 10309
rect 27260 10201 28248 10275
rect 27260 10167 27344 10201
rect 28128 10167 28248 10201
rect 25566 8639 25686 8673
rect 26470 8639 26554 8673
rect 25566 8565 26554 8639
rect 25566 8531 25686 8565
rect 26470 8531 26554 8565
rect 23918 7003 24028 7037
rect 24812 7003 24906 7037
rect 23918 6927 24906 7003
rect 23918 6893 24028 6927
rect 24812 6893 24906 6927
rect 22260 5365 22370 5399
rect 23154 5365 23248 5399
rect 22260 5291 23248 5365
rect 22260 5257 22370 5291
rect 23154 5257 23248 5291
rect 20608 3729 20712 3763
rect 21496 3729 21596 3763
rect 20608 3655 21596 3729
rect 20608 3621 20712 3655
rect 21496 3621 21596 3655
rect 18958 2093 19054 2127
rect 19838 2093 19946 2127
rect 18958 2019 19946 2093
rect 18958 1985 19054 2019
rect 19838 1985 19946 2019
rect 17306 457 17396 491
rect 18180 457 18294 491
rect 17306 442 18294 457
rect 18958 491 19946 1985
rect 20608 2127 21596 3621
rect 22260 3763 23248 5257
rect 23918 5399 24906 6893
rect 25566 7037 26554 8531
rect 27260 8673 28248 10167
rect 28908 10309 29896 11803
rect 30556 11945 31544 13439
rect 32204 13691 33192 15185
rect 33976 13946 35004 15480
rect 32204 13657 32316 13691
rect 33100 13657 33192 13691
rect 32204 13473 33192 13657
rect 32204 13439 32318 13473
rect 33102 13439 33192 13473
rect 30556 11911 30660 11945
rect 31444 11911 31544 11945
rect 30556 11837 31544 11911
rect 30556 11803 30660 11837
rect 31444 11803 31544 11837
rect 28908 10275 29002 10309
rect 29786 10275 29896 10309
rect 28908 10201 29896 10275
rect 28908 10167 29002 10201
rect 29786 10167 29896 10201
rect 27260 8639 27344 8673
rect 28128 8639 28248 8673
rect 27260 8565 28248 8639
rect 27260 8531 27344 8565
rect 28128 8531 28248 8565
rect 25566 7003 25686 7037
rect 26470 7003 26554 7037
rect 25566 6927 26554 7003
rect 25566 6893 25686 6927
rect 26470 6893 26554 6927
rect 23918 5365 24028 5399
rect 24812 5365 24906 5399
rect 23918 5291 24906 5365
rect 23918 5257 24028 5291
rect 24812 5257 24906 5291
rect 22260 3729 22370 3763
rect 23154 3729 23248 3763
rect 22260 3655 23248 3729
rect 22260 3621 22370 3655
rect 23154 3621 23248 3655
rect 20608 2093 20712 2127
rect 21496 2093 21596 2127
rect 20608 2019 21596 2093
rect 20608 1985 20712 2019
rect 21496 1985 21596 2019
rect 18958 457 19054 491
rect 19838 457 19946 491
rect 18958 442 19946 457
rect 20608 491 21596 1985
rect 22260 2127 23248 3621
rect 23918 3763 24906 5257
rect 25566 5399 26554 6893
rect 27260 7037 28248 8531
rect 28908 8673 29896 10167
rect 30556 10309 31544 11803
rect 32204 11945 33192 13439
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 32204 11911 32318 11945
rect 33102 11911 33192 11945
rect 32204 11837 33192 11911
rect 32204 11803 32318 11837
rect 33102 11803 33192 11837
rect 30556 10275 30660 10309
rect 31444 10275 31544 10309
rect 30556 10201 31544 10275
rect 30556 10167 30660 10201
rect 31444 10167 31544 10201
rect 28908 8639 29002 8673
rect 29786 8639 29896 8673
rect 28908 8565 29896 8639
rect 28908 8531 29002 8565
rect 29786 8531 29896 8565
rect 27260 7003 27344 7037
rect 28128 7003 28248 7037
rect 27260 6927 28248 7003
rect 27260 6893 27344 6927
rect 28128 6893 28248 6927
rect 25566 5365 25686 5399
rect 26470 5365 26554 5399
rect 25566 5291 26554 5365
rect 25566 5257 25686 5291
rect 26470 5257 26554 5291
rect 23918 3729 24028 3763
rect 24812 3729 24906 3763
rect 23918 3655 24906 3729
rect 23918 3621 24028 3655
rect 24812 3621 24906 3655
rect 22260 2093 22370 2127
rect 23154 2093 23248 2127
rect 22260 2019 23248 2093
rect 22260 1985 22370 2019
rect 23154 1985 23248 2019
rect 20608 457 20712 491
rect 21496 457 21596 491
rect 20608 442 21596 457
rect 22260 491 23248 1985
rect 23918 2127 24906 3621
rect 25566 3763 26554 5257
rect 27260 5399 28248 6893
rect 28908 7037 29896 8531
rect 30556 8673 31544 10167
rect 32204 10309 33192 11803
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 32204 10275 32318 10309
rect 33102 10275 33192 10309
rect 32204 10201 33192 10275
rect 32204 10167 32318 10201
rect 33102 10167 33192 10201
rect 30556 8639 30660 8673
rect 31444 8639 31544 8673
rect 30556 8565 31544 8639
rect 30556 8531 30660 8565
rect 31444 8531 31544 8565
rect 28908 7003 29002 7037
rect 29786 7003 29896 7037
rect 28908 6927 29896 7003
rect 28908 6893 29002 6927
rect 29786 6893 29896 6927
rect 27260 5365 27344 5399
rect 28128 5365 28248 5399
rect 27260 5291 28248 5365
rect 27260 5257 27344 5291
rect 28128 5257 28248 5291
rect 25566 3729 25686 3763
rect 26470 3729 26554 3763
rect 25566 3655 26554 3729
rect 25566 3621 25686 3655
rect 26470 3621 26554 3655
rect 23918 2093 24028 2127
rect 24812 2093 24906 2127
rect 23918 2019 24906 2093
rect 23918 1985 24028 2019
rect 24812 1985 24906 2019
rect 22260 457 22370 491
rect 23154 457 23248 491
rect 22260 442 23248 457
rect 23918 491 24906 1985
rect 25566 2127 26554 3621
rect 27260 3763 28248 5257
rect 28908 5399 29896 6893
rect 30556 7037 31544 8531
rect 32204 8673 33192 10167
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 32204 8639 32318 8673
rect 33102 8639 33192 8673
rect 32204 8565 33192 8639
rect 32204 8531 32318 8565
rect 33102 8531 33192 8565
rect 30556 7003 30660 7037
rect 31444 7003 31544 7037
rect 30556 6927 31544 7003
rect 30556 6893 30660 6927
rect 31444 6893 31544 6927
rect 28908 5365 29002 5399
rect 29786 5365 29896 5399
rect 28908 5291 29896 5365
rect 28908 5257 29002 5291
rect 29786 5257 29896 5291
rect 27260 3729 27344 3763
rect 28128 3729 28248 3763
rect 27260 3655 28248 3729
rect 27260 3621 27344 3655
rect 28128 3621 28248 3655
rect 25566 2093 25686 2127
rect 26470 2093 26554 2127
rect 25566 2019 26554 2093
rect 25566 1985 25686 2019
rect 26470 1985 26554 2019
rect 23918 457 24028 491
rect 24812 457 24906 491
rect 23918 442 24906 457
rect 25566 491 26554 1985
rect 27260 2127 28248 3621
rect 28908 3763 29896 5257
rect 30556 5399 31544 6893
rect 32204 7037 33192 8531
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 32204 7003 32318 7037
rect 33102 7003 33192 7037
rect 32204 6927 33192 7003
rect 32204 6893 32318 6927
rect 33102 6893 33192 6927
rect 30556 5365 30660 5399
rect 31444 5365 31544 5399
rect 30556 5291 31544 5365
rect 30556 5257 30660 5291
rect 31444 5257 31544 5291
rect 28908 3729 29002 3763
rect 29786 3729 29896 3763
rect 28908 3655 29896 3729
rect 28908 3621 29002 3655
rect 29786 3621 29896 3655
rect 27260 2093 27344 2127
rect 28128 2093 28248 2127
rect 27260 2019 28248 2093
rect 27260 1985 27344 2019
rect 28128 1985 28248 2019
rect 25566 457 25686 491
rect 26470 457 26554 491
rect 25566 442 26554 457
rect 27260 491 28248 1985
rect 28908 2127 29896 3621
rect 30556 3763 31544 5257
rect 32204 5399 33192 6893
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 32204 5365 32318 5399
rect 33102 5365 33192 5399
rect 32204 5291 33192 5365
rect 32204 5257 32318 5291
rect 33102 5257 33192 5291
rect 30556 3729 30660 3763
rect 31444 3729 31544 3763
rect 30556 3655 31544 3729
rect 30556 3621 30660 3655
rect 31444 3621 31544 3655
rect 28908 2093 29002 2127
rect 29786 2093 29896 2127
rect 28908 2019 29896 2093
rect 28908 1985 29002 2019
rect 29786 1985 29896 2019
rect 27260 457 27344 491
rect 28128 457 28248 491
rect 27260 442 28248 457
rect 28908 491 29896 1985
rect 30556 2127 31544 3621
rect 32204 3763 33192 5257
rect 33976 3946 35004 5480
rect 32204 3729 32318 3763
rect 33102 3729 33192 3763
rect 32204 3655 33192 3729
rect 32204 3621 32318 3655
rect 33102 3621 33192 3655
rect 30556 2093 30660 2127
rect 31444 2093 31544 2127
rect 30556 2019 31544 2093
rect 30556 1985 30660 2019
rect 31444 1985 31544 2019
rect 28908 457 29002 491
rect 29786 457 29896 491
rect 28908 442 29896 457
rect 30556 491 31544 1985
rect 32204 2127 33192 3621
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 32204 2093 32318 2127
rect 33102 2093 33192 2127
rect 32204 2019 33192 2093
rect 32204 1985 32318 2019
rect 33102 1985 33192 2019
rect 30556 457 30660 491
rect 31444 457 31544 491
rect 30556 442 31544 457
rect 32204 491 33192 1985
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect 32204 457 32318 491
rect 33102 457 33192 491
rect 32204 442 33192 457
rect 836 436 33192 442
rect 760 318 33192 436
rect 764 308 33192 318
rect 32204 302 33192 308
rect -126 178 20 292
rect -124 138 -30 178
rect 172 177 574 188
rect 168 143 184 177
rect 218 143 376 177
rect 410 143 574 177
rect 172 138 574 143
rect -124 124 -38 138
rect -34586 -54 -734 116
rect -124 90 -94 124
rect -60 90 -38 124
rect -124 70 -38 90
rect 528 132 574 138
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect 528 -312 576 132
rect 33976 52 35004 1480
rect 1532 -54 35054 52
rect 528 -316 578 -312
rect -34586 -828 -734 -520
rect -88 -351 328 -342
rect -88 -385 88 -351
rect 122 -385 280 -351
rect 314 -385 330 -351
rect -88 -404 328 -385
rect -88 -778 -50 -404
rect 530 -462 578 -316
rect 450 -464 578 -462
rect 116 -476 578 -464
rect 116 -510 136 -476
rect 170 -510 328 -476
rect 362 -510 578 -476
rect 116 -516 578 -510
rect 116 -518 456 -516
rect 530 -518 578 -516
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
rect -88 -786 284 -778
rect -88 -820 40 -786
rect 74 -820 232 -786
rect 266 -820 284 -786
rect -88 -830 284 -820
rect -86 -916 518 -900
rect -86 -968 -54 -916
rect 4 -968 346 -916
rect 404 -968 518 -916
rect -86 -982 518 -968
<< viali >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect -32800 16418 -32766 16762
rect -32800 15730 -32766 16418
rect -32800 15386 -32766 15730
rect -31142 16418 -31108 16762
rect -31142 15730 -31108 16418
rect -31142 15386 -31108 15730
rect -34234 13480 -33702 13946
rect -32800 14782 -32766 15126
rect -32800 14094 -32766 14782
rect -32800 13750 -32766 14094
rect -29484 16418 -29450 16762
rect -29484 15730 -29450 16418
rect -29484 15386 -29450 15730
rect -31142 14782 -31108 15126
rect -31142 14094 -31108 14782
rect -31142 13750 -31108 14094
rect -32798 13036 -32764 13380
rect -32798 12348 -32764 13036
rect -32798 12004 -32764 12348
rect -34234 11480 -33702 11946
rect -27826 16418 -27792 16762
rect -27826 15730 -27792 16418
rect -27826 15386 -27792 15730
rect -29484 14782 -29450 15126
rect -29484 14094 -29450 14782
rect -29484 13750 -29450 14094
rect -31140 13036 -31106 13380
rect -31140 12348 -31106 13036
rect -31140 12004 -31106 12348
rect -32798 11400 -32764 11744
rect -32798 10712 -32764 11400
rect -32798 10368 -32764 10712
rect -26168 16418 -26134 16762
rect -26168 15730 -26134 16418
rect -26168 15386 -26134 15730
rect -27826 14782 -27792 15126
rect -27826 14094 -27792 14782
rect -27826 13750 -27792 14094
rect -29482 13036 -29448 13380
rect -29482 12348 -29448 13036
rect -29482 12004 -29448 12348
rect -31140 11400 -31106 11744
rect -31140 10712 -31106 11400
rect -31140 10368 -31106 10712
rect -34234 9480 -33702 9946
rect -32798 9764 -32764 10108
rect -32798 9076 -32764 9764
rect -32798 8732 -32764 9076
rect -24510 16418 -24476 16762
rect -24510 15730 -24476 16418
rect -24510 15386 -24476 15730
rect -26168 14782 -26134 15126
rect -26168 14094 -26134 14782
rect -26168 13750 -26134 14094
rect -27824 13036 -27790 13380
rect -27824 12348 -27790 13036
rect -27824 12004 -27790 12348
rect -29482 11400 -29448 11744
rect -29482 10712 -29448 11400
rect -29482 10368 -29448 10712
rect -31140 9764 -31106 10108
rect -31140 9076 -31106 9764
rect -31140 8732 -31106 9076
rect -34234 7480 -33702 7946
rect -32798 8128 -32764 8472
rect -32798 7440 -32764 8128
rect -32798 7096 -32764 7440
rect -22852 16418 -22818 16762
rect -22852 15730 -22818 16418
rect -22852 15386 -22818 15730
rect -24510 14782 -24476 15126
rect -24510 14094 -24476 14782
rect -24510 13750 -24476 14094
rect -26166 13036 -26132 13380
rect -26166 12348 -26132 13036
rect -26166 12004 -26132 12348
rect -27824 11400 -27790 11744
rect -27824 10712 -27790 11400
rect -27824 10368 -27790 10712
rect -29482 9764 -29448 10108
rect -29482 9076 -29448 9764
rect -29482 8732 -29448 9076
rect -31140 8128 -31106 8472
rect -31140 7440 -31106 8128
rect -31140 7096 -31106 7440
rect -34234 5480 -33702 5946
rect -32798 6490 -32764 6834
rect -32798 5802 -32764 6490
rect -32798 5458 -32764 5802
rect -21194 16418 -21160 16762
rect -21194 15730 -21160 16418
rect -21194 15386 -21160 15730
rect -22852 14782 -22818 15126
rect -22852 14094 -22818 14782
rect -22852 13750 -22818 14094
rect -24508 13036 -24474 13380
rect -24508 12348 -24474 13036
rect -24508 12004 -24474 12348
rect -26166 11400 -26132 11744
rect -26166 10712 -26132 11400
rect -26166 10368 -26132 10712
rect -27824 9764 -27790 10108
rect -27824 9076 -27790 9764
rect -27824 8732 -27790 9076
rect -29482 8128 -29448 8472
rect -29482 7440 -29448 8128
rect -29482 7096 -29448 7440
rect -31140 6490 -31106 6834
rect -31140 5802 -31106 6490
rect -31140 5458 -31106 5802
rect -34234 3480 -33702 3946
rect -32798 4854 -32764 5198
rect -32798 4166 -32764 4854
rect -32798 3822 -32764 4166
rect -19536 16418 -19502 16762
rect -19536 15730 -19502 16418
rect -19536 15386 -19502 15730
rect -21194 14782 -21160 15126
rect -21194 14094 -21160 14782
rect -21194 13750 -21160 14094
rect -22850 13036 -22816 13380
rect -22850 12348 -22816 13036
rect -22850 12004 -22816 12348
rect -24508 11400 -24474 11744
rect -24508 10712 -24474 11400
rect -24508 10368 -24474 10712
rect -26166 9764 -26132 10108
rect -26166 9076 -26132 9764
rect -26166 8732 -26132 9076
rect -27824 8128 -27790 8472
rect -27824 7440 -27790 8128
rect -27824 7096 -27790 7440
rect -29482 6490 -29448 6834
rect -29482 5802 -29448 6490
rect -29482 5458 -29448 5802
rect -31140 4854 -31106 5198
rect -31140 4166 -31106 4854
rect -31140 3822 -31106 4166
rect -32798 3218 -32764 3562
rect -32798 2530 -32764 3218
rect -32798 2186 -32764 2530
rect -34234 1480 -33702 1946
rect -17878 16418 -17844 16762
rect -17878 15730 -17844 16418
rect -17878 15386 -17844 15730
rect -19536 14782 -19502 15126
rect -19536 14094 -19502 14782
rect -19536 13750 -19502 14094
rect -21192 13036 -21158 13380
rect -21192 12348 -21158 13036
rect -21192 12004 -21158 12348
rect -22850 11400 -22816 11744
rect -22850 10712 -22816 11400
rect -22850 10368 -22816 10712
rect -24508 9764 -24474 10108
rect -24508 9076 -24474 9764
rect -24508 8732 -24474 9076
rect -26166 8128 -26132 8472
rect -26166 7440 -26132 8128
rect -26166 7096 -26132 7440
rect -27824 6490 -27790 6834
rect -27824 5802 -27790 6490
rect -27824 5458 -27790 5802
rect -29482 4854 -29448 5198
rect -29482 4166 -29448 4854
rect -29482 3822 -29448 4166
rect -31140 3218 -31106 3562
rect -31140 2530 -31106 3218
rect -31140 2186 -31106 2530
rect -32798 1582 -32764 1926
rect -32798 894 -32764 1582
rect -32798 550 -32764 894
rect -16220 16418 -16186 16762
rect -16220 15730 -16186 16418
rect -16220 15386 -16186 15730
rect -17878 14782 -17844 15126
rect -17878 14094 -17844 14782
rect -17878 13750 -17844 14094
rect -19534 13036 -19500 13380
rect -19534 12348 -19500 13036
rect -19534 12004 -19500 12348
rect -21192 11400 -21158 11744
rect -21192 10712 -21158 11400
rect -21192 10368 -21158 10712
rect -22850 9764 -22816 10108
rect -22850 9076 -22816 9764
rect -22850 8732 -22816 9076
rect -24508 8128 -24474 8472
rect -24508 7440 -24474 8128
rect -24508 7096 -24474 7440
rect -26166 6490 -26132 6834
rect -26166 5802 -26132 6490
rect -26166 5458 -26132 5802
rect -27824 4854 -27790 5198
rect -27824 4166 -27790 4854
rect -27824 3822 -27790 4166
rect -29482 3218 -29448 3562
rect -29482 2530 -29448 3218
rect -29482 2186 -29448 2530
rect -31140 1582 -31106 1926
rect -31140 894 -31106 1582
rect -31140 550 -31106 894
rect -14562 16418 -14528 16762
rect -14562 15730 -14528 16418
rect -14562 15386 -14528 15730
rect -12904 16418 -12870 16762
rect -12904 15730 -12870 16418
rect -12904 15386 -12870 15730
rect -16220 14782 -16186 15126
rect -16220 14094 -16186 14782
rect -16220 13750 -16186 14094
rect -17876 13036 -17842 13380
rect -17876 12348 -17842 13036
rect -17876 12004 -17842 12348
rect -19534 11400 -19500 11744
rect -19534 10712 -19500 11400
rect -19534 10368 -19500 10712
rect -21192 9764 -21158 10108
rect -21192 9076 -21158 9764
rect -21192 8732 -21158 9076
rect -22850 8128 -22816 8472
rect -22850 7440 -22816 8128
rect -22850 7096 -22816 7440
rect -24508 6490 -24474 6834
rect -24508 5802 -24474 6490
rect -24508 5458 -24474 5802
rect -26166 4854 -26132 5198
rect -26166 4166 -26132 4854
rect -26166 3822 -26132 4166
rect -27824 3218 -27790 3562
rect -27824 2530 -27790 3218
rect -27824 2186 -27790 2530
rect -29482 1582 -29448 1926
rect -29482 894 -29448 1582
rect -29482 550 -29448 894
rect -14562 14782 -14528 15126
rect -14562 14094 -14528 14782
rect -14562 13750 -14528 14094
rect -11246 16418 -11212 16762
rect -11246 15730 -11212 16418
rect -11246 15386 -11212 15730
rect -12904 14782 -12870 15126
rect -12904 14094 -12870 14782
rect -12904 13750 -12870 14094
rect -16218 13036 -16184 13380
rect -16218 12348 -16184 13036
rect -16218 12004 -16184 12348
rect -17876 11400 -17842 11744
rect -17876 10712 -17842 11400
rect -17876 10368 -17842 10712
rect -19534 9764 -19500 10108
rect -19534 9076 -19500 9764
rect -19534 8732 -19500 9076
rect -21192 8128 -21158 8472
rect -21192 7440 -21158 8128
rect -21192 7096 -21158 7440
rect -22850 6490 -22816 6834
rect -22850 5802 -22816 6490
rect -22850 5458 -22816 5802
rect -24508 4854 -24474 5198
rect -24508 4166 -24474 4854
rect -24508 3822 -24474 4166
rect -26166 3218 -26132 3562
rect -26166 2530 -26132 3218
rect -26166 2186 -26132 2530
rect -27824 1582 -27790 1926
rect -27824 894 -27790 1582
rect -27824 550 -27790 894
rect -14560 13036 -14526 13380
rect -14560 12348 -14526 13036
rect -14560 12004 -14526 12348
rect -9588 16418 -9554 16762
rect -9588 15730 -9554 16418
rect -9588 15386 -9554 15730
rect -11246 14782 -11212 15126
rect -11246 14094 -11212 14782
rect -11246 13750 -11212 14094
rect -12902 13036 -12868 13380
rect -12902 12348 -12868 13036
rect -12902 12004 -12868 12348
rect -16218 11400 -16184 11744
rect -16218 10712 -16184 11400
rect -16218 10368 -16184 10712
rect -17876 9764 -17842 10108
rect -17876 9076 -17842 9764
rect -17876 8732 -17842 9076
rect -19534 8128 -19500 8472
rect -19534 7440 -19500 8128
rect -19534 7096 -19500 7440
rect -21192 6490 -21158 6834
rect -21192 5802 -21158 6490
rect -21192 5458 -21158 5802
rect -22850 4854 -22816 5198
rect -22850 4166 -22816 4854
rect -22850 3822 -22816 4166
rect -24508 3218 -24474 3562
rect -24508 2530 -24474 3218
rect -24508 2186 -24474 2530
rect -26166 1582 -26132 1926
rect -26166 894 -26132 1582
rect -26166 550 -26132 894
rect -14560 11400 -14526 11744
rect -14560 10712 -14526 11400
rect -14560 10368 -14526 10712
rect -7930 16418 -7896 16762
rect -7930 15730 -7896 16418
rect -7930 15386 -7896 15730
rect -9588 14782 -9554 15126
rect -9588 14094 -9554 14782
rect -9588 13750 -9554 14094
rect -11244 13036 -11210 13380
rect -11244 12348 -11210 13036
rect -11244 12004 -11210 12348
rect -12902 11400 -12868 11744
rect -12902 10712 -12868 11400
rect -12902 10368 -12868 10712
rect -16218 9764 -16184 10108
rect -16218 9076 -16184 9764
rect -16218 8732 -16184 9076
rect -17876 8128 -17842 8472
rect -17876 7440 -17842 8128
rect -17876 7096 -17842 7440
rect -19534 6490 -19500 6834
rect -19534 5802 -19500 6490
rect -19534 5458 -19500 5802
rect -21192 4854 -21158 5198
rect -21192 4166 -21158 4854
rect -21192 3822 -21158 4166
rect -22850 3218 -22816 3562
rect -22850 2530 -22816 3218
rect -22850 2186 -22816 2530
rect -24508 1582 -24474 1926
rect -24508 894 -24474 1582
rect -24508 550 -24474 894
rect -14560 9764 -14526 10108
rect -14560 9076 -14526 9764
rect -14560 8732 -14526 9076
rect -6272 16418 -6238 16762
rect -6272 15730 -6238 16418
rect -6272 15386 -6238 15730
rect -7930 14782 -7896 15126
rect -7930 14094 -7896 14782
rect -7930 13750 -7896 14094
rect -9586 13036 -9552 13380
rect -9586 12348 -9552 13036
rect -9586 12004 -9552 12348
rect -11244 11400 -11210 11744
rect -11244 10712 -11210 11400
rect -11244 10368 -11210 10712
rect -12902 9764 -12868 10108
rect -12902 9076 -12868 9764
rect -12902 8732 -12868 9076
rect -16218 8128 -16184 8472
rect -16218 7440 -16184 8128
rect -16218 7096 -16184 7440
rect -17876 6490 -17842 6834
rect -17876 5802 -17842 6490
rect -17876 5458 -17842 5802
rect -19534 4854 -19500 5198
rect -19534 4166 -19500 4854
rect -19534 3822 -19500 4166
rect -21192 3218 -21158 3562
rect -21192 2530 -21158 3218
rect -21192 2186 -21158 2530
rect -22850 1582 -22816 1926
rect -22850 894 -22816 1582
rect -22850 550 -22816 894
rect -14560 8128 -14526 8472
rect -14560 7440 -14526 8128
rect -14560 7096 -14526 7440
rect -4614 16418 -4580 16762
rect -4614 15730 -4580 16418
rect -4614 15386 -4580 15730
rect -6272 14782 -6238 15126
rect -6272 14094 -6238 14782
rect -6272 13750 -6238 14094
rect -7928 13036 -7894 13380
rect -7928 12348 -7894 13036
rect -7928 12004 -7894 12348
rect -9586 11400 -9552 11744
rect -9586 10712 -9552 11400
rect -9586 10368 -9552 10712
rect -11244 9764 -11210 10108
rect -11244 9076 -11210 9764
rect -11244 8732 -11210 9076
rect -12902 8128 -12868 8472
rect -12902 7440 -12868 8128
rect -12902 7096 -12868 7440
rect -16218 6490 -16184 6834
rect -16218 5802 -16184 6490
rect -16218 5458 -16184 5802
rect -17876 4854 -17842 5198
rect -17876 4166 -17842 4854
rect -17876 3822 -17842 4166
rect -19534 3218 -19500 3562
rect -19534 2530 -19500 3218
rect -19534 2186 -19500 2530
rect -21192 1582 -21158 1926
rect -21192 894 -21158 1582
rect -21192 550 -21158 894
rect -14560 6490 -14526 6834
rect -14560 5802 -14526 6490
rect -14560 5458 -14526 5802
rect -2956 16418 -2922 16762
rect -2956 15730 -2922 16418
rect -2956 15386 -2922 15730
rect -4614 14782 -4580 15126
rect -4614 14094 -4580 14782
rect -4614 13750 -4580 14094
rect -6270 13036 -6236 13380
rect -6270 12348 -6236 13036
rect -6270 12004 -6236 12348
rect -7928 11400 -7894 11744
rect -7928 10712 -7894 11400
rect -7928 10368 -7894 10712
rect -9586 9764 -9552 10108
rect -9586 9076 -9552 9764
rect -9586 8732 -9552 9076
rect -11244 8128 -11210 8472
rect -11244 7440 -11210 8128
rect -11244 7096 -11210 7440
rect -12902 6490 -12868 6834
rect -12902 5802 -12868 6490
rect -12902 5458 -12868 5802
rect -16218 4854 -16184 5198
rect -16218 4166 -16184 4854
rect -16218 3822 -16184 4166
rect -17876 3218 -17842 3562
rect -17876 2530 -17842 3218
rect -17876 2186 -17842 2530
rect -19534 1582 -19500 1926
rect -19534 894 -19500 1582
rect -19534 550 -19500 894
rect -14560 4854 -14526 5198
rect -14560 4166 -14526 4854
rect -14560 3822 -14526 4166
rect -1298 16418 -1264 16762
rect -1298 15730 -1264 16418
rect -1298 15386 -1264 15730
rect -2956 14782 -2922 15126
rect -2956 14094 -2922 14782
rect -2956 13750 -2922 14094
rect -4612 13036 -4578 13380
rect -4612 12348 -4578 13036
rect -4612 12004 -4578 12348
rect -6270 11400 -6236 11744
rect -6270 10712 -6236 11400
rect -6270 10368 -6236 10712
rect -7928 9764 -7894 10108
rect -7928 9076 -7894 9764
rect -7928 8732 -7894 9076
rect -9586 8128 -9552 8472
rect -9586 7440 -9552 8128
rect -9586 7096 -9552 7440
rect -11244 6490 -11210 6834
rect -11244 5802 -11210 6490
rect -11244 5458 -11210 5802
rect -12902 4854 -12868 5198
rect -12902 4166 -12868 4854
rect -12902 3822 -12868 4166
rect -16218 3218 -16184 3562
rect -16218 2530 -16184 3218
rect -16218 2186 -16184 2530
rect -17876 1582 -17842 1926
rect -17876 894 -17842 1582
rect -17876 550 -17842 894
rect -14560 3218 -14526 3562
rect -14560 2530 -14526 3218
rect -14560 2186 -14526 2530
rect 360 16418 394 16762
rect 360 15730 394 16418
rect 360 15386 394 15730
rect -1298 14782 -1264 15126
rect -1298 14094 -1264 14782
rect -1298 13750 -1264 14094
rect -2954 13036 -2920 13380
rect -2954 12348 -2920 13036
rect -2954 12004 -2920 12348
rect -4612 11400 -4578 11744
rect -4612 10712 -4578 11400
rect -4612 10368 -4578 10712
rect -6270 9764 -6236 10108
rect -6270 9076 -6236 9764
rect -6270 8732 -6236 9076
rect -7928 8128 -7894 8472
rect -7928 7440 -7894 8128
rect -7928 7096 -7894 7440
rect -9586 6490 -9552 6834
rect -9586 5802 -9552 6490
rect -9586 5458 -9552 5802
rect -11244 4854 -11210 5198
rect -11244 4166 -11210 4854
rect -11244 3822 -11210 4166
rect -12902 3218 -12868 3562
rect -12902 2530 -12868 3218
rect -12902 2186 -12868 2530
rect -16218 1582 -16184 1926
rect -16218 894 -16184 1582
rect -16218 550 -16184 894
rect -14560 1582 -14526 1926
rect -14560 894 -14526 1582
rect -14560 550 -14526 894
rect 2018 16418 2052 16762
rect 2018 15730 2052 16418
rect 2018 15386 2052 15730
rect 360 14782 394 15126
rect 360 14094 394 14782
rect 360 13750 394 14094
rect -1296 13036 -1262 13380
rect -1296 12348 -1262 13036
rect -1296 12004 -1262 12348
rect -2954 11400 -2920 11744
rect -2954 10712 -2920 11400
rect -2954 10368 -2920 10712
rect -4612 9764 -4578 10108
rect -4612 9076 -4578 9764
rect -4612 8732 -4578 9076
rect -6270 8128 -6236 8472
rect -6270 7440 -6236 8128
rect -6270 7096 -6236 7440
rect -7928 6490 -7894 6834
rect -7928 5802 -7894 6490
rect -7928 5458 -7894 5802
rect -9586 4854 -9552 5198
rect -9586 4166 -9552 4854
rect -9586 3822 -9552 4166
rect -11244 3218 -11210 3562
rect -11244 2530 -11210 3218
rect -11244 2186 -11210 2530
rect -12902 1582 -12868 1926
rect -12902 894 -12868 1582
rect -12902 550 -12868 894
rect 3676 16418 3710 16762
rect 3676 15730 3710 16418
rect 3676 15386 3710 15730
rect 2018 14782 2052 15126
rect 2018 14094 2052 14782
rect 2018 13750 2052 14094
rect 362 13036 396 13380
rect 362 12348 396 13036
rect 362 12004 396 12348
rect -1296 11400 -1262 11744
rect -1296 10712 -1262 11400
rect -1296 10368 -1262 10712
rect -2954 9764 -2920 10108
rect -2954 9076 -2920 9764
rect -2954 8732 -2920 9076
rect -4612 8128 -4578 8472
rect -4612 7440 -4578 8128
rect -4612 7096 -4578 7440
rect -6270 6490 -6236 6834
rect -6270 5802 -6236 6490
rect -6270 5458 -6236 5802
rect -7928 4854 -7894 5198
rect -7928 4166 -7894 4854
rect -7928 3822 -7894 4166
rect -9586 3218 -9552 3562
rect -9586 2530 -9552 3218
rect -9586 2186 -9552 2530
rect -11244 1582 -11210 1926
rect -11244 894 -11210 1582
rect -11244 550 -11210 894
rect 5334 16418 5368 16762
rect 5334 15730 5368 16418
rect 5334 15386 5368 15730
rect 3676 14782 3710 15126
rect 3676 14094 3710 14782
rect 3676 13750 3710 14094
rect 2020 13036 2054 13380
rect 2020 12348 2054 13036
rect 2020 12004 2054 12348
rect 362 11400 396 11744
rect 362 10712 396 11400
rect 362 10368 396 10712
rect -1296 9764 -1262 10108
rect -1296 9076 -1262 9764
rect -1296 8732 -1262 9076
rect -2954 8128 -2920 8472
rect -2954 7440 -2920 8128
rect -2954 7096 -2920 7440
rect -4612 6490 -4578 6834
rect -4612 5802 -4578 6490
rect -4612 5458 -4578 5802
rect -6270 4854 -6236 5198
rect -6270 4166 -6236 4854
rect -6270 3822 -6236 4166
rect -7928 3218 -7894 3562
rect -7928 2530 -7894 3218
rect -7928 2186 -7894 2530
rect -9586 1582 -9552 1926
rect -9586 894 -9552 1582
rect -9586 550 -9552 894
rect 6992 16418 7026 16762
rect 6992 15730 7026 16418
rect 6992 15386 7026 15730
rect 5334 14782 5368 15126
rect 5334 14094 5368 14782
rect 5334 13750 5368 14094
rect 3678 13036 3712 13380
rect 3678 12348 3712 13036
rect 3678 12004 3712 12348
rect 2020 11400 2054 11744
rect 2020 10712 2054 11400
rect 2020 10368 2054 10712
rect 362 9764 396 10108
rect 362 9076 396 9764
rect 362 8732 396 9076
rect -1296 8128 -1262 8472
rect -1296 7440 -1262 8128
rect -1296 7096 -1262 7440
rect -2954 6490 -2920 6834
rect -2954 5802 -2920 6490
rect -2954 5458 -2920 5802
rect -4612 4854 -4578 5198
rect -4612 4166 -4578 4854
rect -4612 3822 -4578 4166
rect -6270 3218 -6236 3562
rect -6270 2530 -6236 3218
rect -6270 2186 -6236 2530
rect -7928 1582 -7894 1926
rect -7928 894 -7894 1582
rect -7928 550 -7894 894
rect 8650 16418 8684 16762
rect 8650 15730 8684 16418
rect 8650 15386 8684 15730
rect 6992 14782 7026 15126
rect 6992 14094 7026 14782
rect 6992 13750 7026 14094
rect 5336 13036 5370 13380
rect 5336 12348 5370 13036
rect 5336 12004 5370 12348
rect 3678 11400 3712 11744
rect 3678 10712 3712 11400
rect 3678 10368 3712 10712
rect 2020 9764 2054 10108
rect 2020 9076 2054 9764
rect 2020 8732 2054 9076
rect 362 8128 396 8472
rect 362 7440 396 8128
rect 362 7096 396 7440
rect -1296 6490 -1262 6834
rect -1296 5802 -1262 6490
rect -1296 5458 -1262 5802
rect -2954 4854 -2920 5198
rect -2954 4166 -2920 4854
rect -2954 3822 -2920 4166
rect -4612 3218 -4578 3562
rect -4612 2530 -4578 3218
rect -4612 2186 -4578 2530
rect -6270 1582 -6236 1926
rect -6270 894 -6236 1582
rect -6270 550 -6236 894
rect 10308 16418 10342 16762
rect 10308 15730 10342 16418
rect 10308 15386 10342 15730
rect 8650 14782 8684 15126
rect 8650 14094 8684 14782
rect 8650 13750 8684 14094
rect 6994 13036 7028 13380
rect 6994 12348 7028 13036
rect 6994 12004 7028 12348
rect 5336 11400 5370 11744
rect 5336 10712 5370 11400
rect 5336 10368 5370 10712
rect 3678 9764 3712 10108
rect 3678 9076 3712 9764
rect 3678 8732 3712 9076
rect 2020 8128 2054 8472
rect 2020 7440 2054 8128
rect 2020 7096 2054 7440
rect 362 6490 396 6834
rect 362 5802 396 6490
rect 362 5458 396 5802
rect -1296 4854 -1262 5198
rect -1296 4166 -1262 4854
rect -1296 3822 -1262 4166
rect -2954 3218 -2920 3562
rect -2954 2530 -2920 3218
rect -2954 2186 -2920 2530
rect -4612 1582 -4578 1926
rect -4612 894 -4578 1582
rect -4612 550 -4578 894
rect 11966 16418 12000 16762
rect 11966 15730 12000 16418
rect 11966 15386 12000 15730
rect 10308 14782 10342 15126
rect 10308 14094 10342 14782
rect 10308 13750 10342 14094
rect 8652 13036 8686 13380
rect 8652 12348 8686 13036
rect 8652 12004 8686 12348
rect 6994 11400 7028 11744
rect 6994 10712 7028 11400
rect 6994 10368 7028 10712
rect 5336 9764 5370 10108
rect 5336 9076 5370 9764
rect 5336 8732 5370 9076
rect 3678 8128 3712 8472
rect 3678 7440 3712 8128
rect 3678 7096 3712 7440
rect 2020 6490 2054 6834
rect 2020 5802 2054 6490
rect 2020 5458 2054 5802
rect 362 4854 396 5198
rect 362 4166 396 4854
rect 362 3822 396 4166
rect -1296 3218 -1262 3562
rect -1296 2530 -1262 3218
rect -1296 2186 -1262 2530
rect -2954 1582 -2920 1926
rect -2954 894 -2920 1582
rect -2954 550 -2920 894
rect 13624 16418 13658 16762
rect 13624 15730 13658 16418
rect 13624 15386 13658 15730
rect 11966 14782 12000 15126
rect 11966 14094 12000 14782
rect 11966 13750 12000 14094
rect 10310 13036 10344 13380
rect 10310 12348 10344 13036
rect 10310 12004 10344 12348
rect 8652 11400 8686 11744
rect 8652 10712 8686 11400
rect 8652 10368 8686 10712
rect 6994 9764 7028 10108
rect 6994 9076 7028 9764
rect 6994 8732 7028 9076
rect 5336 8128 5370 8472
rect 5336 7440 5370 8128
rect 5336 7096 5370 7440
rect 3678 6490 3712 6834
rect 3678 5802 3712 6490
rect 3678 5458 3712 5802
rect 2020 4854 2054 5198
rect 2020 4166 2054 4854
rect 2020 3822 2054 4166
rect 362 3218 396 3562
rect 362 2530 396 3218
rect 362 2186 396 2530
rect -1296 1582 -1262 1926
rect -1296 894 -1262 1582
rect -1296 550 -1262 894
rect 15282 16418 15316 16762
rect 15282 15730 15316 16418
rect 15282 15386 15316 15730
rect 13624 14782 13658 15126
rect 13624 14094 13658 14782
rect 13624 13750 13658 14094
rect 11968 13036 12002 13380
rect 11968 12348 12002 13036
rect 11968 12004 12002 12348
rect 10310 11400 10344 11744
rect 10310 10712 10344 11400
rect 10310 10368 10344 10712
rect 8652 9764 8686 10108
rect 8652 9076 8686 9764
rect 8652 8732 8686 9076
rect 6994 8128 7028 8472
rect 6994 7440 7028 8128
rect 6994 7096 7028 7440
rect 5336 6490 5370 6834
rect 5336 5802 5370 6490
rect 5336 5458 5370 5802
rect 3678 4854 3712 5198
rect 3678 4166 3712 4854
rect 3678 3822 3712 4166
rect 2020 3218 2054 3562
rect 2020 2530 2054 3218
rect 2020 2186 2054 2530
rect 362 1582 396 1926
rect 362 894 396 1582
rect 362 550 396 894
rect 16940 16418 16974 16762
rect 16940 15730 16974 16418
rect 16940 15386 16974 15730
rect 15282 14782 15316 15126
rect 15282 14094 15316 14782
rect 15282 13750 15316 14094
rect 13626 13036 13660 13380
rect 13626 12348 13660 13036
rect 13626 12004 13660 12348
rect 11968 11400 12002 11744
rect 11968 10712 12002 11400
rect 11968 10368 12002 10712
rect 10310 9764 10344 10108
rect 10310 9076 10344 9764
rect 10310 8732 10344 9076
rect 8652 8128 8686 8472
rect 8652 7440 8686 8128
rect 8652 7096 8686 7440
rect 6994 6490 7028 6834
rect 6994 5802 7028 6490
rect 6994 5458 7028 5802
rect 5336 4854 5370 5198
rect 5336 4166 5370 4854
rect 5336 3822 5370 4166
rect 3678 3218 3712 3562
rect 3678 2530 3712 3218
rect 3678 2186 3712 2530
rect 2020 1582 2054 1926
rect 2020 894 2054 1582
rect 2020 550 2054 894
rect 802 457 816 470
rect 816 457 836 470
rect 802 436 836 457
rect 18598 16418 18632 16762
rect 18598 15730 18632 16418
rect 18598 15386 18632 15730
rect 16940 14782 16974 15126
rect 16940 14094 16974 14782
rect 16940 13750 16974 14094
rect 15284 13036 15318 13380
rect 15284 12348 15318 13036
rect 15284 12004 15318 12348
rect 13626 11400 13660 11744
rect 13626 10712 13660 11400
rect 13626 10368 13660 10712
rect 11968 9764 12002 10108
rect 11968 9076 12002 9764
rect 11968 8732 12002 9076
rect 10310 8128 10344 8472
rect 10310 7440 10344 8128
rect 10310 7096 10344 7440
rect 8652 6490 8686 6834
rect 8652 5802 8686 6490
rect 8652 5458 8686 5802
rect 6994 4854 7028 5198
rect 6994 4166 7028 4854
rect 6994 3822 7028 4166
rect 5336 3218 5370 3562
rect 5336 2530 5370 3218
rect 5336 2186 5370 2530
rect 3678 1582 3712 1926
rect 3678 894 3712 1582
rect 3678 550 3712 894
rect 20256 16418 20290 16762
rect 20256 15730 20290 16418
rect 20256 15386 20290 15730
rect 18598 14782 18632 15126
rect 18598 14094 18632 14782
rect 18598 13750 18632 14094
rect 16942 13036 16976 13380
rect 16942 12348 16976 13036
rect 16942 12004 16976 12348
rect 15284 11400 15318 11744
rect 15284 10712 15318 11400
rect 15284 10368 15318 10712
rect 13626 9764 13660 10108
rect 13626 9076 13660 9764
rect 13626 8732 13660 9076
rect 11968 8128 12002 8472
rect 11968 7440 12002 8128
rect 11968 7096 12002 7440
rect 10310 6490 10344 6834
rect 10310 5802 10344 6490
rect 10310 5458 10344 5802
rect 8652 4854 8686 5198
rect 8652 4166 8686 4854
rect 8652 3822 8686 4166
rect 6994 3218 7028 3562
rect 6994 2530 7028 3218
rect 6994 2186 7028 2530
rect 5336 1582 5370 1926
rect 5336 894 5370 1582
rect 5336 550 5370 894
rect 21914 16418 21948 16762
rect 21914 15730 21948 16418
rect 21914 15386 21948 15730
rect 20256 14782 20290 15126
rect 20256 14094 20290 14782
rect 20256 13750 20290 14094
rect 18600 13036 18634 13380
rect 18600 12348 18634 13036
rect 18600 12004 18634 12348
rect 16942 11400 16976 11744
rect 16942 10712 16976 11400
rect 16942 10368 16976 10712
rect 15284 9764 15318 10108
rect 15284 9076 15318 9764
rect 15284 8732 15318 9076
rect 13626 8128 13660 8472
rect 13626 7440 13660 8128
rect 13626 7096 13660 7440
rect 11968 6490 12002 6834
rect 11968 5802 12002 6490
rect 11968 5458 12002 5802
rect 10310 4854 10344 5198
rect 10310 4166 10344 4854
rect 10310 3822 10344 4166
rect 8652 3218 8686 3562
rect 8652 2530 8686 3218
rect 8652 2186 8686 2530
rect 6994 1582 7028 1926
rect 6994 894 7028 1582
rect 6994 550 7028 894
rect 23572 16418 23606 16762
rect 23572 15730 23606 16418
rect 23572 15386 23606 15730
rect 21914 14782 21948 15126
rect 21914 14094 21948 14782
rect 21914 13750 21948 14094
rect 20258 13036 20292 13380
rect 20258 12348 20292 13036
rect 20258 12004 20292 12348
rect 18600 11400 18634 11744
rect 18600 10712 18634 11400
rect 18600 10368 18634 10712
rect 16942 9764 16976 10108
rect 16942 9076 16976 9764
rect 16942 8732 16976 9076
rect 15284 8128 15318 8472
rect 15284 7440 15318 8128
rect 15284 7096 15318 7440
rect 13626 6490 13660 6834
rect 13626 5802 13660 6490
rect 13626 5458 13660 5802
rect 11968 4854 12002 5198
rect 11968 4166 12002 4854
rect 11968 3822 12002 4166
rect 10310 3218 10344 3562
rect 10310 2530 10344 3218
rect 10310 2186 10344 2530
rect 8652 1582 8686 1926
rect 8652 894 8686 1582
rect 8652 550 8686 894
rect 25230 16418 25264 16762
rect 25230 15730 25264 16418
rect 25230 15386 25264 15730
rect 23572 14782 23606 15126
rect 23572 14094 23606 14782
rect 23572 13750 23606 14094
rect 21916 13036 21950 13380
rect 21916 12348 21950 13036
rect 21916 12004 21950 12348
rect 20258 11400 20292 11744
rect 20258 10712 20292 11400
rect 20258 10368 20292 10712
rect 18600 9764 18634 10108
rect 18600 9076 18634 9764
rect 18600 8732 18634 9076
rect 16942 8128 16976 8472
rect 16942 7440 16976 8128
rect 16942 7096 16976 7440
rect 15284 6490 15318 6834
rect 15284 5802 15318 6490
rect 15284 5458 15318 5802
rect 13626 4854 13660 5198
rect 13626 4166 13660 4854
rect 13626 3822 13660 4166
rect 11968 3218 12002 3562
rect 11968 2530 12002 3218
rect 11968 2186 12002 2530
rect 10310 1582 10344 1926
rect 10310 894 10344 1582
rect 10310 550 10344 894
rect 26888 16418 26922 16762
rect 26888 15730 26922 16418
rect 26888 15386 26922 15730
rect 25230 14782 25264 15126
rect 25230 14094 25264 14782
rect 25230 13750 25264 14094
rect 23574 13036 23608 13380
rect 23574 12348 23608 13036
rect 23574 12004 23608 12348
rect 21916 11400 21950 11744
rect 21916 10712 21950 11400
rect 21916 10368 21950 10712
rect 20258 9764 20292 10108
rect 20258 9076 20292 9764
rect 20258 8732 20292 9076
rect 18600 8128 18634 8472
rect 18600 7440 18634 8128
rect 18600 7096 18634 7440
rect 16942 6490 16976 6834
rect 16942 5802 16976 6490
rect 16942 5458 16976 5802
rect 15284 4854 15318 5198
rect 15284 4166 15318 4854
rect 15284 3822 15318 4166
rect 13626 3218 13660 3562
rect 13626 2530 13660 3218
rect 13626 2186 13660 2530
rect 11968 1582 12002 1926
rect 11968 894 12002 1582
rect 11968 550 12002 894
rect 28546 16418 28580 16762
rect 28546 15730 28580 16418
rect 28546 15386 28580 15730
rect 26888 14782 26922 15126
rect 26888 14094 26922 14782
rect 26888 13750 26922 14094
rect 25232 13036 25266 13380
rect 25232 12348 25266 13036
rect 25232 12004 25266 12348
rect 23574 11400 23608 11744
rect 23574 10712 23608 11400
rect 23574 10368 23608 10712
rect 21916 9764 21950 10108
rect 21916 9076 21950 9764
rect 21916 8732 21950 9076
rect 20258 8128 20292 8472
rect 20258 7440 20292 8128
rect 20258 7096 20292 7440
rect 18600 6490 18634 6834
rect 18600 5802 18634 6490
rect 18600 5458 18634 5802
rect 16942 4854 16976 5198
rect 16942 4166 16976 4854
rect 16942 3822 16976 4166
rect 15284 3218 15318 3562
rect 15284 2530 15318 3218
rect 15284 2186 15318 2530
rect 13626 1582 13660 1926
rect 13626 894 13660 1582
rect 13626 550 13660 894
rect 30204 16418 30238 16762
rect 30204 15730 30238 16418
rect 30204 15386 30238 15730
rect 28546 14782 28580 15126
rect 28546 14094 28580 14782
rect 28546 13750 28580 14094
rect 26890 13036 26924 13380
rect 26890 12348 26924 13036
rect 26890 12004 26924 12348
rect 25232 11400 25266 11744
rect 25232 10712 25266 11400
rect 25232 10368 25266 10712
rect 23574 9764 23608 10108
rect 23574 9076 23608 9764
rect 23574 8732 23608 9076
rect 21916 8128 21950 8472
rect 21916 7440 21950 8128
rect 21916 7096 21950 7440
rect 20258 6490 20292 6834
rect 20258 5802 20292 6490
rect 20258 5458 20292 5802
rect 18600 4854 18634 5198
rect 18600 4166 18634 4854
rect 18600 3822 18634 4166
rect 16942 3218 16976 3562
rect 16942 2530 16976 3218
rect 16942 2186 16976 2530
rect 15284 1582 15318 1926
rect 15284 894 15318 1582
rect 15284 550 15318 894
rect 31862 16418 31896 16762
rect 31862 15730 31896 16418
rect 31862 15386 31896 15730
rect 30204 14782 30238 15126
rect 30204 14094 30238 14782
rect 30204 13750 30238 14094
rect 28548 13036 28582 13380
rect 28548 12348 28582 13036
rect 28548 12004 28582 12348
rect 26890 11400 26924 11744
rect 26890 10712 26924 11400
rect 26890 10368 26924 10712
rect 25232 9764 25266 10108
rect 25232 9076 25266 9764
rect 25232 8732 25266 9076
rect 23574 8128 23608 8472
rect 23574 7440 23608 8128
rect 23574 7096 23608 7440
rect 21916 6490 21950 6834
rect 21916 5802 21950 6490
rect 21916 5458 21950 5802
rect 20258 4854 20292 5198
rect 20258 4166 20292 4854
rect 20258 3822 20292 4166
rect 18600 3218 18634 3562
rect 18600 2530 18634 3218
rect 18600 2186 18634 2530
rect 16942 1582 16976 1926
rect 16942 894 16976 1582
rect 16942 550 16976 894
rect 33520 16418 33554 16762
rect 33520 15730 33554 16418
rect 33520 15386 33554 15730
rect 34166 15480 34698 15946
rect 31862 14782 31896 15126
rect 31862 14094 31896 14782
rect 31862 13750 31896 14094
rect 30206 13036 30240 13380
rect 30206 12348 30240 13036
rect 30206 12004 30240 12348
rect 28548 11400 28582 11744
rect 28548 10712 28582 11400
rect 28548 10368 28582 10712
rect 26890 9764 26924 10108
rect 26890 9076 26924 9764
rect 26890 8732 26924 9076
rect 25232 8128 25266 8472
rect 25232 7440 25266 8128
rect 25232 7096 25266 7440
rect 23574 6490 23608 6834
rect 23574 5802 23608 6490
rect 23574 5458 23608 5802
rect 21916 4854 21950 5198
rect 21916 4166 21950 4854
rect 21916 3822 21950 4166
rect 20258 3218 20292 3562
rect 20258 2530 20292 3218
rect 20258 2186 20292 2530
rect 18600 1582 18634 1926
rect 18600 894 18634 1582
rect 18600 550 18634 894
rect 33520 14782 33554 15126
rect 33520 14094 33554 14782
rect 33520 13750 33554 14094
rect 31864 13036 31898 13380
rect 31864 12348 31898 13036
rect 31864 12004 31898 12348
rect 30206 11400 30240 11744
rect 30206 10712 30240 11400
rect 30206 10368 30240 10712
rect 28548 9764 28582 10108
rect 28548 9076 28582 9764
rect 28548 8732 28582 9076
rect 26890 8128 26924 8472
rect 26890 7440 26924 8128
rect 26890 7096 26924 7440
rect 25232 6490 25266 6834
rect 25232 5802 25266 6490
rect 25232 5458 25266 5802
rect 23574 4854 23608 5198
rect 23574 4166 23608 4854
rect 23574 3822 23608 4166
rect 21916 3218 21950 3562
rect 21916 2530 21950 3218
rect 21916 2186 21950 2530
rect 20258 1582 20292 1926
rect 20258 894 20292 1582
rect 20258 550 20292 894
rect 34166 13480 34698 13946
rect 33522 13036 33556 13380
rect 33522 12348 33556 13036
rect 33522 12004 33556 12348
rect 31864 11400 31898 11744
rect 31864 10712 31898 11400
rect 31864 10368 31898 10712
rect 30206 9764 30240 10108
rect 30206 9076 30240 9764
rect 30206 8732 30240 9076
rect 28548 8128 28582 8472
rect 28548 7440 28582 8128
rect 28548 7096 28582 7440
rect 26890 6490 26924 6834
rect 26890 5802 26924 6490
rect 26890 5458 26924 5802
rect 25232 4854 25266 5198
rect 25232 4166 25266 4854
rect 25232 3822 25266 4166
rect 23574 3218 23608 3562
rect 23574 2530 23608 3218
rect 23574 2186 23608 2530
rect 21916 1582 21950 1926
rect 21916 894 21950 1582
rect 21916 550 21950 894
rect 33522 11400 33556 11744
rect 33522 10712 33556 11400
rect 33522 10368 33556 10712
rect 34166 11480 34698 11946
rect 31864 9764 31898 10108
rect 31864 9076 31898 9764
rect 31864 8732 31898 9076
rect 30206 8128 30240 8472
rect 30206 7440 30240 8128
rect 30206 7096 30240 7440
rect 28548 6490 28582 6834
rect 28548 5802 28582 6490
rect 28548 5458 28582 5802
rect 26890 4854 26924 5198
rect 26890 4166 26924 4854
rect 26890 3822 26924 4166
rect 25232 3218 25266 3562
rect 25232 2530 25266 3218
rect 25232 2186 25266 2530
rect 23574 1582 23608 1926
rect 23574 894 23608 1582
rect 23574 550 23608 894
rect 33522 9764 33556 10108
rect 33522 9076 33556 9764
rect 33522 8732 33556 9076
rect 34166 9480 34698 9946
rect 31864 8128 31898 8472
rect 31864 7440 31898 8128
rect 31864 7096 31898 7440
rect 30206 6490 30240 6834
rect 30206 5802 30240 6490
rect 30206 5458 30240 5802
rect 28548 4854 28582 5198
rect 28548 4166 28582 4854
rect 28548 3822 28582 4166
rect 26890 3218 26924 3562
rect 26890 2530 26924 3218
rect 26890 2186 26924 2530
rect 25232 1582 25266 1926
rect 25232 894 25266 1582
rect 25232 550 25266 894
rect 33522 8128 33556 8472
rect 33522 7440 33556 8128
rect 33522 7096 33556 7440
rect 34166 7480 34698 7946
rect 31864 6490 31898 6834
rect 31864 5802 31898 6490
rect 31864 5458 31898 5802
rect 30206 4854 30240 5198
rect 30206 4166 30240 4854
rect 30206 3822 30240 4166
rect 28548 3218 28582 3562
rect 28548 2530 28582 3218
rect 28548 2186 28582 2530
rect 26890 1582 26924 1926
rect 26890 894 26924 1582
rect 26890 550 26924 894
rect 33522 6490 33556 6834
rect 33522 5802 33556 6490
rect 33522 5458 33556 5802
rect 34166 5480 34698 5946
rect 31864 4854 31898 5198
rect 31864 4166 31898 4854
rect 31864 3822 31898 4166
rect 30206 3218 30240 3562
rect 30206 2530 30240 3218
rect 30206 2186 30240 2530
rect 28548 1582 28582 1926
rect 28548 894 28582 1582
rect 28548 550 28582 894
rect 33522 4854 33556 5198
rect 33522 4166 33556 4854
rect 33522 3822 33556 4166
rect 31864 3218 31898 3562
rect 31864 2530 31898 3218
rect 31864 2186 31898 2530
rect 30206 1582 30240 1926
rect 30206 894 30240 1582
rect 30206 550 30240 894
rect 33522 3218 33556 3562
rect 33522 2530 33556 3218
rect 33522 2186 33556 2530
rect 34166 3480 34698 3946
rect 31864 1582 31898 1926
rect 31864 894 31898 1582
rect 31864 550 31898 894
rect 33522 1582 33556 1926
rect 33522 894 33556 1582
rect 33522 550 33556 894
rect 34166 1480 34698 1946
rect -94 90 -60 124
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 40 -10 74 84
rect 40 -198 74 -10
rect 40 -292 74 -198
rect 136 -10 170 84
rect 136 -198 170 -10
rect 136 -292 170 -198
rect 232 -10 266 84
rect 232 -198 266 -10
rect 232 -292 266 -198
rect 328 -10 362 84
rect 328 -198 362 -10
rect 328 -292 362 -198
rect 424 -10 458 84
rect 424 -198 458 -10
rect 424 -292 458 -198
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
rect -8 -604 26 -560
rect -8 -692 26 -604
rect -8 -736 26 -692
rect 88 -604 122 -560
rect 88 -692 122 -604
rect 88 -736 122 -692
rect 184 -604 218 -560
rect 184 -692 218 -604
rect 184 -736 218 -692
rect 280 -604 314 -560
rect 280 -692 314 -604
rect 280 -736 314 -692
rect 376 -604 410 -560
rect 376 -692 410 -604
rect 376 -736 410 -692
rect -54 -968 4 -916
rect 346 -968 404 -916
<< metal1 >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect 178 17330 548 17406
rect 176 17314 548 17330
rect -32806 16762 -32760 16774
rect -32806 16710 -32800 16762
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect -32980 15386 -32800 16710
rect -32766 16710 -32760 16762
rect -31148 16762 -31102 16774
rect -31148 16710 -31142 16762
rect -32766 15386 -31142 16710
rect -31108 16710 -31102 16762
rect -29490 16762 -29444 16774
rect -29490 16710 -29484 16762
rect -31108 15386 -29484 16710
rect -29450 16710 -29444 16762
rect -27832 16762 -27786 16774
rect -27832 16710 -27826 16762
rect -29450 15386 -27826 16710
rect -27792 16710 -27786 16762
rect -26174 16762 -26128 16774
rect -26174 16710 -26168 16762
rect -27792 15386 -26168 16710
rect -26134 16710 -26128 16762
rect -24516 16762 -24470 16774
rect -24516 16710 -24510 16762
rect -26134 15386 -24510 16710
rect -24476 16710 -24470 16762
rect -22858 16762 -22812 16774
rect -22858 16710 -22852 16762
rect -24476 15386 -22852 16710
rect -22818 16710 -22812 16762
rect -21200 16762 -21154 16774
rect -21200 16710 -21194 16762
rect -22818 15386 -21194 16710
rect -21160 16710 -21154 16762
rect -19542 16762 -19496 16774
rect -19542 16710 -19536 16762
rect -21160 15386 -19536 16710
rect -19502 16710 -19496 16762
rect -17884 16762 -17838 16774
rect -17884 16710 -17878 16762
rect -19502 15386 -17878 16710
rect -17844 16710 -17838 16762
rect -16226 16762 -16180 16774
rect -16226 16710 -16220 16762
rect -17844 15386 -16220 16710
rect -16186 16710 -16180 16762
rect -14568 16762 -14522 16774
rect -14568 16710 -14562 16762
rect -16186 15386 -14562 16710
rect -14528 16710 -14522 16762
rect -12910 16762 -12864 16774
rect -12910 16710 -12904 16762
rect -14528 15386 -12904 16710
rect -12870 16710 -12864 16762
rect -11252 16762 -11206 16774
rect -11252 16710 -11246 16762
rect -12870 15386 -11246 16710
rect -11212 16710 -11206 16762
rect -9594 16762 -9548 16774
rect -9594 16710 -9588 16762
rect -11212 15386 -9588 16710
rect -9554 16710 -9548 16762
rect -7936 16762 -7890 16774
rect -7936 16710 -7930 16762
rect -9554 15386 -7930 16710
rect -7896 16710 -7890 16762
rect -6278 16762 -6232 16774
rect -6278 16710 -6272 16762
rect -7896 15386 -6272 16710
rect -6238 16710 -6232 16762
rect -4620 16762 -4574 16774
rect -4620 16710 -4614 16762
rect -6238 15386 -4614 16710
rect -4580 16710 -4574 16762
rect -2962 16762 -2916 16774
rect -2962 16710 -2956 16762
rect -4580 15386 -2956 16710
rect -2922 16710 -2916 16762
rect -1304 16762 -1258 16774
rect -1304 16710 -1298 16762
rect -2922 15386 -1298 16710
rect -1264 16710 -1258 16762
rect 176 16762 544 17314
rect 176 16710 360 16762
rect -1264 15386 360 16710
rect 394 16710 544 16762
rect 2012 16762 2058 16774
rect 2012 16710 2018 16762
rect 394 15386 2018 16710
rect 2052 16710 2058 16762
rect 3670 16762 3716 16774
rect 3670 16710 3676 16762
rect 2052 15386 3676 16710
rect 3710 16710 3716 16762
rect 5328 16762 5374 16774
rect 5328 16710 5334 16762
rect 3710 15386 5334 16710
rect 5368 16710 5374 16762
rect 6986 16762 7032 16774
rect 6986 16710 6992 16762
rect 5368 15386 6992 16710
rect 7026 16710 7032 16762
rect 8644 16762 8690 16774
rect 8644 16710 8650 16762
rect 7026 15386 8650 16710
rect 8684 16710 8690 16762
rect 10302 16762 10348 16774
rect 10302 16710 10308 16762
rect 8684 15386 10308 16710
rect 10342 16710 10348 16762
rect 11960 16762 12006 16774
rect 11960 16710 11966 16762
rect 10342 15386 11966 16710
rect 12000 16710 12006 16762
rect 13618 16762 13664 16774
rect 13618 16710 13624 16762
rect 12000 15386 13624 16710
rect 13658 16710 13664 16762
rect 15276 16762 15322 16774
rect 15276 16710 15282 16762
rect 13658 15386 15282 16710
rect 15316 16710 15322 16762
rect 16934 16762 16980 16774
rect 16934 16710 16940 16762
rect 15316 15386 16940 16710
rect 16974 16710 16980 16762
rect 18592 16762 18638 16774
rect 18592 16710 18598 16762
rect 16974 15386 18598 16710
rect 18632 16710 18638 16762
rect 20250 16762 20296 16774
rect 20250 16710 20256 16762
rect 18632 15386 20256 16710
rect 20290 16710 20296 16762
rect 21908 16762 21954 16774
rect 21908 16710 21914 16762
rect 20290 15386 21914 16710
rect 21948 16710 21954 16762
rect 23566 16762 23612 16774
rect 23566 16710 23572 16762
rect 21948 15386 23572 16710
rect 23606 16710 23612 16762
rect 25224 16762 25270 16774
rect 25224 16710 25230 16762
rect 23606 15386 25230 16710
rect 25264 16710 25270 16762
rect 26882 16762 26928 16774
rect 26882 16710 26888 16762
rect 25264 15386 26888 16710
rect 26922 16710 26928 16762
rect 28540 16762 28586 16774
rect 28540 16710 28546 16762
rect 26922 15386 28546 16710
rect 28580 16710 28586 16762
rect 30198 16762 30244 16774
rect 30198 16710 30204 16762
rect 28580 15386 30204 16710
rect 30238 16710 30244 16762
rect 31856 16762 31902 16774
rect 31856 16710 31862 16762
rect 30238 15386 31862 16710
rect 31896 16710 31902 16762
rect 33514 16762 33560 16774
rect 33514 16710 33520 16762
rect 31896 15386 33520 16710
rect 33554 16710 33560 16762
rect 33554 15386 33630 16710
rect -32980 15126 33630 15386
rect -32980 13750 -32800 15126
rect -32766 13750 -31142 15126
rect -31108 13750 -29484 15126
rect -29450 13750 -27826 15126
rect -27792 13750 -26168 15126
rect -26134 13750 -24510 15126
rect -24476 13750 -22852 15126
rect -22818 13750 -21194 15126
rect -21160 13750 -19536 15126
rect -19502 13750 -17878 15126
rect -17844 13750 -16220 15126
rect -16186 13750 -14562 15126
rect -14528 13750 -12904 15126
rect -12870 13750 -11246 15126
rect -11212 13750 -9588 15126
rect -9554 13750 -7930 15126
rect -7896 13750 -6272 15126
rect -6238 13750 -4614 15126
rect -4580 13750 -2956 15126
rect -2922 13750 -1298 15126
rect -1264 13750 360 15126
rect 394 13750 2018 15126
rect 2052 13750 3676 15126
rect 3710 13750 5334 15126
rect 5368 13750 6992 15126
rect 7026 13750 8650 15126
rect 8684 13750 10308 15126
rect 10342 13750 11966 15126
rect 12000 13750 13624 15126
rect 13658 13750 15282 15126
rect 15316 13750 16940 15126
rect 16974 13750 18598 15126
rect 18632 13750 20256 15126
rect 20290 13750 21914 15126
rect 21948 13750 23572 15126
rect 23606 13750 25230 15126
rect 25264 13750 26888 15126
rect 26922 13750 28546 15126
rect 28580 13750 30204 15126
rect 30238 13750 31862 15126
rect 31896 13750 33520 15126
rect 33554 13750 33630 15126
rect -32980 13380 33630 13750
rect -32980 12004 -32798 13380
rect -32764 12004 -31140 13380
rect -31106 12004 -29482 13380
rect -29448 12004 -27824 13380
rect -27790 12004 -26166 13380
rect -26132 12004 -24508 13380
rect -24474 12004 -22850 13380
rect -22816 12004 -21192 13380
rect -21158 12004 -19534 13380
rect -19500 12004 -17876 13380
rect -17842 12004 -16218 13380
rect -16184 12004 -14560 13380
rect -14526 12004 -12902 13380
rect -12868 12004 -11244 13380
rect -11210 12004 -9586 13380
rect -9552 12004 -7928 13380
rect -7894 12004 -6270 13380
rect -6236 12004 -4612 13380
rect -4578 12004 -2954 13380
rect -2920 12004 -1296 13380
rect -1262 12004 362 13380
rect 396 12004 2020 13380
rect 2054 12004 3678 13380
rect 3712 12004 5336 13380
rect 5370 12004 6994 13380
rect 7028 12004 8652 13380
rect 8686 12004 10310 13380
rect 10344 12004 11968 13380
rect 12002 12004 13626 13380
rect 13660 12004 15284 13380
rect 15318 12004 16942 13380
rect 16976 12004 18600 13380
rect 18634 12004 20258 13380
rect 20292 12004 21916 13380
rect 21950 12004 23574 13380
rect 23608 12004 25232 13380
rect 25266 12004 26890 13380
rect 26924 12004 28548 13380
rect 28582 12004 30206 13380
rect 30240 12004 31864 13380
rect 31898 12004 33522 13380
rect 33556 12004 33630 13380
rect -32980 11744 33630 12004
rect -32980 10368 -32798 11744
rect -32764 10368 -31140 11744
rect -31106 10368 -29482 11744
rect -29448 10368 -27824 11744
rect -27790 10368 -26166 11744
rect -26132 10368 -24508 11744
rect -24474 10368 -22850 11744
rect -22816 10368 -21192 11744
rect -21158 10368 -19534 11744
rect -19500 10368 -17876 11744
rect -17842 10368 -16218 11744
rect -16184 10368 -14560 11744
rect -14526 10368 -12902 11744
rect -12868 10368 -11244 11744
rect -11210 10368 -9586 11744
rect -9552 10368 -7928 11744
rect -7894 10368 -6270 11744
rect -6236 10368 -4612 11744
rect -4578 10368 -2954 11744
rect -2920 10368 -1296 11744
rect -1262 10368 362 11744
rect 396 10368 2020 11744
rect 2054 10368 3678 11744
rect 3712 10368 5336 11744
rect 5370 10368 6994 11744
rect 7028 10368 8652 11744
rect 8686 10368 10310 11744
rect 10344 10368 11968 11744
rect 12002 10368 13626 11744
rect 13660 10368 15284 11744
rect 15318 10368 16942 11744
rect 16976 10368 18600 11744
rect 18634 10368 20258 11744
rect 20292 10368 21916 11744
rect 21950 10368 23574 11744
rect 23608 10368 25232 11744
rect 25266 10368 26890 11744
rect 26924 10368 28548 11744
rect 28582 10368 30206 11744
rect 30240 10368 31864 11744
rect 31898 10368 33522 11744
rect 33556 10368 33630 11744
rect -32980 10108 33630 10368
rect -32980 8732 -32798 10108
rect -32764 8732 -31140 10108
rect -31106 8732 -29482 10108
rect -29448 8732 -27824 10108
rect -27790 8732 -26166 10108
rect -26132 8732 -24508 10108
rect -24474 8732 -22850 10108
rect -22816 8732 -21192 10108
rect -21158 8732 -19534 10108
rect -19500 8732 -17876 10108
rect -17842 8732 -16218 10108
rect -16184 8732 -14560 10108
rect -14526 8732 -12902 10108
rect -12868 8732 -11244 10108
rect -11210 8732 -9586 10108
rect -9552 8732 -7928 10108
rect -7894 8732 -6270 10108
rect -6236 8732 -4612 10108
rect -4578 8732 -2954 10108
rect -2920 8732 -1296 10108
rect -1262 8732 362 10108
rect 396 8732 2020 10108
rect 2054 8732 3678 10108
rect 3712 8732 5336 10108
rect 5370 8732 6994 10108
rect 7028 8732 8652 10108
rect 8686 8732 10310 10108
rect 10344 8732 11968 10108
rect 12002 8732 13626 10108
rect 13660 8732 15284 10108
rect 15318 8732 16942 10108
rect 16976 8732 18600 10108
rect 18634 8732 20258 10108
rect 20292 8732 21916 10108
rect 21950 8732 23574 10108
rect 23608 8732 25232 10108
rect 25266 8732 26890 10108
rect 26924 8732 28548 10108
rect 28582 8732 30206 10108
rect 30240 8732 31864 10108
rect 31898 8732 33522 10108
rect 33556 8732 33630 10108
rect -32980 8472 33630 8732
rect -32980 7096 -32798 8472
rect -32764 7096 -31140 8472
rect -31106 7096 -29482 8472
rect -29448 7096 -27824 8472
rect -27790 7096 -26166 8472
rect -26132 7096 -24508 8472
rect -24474 7096 -22850 8472
rect -22816 7096 -21192 8472
rect -21158 7096 -19534 8472
rect -19500 7096 -17876 8472
rect -17842 7096 -16218 8472
rect -16184 7096 -14560 8472
rect -14526 7096 -12902 8472
rect -12868 7096 -11244 8472
rect -11210 7096 -9586 8472
rect -9552 7096 -7928 8472
rect -7894 7096 -6270 8472
rect -6236 7096 -4612 8472
rect -4578 7096 -2954 8472
rect -2920 7096 -1296 8472
rect -1262 7096 362 8472
rect 396 7096 2020 8472
rect 2054 7096 3678 8472
rect 3712 7096 5336 8472
rect 5370 7096 6994 8472
rect 7028 7096 8652 8472
rect 8686 7096 10310 8472
rect 10344 7096 11968 8472
rect 12002 7096 13626 8472
rect 13660 7096 15284 8472
rect 15318 7096 16942 8472
rect 16976 7096 18600 8472
rect 18634 7096 20258 8472
rect 20292 7096 21916 8472
rect 21950 7096 23574 8472
rect 23608 7096 25232 8472
rect 25266 7096 26890 8472
rect 26924 7096 28548 8472
rect 28582 7096 30206 8472
rect 30240 7096 31864 8472
rect 31898 7096 33522 8472
rect 33556 7096 33630 8472
rect -32980 6834 33630 7096
rect -32980 5458 -32798 6834
rect -32764 5458 -31140 6834
rect -31106 5458 -29482 6834
rect -29448 5458 -27824 6834
rect -27790 5458 -26166 6834
rect -26132 5458 -24508 6834
rect -24474 5458 -22850 6834
rect -22816 5458 -21192 6834
rect -21158 5458 -19534 6834
rect -19500 5458 -17876 6834
rect -17842 5458 -16218 6834
rect -16184 5458 -14560 6834
rect -14526 5458 -12902 6834
rect -12868 5458 -11244 6834
rect -11210 5458 -9586 6834
rect -9552 5458 -7928 6834
rect -7894 5458 -6270 6834
rect -6236 5458 -4612 6834
rect -4578 5458 -2954 6834
rect -2920 5458 -1296 6834
rect -1262 5458 362 6834
rect 396 5458 2020 6834
rect 2054 5458 3678 6834
rect 3712 5458 5336 6834
rect 5370 5458 6994 6834
rect 7028 5458 8652 6834
rect 8686 5458 10310 6834
rect 10344 5458 11968 6834
rect 12002 5458 13626 6834
rect 13660 5458 15284 6834
rect 15318 5458 16942 6834
rect 16976 5458 18600 6834
rect 18634 5458 20258 6834
rect 20292 5458 21916 6834
rect 21950 5458 23574 6834
rect 23608 5458 25232 6834
rect 25266 5458 26890 6834
rect 26924 5458 28548 6834
rect 28582 5458 30206 6834
rect 30240 5458 31864 6834
rect 31898 5458 33522 6834
rect 33556 5458 33630 6834
rect -32980 5198 33630 5458
rect -32980 3822 -32798 5198
rect -32764 3822 -31140 5198
rect -31106 3822 -29482 5198
rect -29448 3822 -27824 5198
rect -27790 3822 -26166 5198
rect -26132 3822 -24508 5198
rect -24474 3822 -22850 5198
rect -22816 3822 -21192 5198
rect -21158 3822 -19534 5198
rect -19500 3822 -17876 5198
rect -17842 3822 -16218 5198
rect -16184 3822 -14560 5198
rect -14526 3822 -12902 5198
rect -12868 3822 -11244 5198
rect -11210 3822 -9586 5198
rect -9552 3822 -7928 5198
rect -7894 3822 -6270 5198
rect -6236 3822 -4612 5198
rect -4578 3822 -2954 5198
rect -2920 3822 -1296 5198
rect -1262 3822 362 5198
rect 396 3822 2020 5198
rect 2054 3822 3678 5198
rect 3712 3822 5336 5198
rect 5370 3822 6994 5198
rect 7028 3822 8652 5198
rect 8686 3822 10310 5198
rect 10344 3822 11968 5198
rect 12002 3822 13626 5198
rect 13660 3822 15284 5198
rect 15318 3822 16942 5198
rect 16976 3822 18600 5198
rect 18634 3822 20258 5198
rect 20292 3822 21916 5198
rect 21950 3822 23574 5198
rect 23608 3822 25232 5198
rect 25266 3822 26890 5198
rect 26924 3822 28548 5198
rect 28582 3822 30206 5198
rect 30240 3822 31864 5198
rect 31898 3822 33522 5198
rect 33556 3822 33630 5198
rect -32980 3562 33630 3822
rect -32980 2186 -32798 3562
rect -32764 2186 -31140 3562
rect -31106 2186 -29482 3562
rect -29448 2186 -27824 3562
rect -27790 2186 -26166 3562
rect -26132 2186 -24508 3562
rect -24474 2186 -22850 3562
rect -22816 2186 -21192 3562
rect -21158 2186 -19534 3562
rect -19500 2186 -17876 3562
rect -17842 2186 -16218 3562
rect -16184 2186 -14560 3562
rect -14526 2186 -12902 3562
rect -12868 2186 -11244 3562
rect -11210 2186 -9586 3562
rect -9552 2186 -7928 3562
rect -7894 2186 -6270 3562
rect -6236 2186 -4612 3562
rect -4578 2186 -2954 3562
rect -2920 2186 -1296 3562
rect -1262 2186 362 3562
rect 396 2186 2020 3562
rect 2054 2186 3678 3562
rect 3712 2186 5336 3562
rect 5370 2186 6994 3562
rect 7028 2186 8652 3562
rect 8686 2186 10310 3562
rect 10344 2186 11968 3562
rect 12002 2186 13626 3562
rect 13660 2186 15284 3562
rect 15318 2186 16942 3562
rect 16976 2186 18600 3562
rect 18634 2186 20258 3562
rect 20292 2186 21916 3562
rect 21950 2186 23574 3562
rect 23608 2186 25232 3562
rect 25266 2186 26890 3562
rect 26924 2186 28548 3562
rect 28582 2186 30206 3562
rect 30240 2186 31864 3562
rect 31898 2186 33522 3562
rect 33556 2186 33630 3562
rect -32980 1926 33630 2186
rect -32980 634 -32798 1926
rect -32804 550 -32798 634
rect -32764 634 -31140 1926
rect -32764 550 -32758 634
rect -32804 538 -32758 550
rect -31146 550 -31140 634
rect -31106 634 -29482 1926
rect -31106 550 -31100 634
rect -31146 538 -31100 550
rect -29488 550 -29482 634
rect -29448 634 -27824 1926
rect -29448 550 -29442 634
rect -29488 538 -29442 550
rect -27830 550 -27824 634
rect -27790 634 -26166 1926
rect -27790 550 -27784 634
rect -27830 538 -27784 550
rect -26172 550 -26166 634
rect -26132 634 -24508 1926
rect -26132 550 -26126 634
rect -26172 538 -26126 550
rect -24514 550 -24508 634
rect -24474 634 -22850 1926
rect -24474 550 -24468 634
rect -24514 538 -24468 550
rect -22856 550 -22850 634
rect -22816 634 -21192 1926
rect -22816 550 -22810 634
rect -22856 538 -22810 550
rect -21198 550 -21192 634
rect -21158 634 -19534 1926
rect -21158 550 -21152 634
rect -21198 538 -21152 550
rect -19540 550 -19534 634
rect -19500 634 -17876 1926
rect -19500 550 -19494 634
rect -19540 538 -19494 550
rect -17882 550 -17876 634
rect -17842 634 -16218 1926
rect -17842 550 -17836 634
rect -17882 538 -17836 550
rect -16224 550 -16218 634
rect -16184 634 -14560 1926
rect -16184 550 -16178 634
rect -16224 538 -16178 550
rect -14566 550 -14560 634
rect -14526 634 -12902 1926
rect -14526 550 -14520 634
rect -14566 538 -14520 550
rect -12908 550 -12902 634
rect -12868 634 -11244 1926
rect -12868 550 -12862 634
rect -12908 538 -12862 550
rect -11250 550 -11244 634
rect -11210 634 -9586 1926
rect -11210 550 -11204 634
rect -11250 538 -11204 550
rect -9592 550 -9586 634
rect -9552 634 -7928 1926
rect -9552 550 -9546 634
rect -9592 538 -9546 550
rect -7934 550 -7928 634
rect -7894 634 -6270 1926
rect -7894 550 -7888 634
rect -7934 538 -7888 550
rect -6276 550 -6270 634
rect -6236 634 -4612 1926
rect -6236 550 -6230 634
rect -6276 538 -6230 550
rect -4618 550 -4612 634
rect -4578 634 -2954 1926
rect -4578 550 -4572 634
rect -4618 538 -4572 550
rect -2960 550 -2954 634
rect -2920 634 -1296 1926
rect -2920 550 -2914 634
rect -2960 538 -2914 550
rect -1302 550 -1296 634
rect -1262 634 362 1926
rect -1262 550 -1256 634
rect -1302 538 -1256 550
rect 356 550 362 634
rect 396 634 2020 1926
rect 396 550 402 634
rect 356 538 402 550
rect 2014 550 2020 634
rect 2054 634 3678 1926
rect 2054 550 2060 634
rect 2014 538 2060 550
rect 3672 550 3678 634
rect 3712 634 5336 1926
rect 3712 550 3718 634
rect 3672 538 3718 550
rect 5330 550 5336 634
rect 5370 634 6994 1926
rect 5370 550 5376 634
rect 5330 538 5376 550
rect 6988 550 6994 634
rect 7028 634 8652 1926
rect 7028 550 7034 634
rect 6988 538 7034 550
rect 8646 550 8652 634
rect 8686 634 10310 1926
rect 8686 550 8692 634
rect 8646 538 8692 550
rect 10304 550 10310 634
rect 10344 634 11968 1926
rect 10344 550 10350 634
rect 10304 538 10350 550
rect 11962 550 11968 634
rect 12002 634 13626 1926
rect 12002 550 12008 634
rect 11962 538 12008 550
rect 13620 550 13626 634
rect 13660 634 15284 1926
rect 13660 550 13666 634
rect 13620 538 13666 550
rect 15278 550 15284 634
rect 15318 634 16942 1926
rect 15318 550 15324 634
rect 15278 538 15324 550
rect 16936 550 16942 634
rect 16976 634 18600 1926
rect 16976 550 16982 634
rect 16936 538 16982 550
rect 18594 550 18600 634
rect 18634 634 20258 1926
rect 18634 550 18640 634
rect 18594 538 18640 550
rect 20252 550 20258 634
rect 20292 634 21916 1926
rect 20292 550 20298 634
rect 20252 538 20298 550
rect 21910 550 21916 634
rect 21950 634 23574 1926
rect 21950 550 21956 634
rect 21910 538 21956 550
rect 23568 550 23574 634
rect 23608 634 25232 1926
rect 23608 550 23614 634
rect 23568 538 23614 550
rect 25226 550 25232 634
rect 25266 634 26890 1926
rect 25266 550 25272 634
rect 25226 538 25272 550
rect 26884 550 26890 634
rect 26924 634 28548 1926
rect 26924 550 26930 634
rect 26884 538 26930 550
rect 28542 550 28548 634
rect 28582 634 30206 1926
rect 28582 550 28588 634
rect 28542 538 28588 550
rect 30200 550 30206 634
rect 30240 634 31864 1926
rect 30240 550 30246 634
rect 30200 538 30246 550
rect 31858 550 31864 634
rect 31898 634 33522 1926
rect 31898 550 31904 634
rect 31858 538 31904 550
rect 33516 550 33522 634
rect 33556 634 33630 1926
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 33976 13946 35004 15480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 33976 3946 35004 5480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect 33556 550 33562 634
rect 33516 538 33562 550
rect 788 470 848 486
rect 788 460 802 470
rect 614 436 802 460
rect 836 436 848 470
rect 614 424 848 436
rect 614 398 674 424
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect 612 256 674 398
rect 326 236 674 256
rect 326 216 676 236
rect 328 212 676 216
rect 328 184 358 212
rect 574 204 676 212
rect 326 182 358 184
rect -114 136 158 166
rect -114 124 -38 136
rect -34586 -54 -734 116
rect -114 90 -94 124
rect -60 90 -38 124
rect 130 96 158 136
rect 326 96 356 182
rect 34 94 80 96
rect -114 70 -38 90
rect -6 84 80 94
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -92 -486 -42 70
rect -6 -72 40 84
rect -6 -124 22 -72
rect -6 -292 40 -124
rect 74 -292 80 84
rect -6 -304 80 -292
rect 130 84 176 96
rect 130 -292 136 84
rect 170 -292 176 84
rect 130 -304 176 -292
rect 226 84 272 96
rect 226 -292 232 84
rect 266 -292 272 84
rect 226 -304 272 -292
rect 322 84 368 96
rect 322 -292 328 84
rect 362 -292 368 84
rect 322 -304 368 -292
rect 418 84 514 96
rect 418 -292 424 84
rect 458 -76 514 84
rect 492 -128 514 -76
rect 458 -292 514 -128
rect 418 -302 514 -292
rect 418 -304 494 -302
rect 30 -428 66 -304
rect 226 -426 262 -304
rect 30 -458 196 -428
rect 226 -454 420 -426
rect 226 -456 312 -454
rect 226 -458 272 -456
rect -92 -514 100 -486
rect -34586 -828 -734 -520
rect 72 -548 100 -514
rect 168 -548 196 -458
rect 384 -548 420 -454
rect -14 -552 32 -548
rect -48 -560 32 -552
rect -48 -610 -8 -560
rect -48 -706 -34 -610
rect -48 -736 -8 -706
rect 26 -736 32 -560
rect -48 -744 32 -736
rect -14 -748 32 -744
rect 72 -560 128 -548
rect 72 -736 88 -560
rect 122 -736 128 -560
rect 72 -748 128 -736
rect 168 -560 224 -548
rect 168 -736 184 -560
rect 218 -736 224 -560
rect 168 -744 224 -736
rect 178 -748 224 -744
rect 274 -560 320 -548
rect 274 -736 280 -560
rect 314 -734 320 -560
rect 370 -552 420 -548
rect 370 -560 452 -552
rect 314 -736 326 -734
rect 274 -748 326 -736
rect 370 -736 376 -560
rect 410 -610 452 -560
rect 436 -696 452 -610
rect 410 -736 452 -696
rect 370 -742 452 -736
rect 370 -748 416 -742
rect 286 -820 326 -748
rect 614 -816 676 204
rect 33976 52 35004 1480
rect 1532 -54 35054 52
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
rect 610 -818 678 -816
rect 576 -820 678 -818
rect 286 -866 678 -820
rect 576 -870 678 -866
rect 576 -872 616 -870
rect -86 -916 518 -900
rect -86 -968 -54 -916
rect 4 -968 346 -916
rect 404 -968 518 -916
rect -86 -982 518 -968
<< via1 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect 34166 15480 34698 15946
rect 34166 13480 34698 13946
rect 34166 11480 34698 11946
rect 34166 9480 34698 9946
rect 34166 7480 34698 7946
rect 34166 5480 34698 5946
rect 34166 3480 34698 3946
rect 34166 1480 34698 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 22 -124 40 -72
rect 40 -124 74 -72
rect 440 -128 458 -76
rect 458 -128 492 -76
rect -34 -706 -8 -610
rect -8 -706 22 -610
rect 384 -696 410 -610
rect 410 -696 436 -610
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
rect -54 -968 4 -916
rect 346 -968 404 -916
<< metal2 >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 33976 13946 35004 15480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 33976 3946 35004 5480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -6 -72 514 98
rect 33976 52 35004 1480
rect -6 -124 22 -72
rect 74 -76 514 -72
rect 74 -124 440 -76
rect -6 -128 440 -124
rect 492 -128 514 -76
rect -6 -304 514 -128
rect 1532 -54 35054 52
rect -34586 -828 -734 -520
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect -48 -610 452 -550
rect 1532 -570 35054 -520
rect -48 -706 -34 -610
rect 22 -696 384 -610
rect 436 -696 452 -610
rect 22 -706 452 -696
rect -48 -748 452 -706
rect -86 -912 518 -900
rect -86 -968 -54 -912
rect 4 -968 346 -912
rect 404 -968 518 -912
rect -86 -982 518 -968
<< via2 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect 34166 15480 34698 15946
rect 34166 13480 34698 13946
rect 34166 11480 34698 11946
rect 34166 9480 34698 9946
rect 34166 7480 34698 7946
rect 34166 5480 34698 5946
rect 34166 3480 34698 3946
rect 34166 1480 34698 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
rect -54 -916 4 -912
rect -54 -968 4 -916
rect 346 -916 404 -912
rect 346 -968 404 -916
<< metal3 >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 33976 13946 35004 15480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 33976 3946 35004 5480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect 33976 52 35004 1480
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
rect 1532 -54 35054 52
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
rect -86 -904 518 -900
rect -86 -968 -54 -904
rect 10 -968 346 -904
rect 410 -968 518 -904
rect -86 -982 518 -968
<< via3 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect 34166 15480 34698 15946
rect 34166 13480 34698 13946
rect 34166 11480 34698 11946
rect 34166 9480 34698 9946
rect 34166 7480 34698 7946
rect 34166 5480 34698 5946
rect 34166 3480 34698 3946
rect 34166 1480 34698 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
rect -54 -912 10 -904
rect -54 -968 4 -912
rect 4 -968 10 -912
rect 346 -912 410 -904
rect 346 -968 404 -912
rect 404 -968 410 -912
<< metal4 >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 388 -33510 1480
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 33976 13946 35004 15480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 33976 3946 35004 5480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect -34456 384 -33512 388
rect -34586 116 -33512 384
rect -34586 -54 -734 116
rect 33976 52 35004 1480
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
rect 1532 -54 35054 52
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
rect -86 -904 518 -900
rect -86 -968 -54 -904
rect 10 -968 346 -904
rect 410 -968 518 -904
rect -86 -982 518 -968
<< via4 >>
rect -34234 17480 -33702 17946
rect -32234 17480 -31702 17946
rect -30234 17480 -29702 17946
rect -28234 17480 -27702 17946
rect -26234 17480 -25702 17946
rect -24234 17480 -23702 17946
rect -22234 17480 -21702 17946
rect -20234 17480 -19702 17946
rect -18234 17480 -17702 17946
rect -16234 17480 -15702 17946
rect -14234 17480 -13702 17946
rect -12234 17480 -11702 17946
rect -10234 17480 -9702 17946
rect -8234 17480 -7702 17946
rect -6234 17480 -5702 17946
rect -4234 17480 -3702 17946
rect -2234 17480 -1702 17946
rect -234 17480 298 17946
rect 1766 17480 2298 17946
rect 3766 17480 4298 17946
rect 5766 17480 6298 17946
rect 7766 17480 8298 17946
rect 9766 17480 10298 17946
rect 11766 17480 12298 17946
rect 13766 17480 14298 17946
rect 15766 17480 16298 17946
rect 17766 17480 18298 17946
rect 19766 17480 20298 17946
rect 21766 17480 22298 17946
rect 23766 17480 24298 17946
rect 25766 17480 26298 17946
rect 27766 17480 28298 17946
rect 29766 17480 30298 17946
rect 31766 17480 32298 17946
rect 34166 17480 34698 17946
rect -34234 15480 -33702 15946
rect -34234 13480 -33702 13946
rect -34234 11480 -33702 11946
rect -34234 9480 -33702 9946
rect -34234 7480 -33702 7946
rect -34234 5480 -33702 5946
rect -34234 3480 -33702 3946
rect -34234 1480 -33702 1946
rect 34166 15480 34698 15946
rect 34166 13480 34698 13946
rect 34166 11480 34698 11946
rect 34166 9480 34698 9946
rect 34166 7480 34698 7946
rect 34166 5480 34698 5946
rect 34166 3480 34698 3946
rect 34166 1480 34698 1946
rect -33834 -520 -33302 -54
rect -31834 -520 -31302 -54
rect -29834 -520 -29302 -54
rect -27834 -520 -27302 -54
rect -25834 -520 -25302 -54
rect -23834 -520 -23302 -54
rect -21834 -520 -21302 -54
rect -19834 -520 -19302 -54
rect -17834 -520 -17302 -54
rect -15834 -520 -15302 -54
rect -13834 -520 -13302 -54
rect -11834 -520 -11302 -54
rect -9834 -520 -9302 -54
rect -7834 -520 -7302 -54
rect -5834 -520 -5302 -54
rect -3834 -520 -3302 -54
rect -1834 -520 -1302 -54
rect 2166 -520 2698 -54
rect 4166 -520 4698 -54
rect 6166 -520 6698 -54
rect 8166 -520 8698 -54
rect 10166 -520 10698 -54
rect 12166 -520 12698 -54
rect 14166 -520 14698 -54
rect 16166 -520 16698 -54
rect 18166 -520 18698 -54
rect 20166 -520 20698 -54
rect 22166 -520 22698 -54
rect 24166 -520 24698 -54
rect 26166 -520 26698 -54
rect 28166 -520 28698 -54
rect 30166 -520 30698 -54
rect 32166 -520 32698 -54
rect 34166 -520 34698 -54
<< metal5 >>
rect -34456 18152 -32822 18174
rect -34456 18112 34986 18152
rect -34456 17946 35004 18112
rect -34456 17480 -34234 17946
rect -33702 17480 -32234 17946
rect -31702 17480 -30234 17946
rect -29702 17480 -28234 17946
rect -27702 17480 -26234 17946
rect -25702 17480 -24234 17946
rect -23702 17480 -22234 17946
rect -21702 17480 -20234 17946
rect -19702 17480 -18234 17946
rect -17702 17480 -16234 17946
rect -15702 17480 -14234 17946
rect -13702 17480 -12234 17946
rect -11702 17480 -10234 17946
rect -9702 17480 -8234 17946
rect -7702 17480 -6234 17946
rect -5702 17480 -4234 17946
rect -3702 17480 -2234 17946
rect -1702 17480 -234 17946
rect 298 17480 1766 17946
rect 2298 17480 3766 17946
rect 4298 17480 5766 17946
rect 6298 17480 7766 17946
rect 8298 17480 9766 17946
rect 10298 17480 11766 17946
rect 12298 17480 13766 17946
rect 14298 17480 15766 17946
rect 16298 17480 17766 17946
rect 18298 17480 19766 17946
rect 20298 17480 21766 17946
rect 22298 17480 23766 17946
rect 24298 17480 25766 17946
rect 26298 17480 27766 17946
rect 28298 17480 29766 17946
rect 30298 17480 31766 17946
rect 32298 17480 34166 17946
rect 34698 17480 35004 17946
rect -34456 17406 35004 17480
rect -34456 17378 -32822 17406
rect -34456 17376 -33498 17378
rect -34456 15946 -33510 17376
rect -34456 15480 -34234 15946
rect -33702 15480 -33510 15946
rect -34456 13946 -33510 15480
rect -34456 13480 -34234 13946
rect -33702 13480 -33510 13946
rect -34456 11946 -33510 13480
rect -34456 11480 -34234 11946
rect -33702 11480 -33510 11946
rect -34456 9946 -33510 11480
rect -34456 9480 -34234 9946
rect -33702 9480 -33510 9946
rect -34456 7946 -33510 9480
rect -34456 7480 -34234 7946
rect -33702 7480 -33510 7946
rect -34456 5946 -33510 7480
rect -34456 5480 -34234 5946
rect -33702 5480 -33510 5946
rect -34456 3946 -33510 5480
rect -34456 3480 -34234 3946
rect -33702 3480 -33510 3946
rect -34456 1946 -33510 3480
rect -34456 1480 -34234 1946
rect -33702 1480 -33510 1946
rect -34456 384 -33510 1480
rect -34586 116 -33510 384
rect 33976 15946 35004 17406
rect 33976 15480 34166 15946
rect 34698 15480 35004 15946
rect 33976 13946 35004 15480
rect 33976 13480 34166 13946
rect 34698 13480 35004 13946
rect 33976 11946 35004 13480
rect 33976 11480 34166 11946
rect 34698 11480 35004 11946
rect 33976 9946 35004 11480
rect 33976 9480 34166 9946
rect 34698 9480 35004 9946
rect 33976 7946 35004 9480
rect 33976 7480 34166 7946
rect 34698 7480 35004 7946
rect 33976 5946 35004 7480
rect 33976 5480 34166 5946
rect 34698 5480 35004 5946
rect 33976 3946 35004 5480
rect 33976 3480 34166 3946
rect 34698 3480 35004 3946
rect 33976 1946 35004 3480
rect 33976 1480 34166 1946
rect 34698 1480 35004 1946
rect -34586 -54 -734 116
rect 33976 52 35004 1480
rect -34586 -520 -33834 -54
rect -33302 -520 -31834 -54
rect -31302 -520 -29834 -54
rect -29302 -520 -27834 -54
rect -27302 -520 -25834 -54
rect -25302 -520 -23834 -54
rect -23302 -520 -21834 -54
rect -21302 -520 -19834 -54
rect -19302 -520 -17834 -54
rect -17302 -520 -15834 -54
rect -15302 -520 -13834 -54
rect -13302 -520 -11834 -54
rect -11302 -520 -9834 -54
rect -9302 -520 -7834 -54
rect -7302 -520 -5834 -54
rect -5302 -520 -3834 -54
rect -3302 -520 -1834 -54
rect -1302 -520 -734 -54
rect -34586 -828 -734 -520
rect 1532 -54 35054 52
rect 1532 -520 2166 -54
rect 2698 -520 4166 -54
rect 4698 -520 6166 -54
rect 6698 -520 8166 -54
rect 8698 -520 10166 -54
rect 10698 -520 12166 -54
rect 12698 -520 14166 -54
rect 14698 -520 16166 -54
rect 16698 -520 18166 -54
rect 18698 -520 20166 -54
rect 20698 -520 22166 -54
rect 22698 -520 24166 -54
rect 24698 -520 26166 -54
rect 26698 -520 28166 -54
rect 28698 -520 30166 -54
rect 30698 -520 32166 -54
rect 32698 -520 34166 -54
rect 34698 -520 35054 -54
rect 1532 -570 35054 -520
<< labels >>
flabel locali 1074 346 1074 346 0 FreeSans 320 0 0 0 net2
flabel locali -424 370 -424 370 0 FreeSans 320 0 0 0 net1
flabel metal1 374 17216 374 17216 0 FreeSans 1600 0 0 0 VDD!
flabel metal1 60 -450 60 -450 0 FreeSans 320 0 0 0 in
flabel metal1 268 -436 268 -436 0 FreeSans 320 0 0 0 out
flabel locali 492 -496 492 -496 0 FreeSans 480 0 0 0 clkb_in
flabel locali -70 -794 -70 -794 0 FreeSans 480 0 0 0 cl_in
flabel metal4 178 -960 178 -952 0 FreeSans 1600 0 0 0 GND!
<< end >>
