* NGSPICE file created from 20bitCounter_flat.ext - technology: sky130A


* Top level circuit 20bitCounter_flat

X0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41487_21# a_41474_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20327_21# a_20314_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_9681_47# a_8491_47# a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22268_47# a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15617_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_32379_47# a_31933_47# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9747_21# a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30907_21# a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_24384_47# a_23469_47# a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_30167_47# a_29651_47# a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_19237_47# a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_805_47# a_761_289# a_639_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_38631_47# a_38115_47# a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5515_21# a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37255_21# a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_11219_47# a_10773_47# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28616_47# a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24081_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_19683_47# a_19237_47# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_16095_21# a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_17471_47# a_16955_47# a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3399_21# a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13979_21# a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35139_21# a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1283_21# a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 a_28791_21# a_28616_47# a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X43 a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1108_47# a_193_47# a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11863_21# a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X46 a_15005_47# a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33023_21# a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X48 a_9572_47# a_8657_47# a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X49 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 a_1283_21# a_1108_47# a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_17121_47# a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X53 a_38281_47# a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X54 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_4425_47# a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X56 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7631_21# a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39371_21# a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X58 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_37255_21# a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X59 a_36165_47# a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X60 a_2309_47# a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X61 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9269_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X62 a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X63 a_34049_47# a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X64 a_24384_47# a_23303_47# a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X65 a_41474_413# a_40397_47# a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X66 a_20314_413# a_19237_47# a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X67 a_30841_47# a_29651_47# a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X68 a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X69 a_26609_47# a_25419_47# a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X70 a_22268_47# a_21187_47# a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X71 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_11863_21# a_11797_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X72 a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X73 a_651_413# a_27_47# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_37255_21# a_37189_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X75 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 a_28616_47# a_27535_47# a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X77 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X78 a_35073_47# a_33883_47# a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X79 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X80 a_34617_289# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X81 a_26500_47# a_25419_47# a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X82 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_16095_21# a_16029_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X83 a_32545_47# a_32501_289# a_32379_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X84 a_13457_289# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X85 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11341_289# a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 a_38849_289# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X88 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32501_289# a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X89 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X90 a_11385_47# a_11341_289# a_11219_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X92 a_30732_47# a_29817_47# a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4993_289# a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X95 a_26675_21# a_26500_47# a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15573_289# a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36733_289# a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X99 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_2877_289# a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X101 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26197_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X102 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_18211_21# a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_19587_47# a_19071_47# a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X105 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13457_289# a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X107 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34617_289# a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9225_289# a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X111 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_805_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 a_28051_47# a_27535_47# a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X115 a_3399_21# a_3224_47# a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7109_289# a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17689_289# a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38849_289# a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X120 a_2755_47# a_2309_47# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X121 a_25585_47# a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X122 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X123 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_39371_21# a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X125 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30429_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X126 a_32391_413# a_31767_47# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_3399_21# a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X128 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X129 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_30275_413# a_29651_47# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X131 a_32957_47# a_31767_47# a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X132 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_26675_21# a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X133 a_2309_47# a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_36623_413# a_35999_47# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_13979_21# a_13913_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 a_11797_47# a_10607_47# a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X138 a_37189_47# a_35999_47# a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X139 a_34507_413# a_33883_47# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_22443_21# a_22377_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X141 a_9115_413# a_8491_47# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 a_13457_289# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X143 a_34617_289# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X144 a_20261_47# a_19071_47# a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X145 a_11341_289# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X146 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 a_7109_289# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_32848_47# a_31933_47# a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X149 a_24037_289# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X150 a_17689_289# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X151 a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24559_21# a_24546_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_11688_47# a_10773_47# a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X154 a_15573_289# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X155 a_41421_47# a_40231_47# a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X156 a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X157 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_7631_21# a_7565_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X159 a_25935_47# a_25419_47# a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X160 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11385_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X162 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X164 a_20152_47# a_19237_47# a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28791_21# a_28778_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 a_9225_289# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X167 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_28791_21# a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X168 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X169 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_16095_21# a_15920_47# a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_9225_289# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X173 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26675_21# a_26662_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X175 a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X176 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 a_15451_47# a_15005_47# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X178 a_31933_47# a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X179 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 a_7153_47# a_7109_289# a_6987_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X182 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X183 a_2659_47# a_2143_47# a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16095_21# a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X185 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 a_21703_47# a_21353_47# a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X188 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32545_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26500_47# a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X190 a_10773_47# a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 a_41312_47# a_40397_47# a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X192 a_10773_47# a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X193 a_36165_47# a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 a_40747_47# a_40397_47# a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 a_31933_47# a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X196 a_5340_47# a_4425_47# a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X197 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X198 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 a_37255_21# a_37080_47# a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X200 a_28051_47# a_27701_47# a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X201 a_6541_47# a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X202 a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41009_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X204 a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19849_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X207 a_2921_47# a_2877_289# a_2755_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_36611_47# a_36165_47# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X209 a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X210 a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X211 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X212 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_15005_47# a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X214 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 a_23819_47# a_23469_47# a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18211_21# a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X217 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_1283_21# a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 a_12889_47# a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X221 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_24559_21# a_24493_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 a_22377_47# a_21187_47# a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X223 a_22430_413# a_21353_47# a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 a_8657_47# a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X226 a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X227 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X228 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_33023_21# a_32957_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 a_19237_47# a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X230 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 a_30385_289# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X232 a_26662_413# a_25585_47# a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X233 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X234 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X235 a_19805_289# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X236 a_40965_289# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30732_47# a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X238 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X239 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X240 a_24546_413# a_23469_47# a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_9747_21# a_9681_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35139_21# a_35126_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 a_7565_47# a_6375_47# a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X245 a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X246 a_761_289# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X247 a_41009_47# a_40965_289# a_40843_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33023_21# a_33010_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X249 a_22268_47# a_21353_47# a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X250 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X251 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34964_47# a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X254 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X255 a_28778_413# a_27701_47# a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X256 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11688_47# a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32848_47# a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X259 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21965_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X260 a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X262 a_17567_47# a_17121_47# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X265 a_15355_47# a_14839_47# a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37255_21# a_37242_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X267 a_9269_47# a_9225_289# a_9103_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41487_21# a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X271 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_12889_47# a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26675_21# a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X274 a_26031_47# a_25585_47# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X275 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37080_47# a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X278 a_7456_47# a_6541_47# a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X281 a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24559_21# a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X283 a_21353_47# a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19805_289# a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_35139_21# a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X286 a_38727_47# a_38281_47# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X289 a_22443_21# a_22268_47# a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X290 a_36515_47# a_35999_47# a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X291 a_40397_47# a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22443_21# a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X293 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_13979_21# a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X295 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X297 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_30907_21# a_30841_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_3224_47# a_2143_47# a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X299 a_11231_413# a_10607_47# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X300 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2921_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 a_6541_47# a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X302 a_193_47# a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 a_4883_413# a_4259_47# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X304 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_35139_21# a_35073_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X305 a_34964_47# a_33883_47# a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X306 a_1108_47# a_27_47# a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 a_7631_21# a_7456_47# a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 a_32848_47# a_31767_47# a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X309 a_32501_289# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X310 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7153_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X311 a_15463_413# a_14839_47# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X312 a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X313 a_2767_413# a_2143_47# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X314 a_30732_47# a_29651_47# a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X315 a_11341_289# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X316 a_39196_47# a_38115_47# a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 a_18036_47# a_16955_47# a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 a_13347_413# a_12723_47# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X319 a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X320 a_5340_47# a_4259_47# a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 a_35126_413# a_34049_47# a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X322 a_19695_413# a_19071_47# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_6999_413# a_6375_47# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X324 a_37080_47# a_35999_47# a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X325 a_19805_289# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X326 a_17733_47# a_17689_289# a_17567_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X327 a_17579_413# a_16955_47# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 a_38739_413# a_38115_47# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X330 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40965_289# a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X333 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X334 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 a_30429_47# a_30385_289# a_30263_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X336 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 a_38893_47# a_38849_289# a_38727_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 a_40965_289# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X339 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X340 a_28147_47# a_27701_47# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X341 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26153_289# a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X343 a_11863_21# a_11688_47# a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X344 a_4993_289# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X345 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24037_289# a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X347 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X348 a_23469_47# a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X349 a_24559_21# a_24384_47# a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X350 a_543_47# a_27_47# a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X351 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_20327_21# a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X352 a_15920_47# a_15005_47# a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X353 a_23915_47# a_23469_47# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X354 a_21703_47# a_21187_47# a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X355 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28269_289# a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X357 a_33023_21# a_32848_47# a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X358 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_24559_21# a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X361 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X363 a_8657_47# a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X364 a_25935_47# a_25585_47# a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X365 a_9747_21# a_9572_47# a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X366 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_20327_21# a_20261_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X368 a_543_47# a_193_47# a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X369 a_6891_47# a_6375_47# a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X370 a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X371 a_21921_289# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X372 a_24037_289# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X373 a_19849_47# a_19805_289# a_19683_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_41487_21# a_41421_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X376 a_21921_289# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X377 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X378 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_5515_21# a_5449_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 a_3333_47# a_2143_47# a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3399_21# a_3386_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X381 a_28269_289# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X382 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X383 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X384 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_28791_21# a_28725_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X385 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13979_21# a_13966_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1283_21# a_1270_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X388 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X389 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X390 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X391 a_26153_289# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X392 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3224_47# a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_13979_21# a_13804_47# a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 a_7109_289# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7631_21# a_7618_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 a_13335_47# a_12889_47# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X398 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X399 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X401 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30907_21# a_30894_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9572_47# a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X405 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13804_47# a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X407 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1108_47# a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X410 a_5037_47# a_4993_289# a_4871_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39371_21# a_39358_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18211_21# a_18198_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5515_21# a_5502_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X414 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20327_21# a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X417 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7456_47# a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 a_28313_47# a_28269_289# a_28147_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X421 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16095_21# a_16082_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X423 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38893_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X424 a_34049_47# a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X425 a_23819_47# a_23303_47# a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X426 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X427 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X428 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X429 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39196_47# a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18036_47# a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5340_47# a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 a_35139_21# a_34964_47# a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X434 a_32283_47# a_31933_47# a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9747_21# a_9734_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X436 a_34495_47# a_34049_47# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X437 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_30907_21# a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X438 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17733_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X440 a_26500_47# a_25585_47# a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15920_47# a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X442 a_32283_47# a_31767_47# a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X443 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_9747_21# a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 a_30167_47# a_29817_47# a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X446 a_21353_47# a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X447 a_11123_47# a_10607_47# a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X448 a_36515_47# a_36165_47# a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X449 a_27701_47# a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X450 a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X452 a_9007_47# a_8491_47# a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X453 a_34399_47# a_34049_47# a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28791_21# a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X456 a_25585_47# a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X457 a_3224_47# a_2309_47# a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X458 a_1270_413# a_193_47# a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 a_33010_413# a_31933_47# a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X460 a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X461 a_193_47# a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X462 a_23469_47# a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X463 a_13804_47# a_12723_47# a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X464 a_30894_413# a_29817_47# a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X465 a_29817_47# a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X466 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X467 a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X468 a_11688_47# a_10607_47# a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X469 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_18211_21# a_18145_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X470 a_5502_413# a_4425_47# a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X471 a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X472 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X473 a_5449_47# a_4259_47# a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X474 a_7456_47# a_6375_47# a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X475 a_16082_413# a_15005_47# a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X476 a_37242_413# a_36165_47# a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X477 a_3386_413# a_2309_47# a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X478 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X479 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X480 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X482 a_15920_47# a_14839_47# a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X483 a_28725_47# a_27535_47# a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X484 a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X486 a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X487 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_39371_21# a_39305_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X489 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 a_7618_413# a_6541_47# a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X491 a_13239_47# a_12723_47# a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21921_289# a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X493 a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X494 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X495 a_36733_289# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X496 a_9572_47# a_8491_47# a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X497 a_39358_413# a_38281_47# a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X498 a_18198_413# a_17121_47# a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 a_34661_47# a_34617_289# a_34495_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X501 a_15573_289# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X502 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X504 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X505 a_41487_21# a_41312_47# a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_13501_47# a_13457_289# a_13335_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X507 a_40843_47# a_40397_47# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X508 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_33023_21# a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_761_289# a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X510 a_34399_47# a_33883_47# a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X511 a_28616_47# a_27701_47# a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X513 a_20327_21# a_20152_47# a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X515 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X516 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_11863_21# a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X518 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_41487_21# a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X519 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28313_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X520 a_37080_47# a_36165_47# a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X521 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X522 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X524 a_40397_47# a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X525 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X526 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 a_21811_413# a_21187_47# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X528 a_5515_21# a_5340_47# a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X529 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5037_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X530 a_27701_47# a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X531 a_4871_47# a_4425_47# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X532 a_40855_413# a_40231_47# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X533 a_18145_47# a_16955_47# a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X534 a_17689_289# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X535 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_5515_21# a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 a_9103_47# a_8657_47# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X537 a_26043_413# a_25419_47# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 a_23927_413# a_23303_47# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 a_41312_47# a_40231_47# a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X540 a_20152_47# a_19071_47# a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X541 a_4425_47# a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 a_13913_47# a_12723_47# a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X543 a_39305_47# a_38115_47# a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X544 a_28159_413# a_27535_47# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X545 a_36777_47# a_36733_289# a_36611_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X546 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X547 a_18036_47# a_17121_47# a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30385_289# a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X549 a_15617_47# a_15573_289# a_15451_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11863_21# a_11850_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X551 a_34964_47# a_34049_47# a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X552 a_26153_289# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X553 a_40747_47# a_40231_47# a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X554 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X555 a_639_47# a_193_47# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X556 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X557 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_1283_21# a_1217_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 a_24081_47# a_24037_289# a_23915_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X559 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X560 a_13804_47# a_12889_47# a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X561 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_21799_47# a_21353_47# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X563 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34661_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X564 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X565 a_39196_47# a_38281_47# a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X566 a_30907_21# a_30732_47# a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X567 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13501_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 a_39371_21# a_39196_47# a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X569 a_30263_47# a_29817_47# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X570 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_22443_21# a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_2877_289# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X575 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X576 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X577 a_18211_21# a_18036_47# a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X578 a_6891_47# a_6541_47# a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X579 a_11123_47# a_10773_47# a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X580 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X583 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X584 a_6987_47# a_6541_47# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X585 a_17471_47# a_17121_47# a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 a_38631_47# a_38281_47# a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X587 a_29817_47# a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X589 a_4775_47# a_4425_47# a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X590 a_4775_47# a_4259_47# a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X591 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X593 a_15355_47# a_15005_47# a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 a_2659_47# a_2309_47# a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X595 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_38281_47# a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_7631_21# a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X598 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 a_9007_47# a_8657_47# a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X600 a_13239_47# a_12889_47# a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X601 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X602 a_17121_47# a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X604 a_11850_413# a_10773_47# a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 a_19587_47# a_19237_47# a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 a_2877_289# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X607 a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X608 a_16029_47# a_14839_47# a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X609 a_761_289# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X610 a_32501_289# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X611 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X612 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_26675_21# a_26609_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X613 a_24493_47# a_23303_47# a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X614 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X615 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X616 a_30385_289# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20152_47# a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X618 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41312_47# a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X620 a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X621 a_13966_413# a_12889_47# a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 a_38849_289# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X623 a_21965_47# a_21921_289# a_21799_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_4993_289# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X625 a_9734_413# a_8657_47# a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X626 a_28269_289# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X627 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X628 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 a_36733_289# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22443_21# a_22430_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24384_47# a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_3399_21# a_3333_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X633 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X634 a_26197_47# a_26153_289# a_26031_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X635 a_1217_47# a_27_47# a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X636 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36777_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X638 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X639 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30732_47# 0.02fF
C1 a_36165_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C2 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6999_413# 0.17fF
C3 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.53fF
C4 a_30732_47# a_30841_47# 0.04fF
C5 a_30907_21# a_31086_47# 0.04fF
C6 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# 0.27fF
C7 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35703_47# 0.27fF
C8 a_2309_47# a_2877_289# 0.41fF
C9 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0.02fF
C10 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15463_413# 0.26fF
C11 a_32501_289# a_32283_47# 0.50fF
C12 a_31933_47# a_33023_21# 0.10fF
C13 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4259_47# 0.71fF
C14 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15573_289# 0.46fF
C15 a_36165_47# a_36515_47# 0.49fF
C16 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38281_47# 0.72fF
C17 a_34399_47# a_34049_47# 0.49fF
C18 a_32501_289# a_32188_47# 0.00fF
C19 a_31933_47# a_32391_413# 0.12fF
C20 a_33023_21# a_32848_47# 0.62fF
C21 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23007_47# 0.09fF
C22 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# 0.27fF
C23 a_9926_47# a_9747_21# 0.04fF
C24 a_9681_47# a_9572_47# 0.04fF
C25 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38739_413# 0.17fF
C26 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29817_47# 0.08fF
C27 a_32848_47# a_32391_413# 0.01fF
C28 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6796_47# 0.06fF
C29 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# 0.27fF
C30 a_8912_47# a_8491_47# 0.23fF
C31 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.24fF
C32 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26043_413# 0.17fF
C33 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[14]/D 1.68fF
C34 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15005_47# 1.17fF
C35 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15260_47# 0.15fF
C36 a_31933_47# a_32283_47# 0.49fF
C37 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37255_21# 0.22fF
C38 a_35999_47# a_37080_47# 0.27fF
C39 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[2]/D 1.68fF
C40 a_34964_47# a_33883_47# 0.27fF
C41 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.22fF
C42 a_32283_47# a_32848_47# 0.01fF
C43 a_31933_47# a_32188_47# 0.22fF
C44 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38631_47# 0.09fF
C45 a_38115_47# a_39371_21# 0.12fF
C46 a_5340_47# a_4883_413# 0.01fF
C47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22430_413# 0.01fF
C48 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5694_47# 0.01fF
C49 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22268_47# 0.68fF
C50 a_22622_47# a_22443_21# 0.04fF
C51 a_22377_47# a_22268_47# 0.04fF
C52 a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.63fF
C53 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8195_47# 0.09fF
C54 a_8657_47# a_8195_47# 0.01fF
C55 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25840_47# 0.06fF
C56 a_7618_413# a_7456_47# 0.04fF
C57 a_10773_47# a_11341_289# 0.41fF
C58 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_29651_47# 0.99fF
C59 a_31933_47# a_32501_289# 0.41fF
C60 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16659_47# 0.27fF
C61 a_448_47# a_651_413# 0.02fF
C62 a_40652_47# a_40965_289# 0.00fF
C63 a_40855_413# a_40397_47# 0.12fF
C64 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11850_413# 0.01fF
C65 a_37255_21# a_37434_47# 0.04fF
C66 a_37080_47# a_37189_47# 0.04fF
C67 a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C68 a_32501_289# a_32848_47# 0.13fF
C69 a_34964_47# a_35703_47# 0.00fF
C70 a_26662_413# a_26500_47# 0.04fF
C71 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.45fF
C72 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22443_21# 0.73fF
C73 a_34399_47# a_34507_413# 0.21fF
C74 a_27701_47# a_27239_47# 0.01fF
C75 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.27fF
C76 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.45fF
C77 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5449_47# 0.01fF
C78 a_32848_47# a_33587_47# 0.00fF
C79 a_31933_47# a_31471_47# 0.01fF
C80 a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.36fF
C81 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7456_47# 0.68fF
C82 a_30894_413# a_30732_47# 0.04fF
C83 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.11fF
C84 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.45fF
C85 a_2877_289# a_2767_413# 0.23fF
C86 a_6987_47# a_6891_47# 0.07fF
C87 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_27239_47# 0.09fF
C88 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.36fF
C89 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.27fF
C90 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15920_47# 0.39fF
C91 a_1108_47# a_1270_413# 0.04fF
C92 a_1847_47# a_2309_47# 0.01fF
C93 a_30732_47# a_31471_47# 0.00fF
C94 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.19fF
C95 a_38739_413# a_39196_47# 0.01fF
C96 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9926_47# 0.01fF
C97 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.12fF
C98 a_18775_47# a_19071_47# 0.07fF
C99 a_31933_47# a_32848_47# 0.29fF
C100 a_5340_47# a_6079_47# 0.00fF
C101 a_4775_47# a_4883_413# 0.21fF
C102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34399_47# 0.28fF
C103 a_26031_47# a_25935_47# 0.07fF
C104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_10607_47# 0.56fF
C105 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21703_47# 0.36fF
C106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_31767_47# 0.56fF
C107 a_30263_47# a_30167_47# 0.07fF
C108 a_19587_47# a_19683_47# 0.07fF
C109 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36733_289# 0.10fF
C110 a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.02fF
C111 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7631_21# 0.73fF
C112 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28159_413# 0.01fF
C113 a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.10fF
C114 a_38115_47# a_38849_289# 0.16fF
C115 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38281_47# 0.65fF
C116 a_2877_289# a_2564_47# 0.00fF
C117 a_2309_47# a_2767_413# 0.12fF
C118 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26500_47# 0.68fF
C119 a_24559_21# a_24738_47# 0.04fF
C120 a_24384_47# a_24493_47# 0.04fF
C121 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.11fF
C122 a_30907_21# a_31471_47# 0.30fF
C123 a_1108_47# a_651_413# 0.01fF
C124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16095_21# 0.37fF
C125 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[6]/D 1.68fF
C126 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17733_47# 0.01fF
C127 a_13804_47# a_13966_413# 0.04fF
C128 a_4993_289# a_4883_413# 0.23fF
C129 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21921_289# 0.46fF
C130 a_4775_47# a_4680_47# 0.13fF
C131 a_5515_21# a_6079_47# 0.30fF
C132 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21811_413# 0.26fF
C133 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.27fF
C134 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6891_47# 0.36fF
C135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.19fF
C136 a_20891_47# a_21353_47# 0.01fF
C137 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_27956_47# 0.53fF
C138 a_2309_47# a_2564_47# 0.22fF
C139 a_41312_47# a_41474_413# 0.04fF
C140 a_34617_289# a_34304_47# 0.00fF
C141 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26675_21# 0.73fF
C142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15355_47# 0.28fF
C143 a_30907_21# a_30732_47# 0.62fF
C144 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39550_47# 0.01fF
C145 a_38727_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.02fF
C146 a_35703_47# a_35999_47# 0.07fF
C147 a_18211_21# a_19071_47# 0.02fF
C148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.19fF
C149 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11231_413# 0.17fF
C150 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17567_47# 0.02fF
C151 a_13239_47# a_13335_47# 0.07fF
C152 a_13144_47# a_13347_413# 0.02fF
C153 a_4993_289# a_4680_47# 0.00fF
C154 a_5515_21# a_5340_47# 0.62fF
C155 a_4425_47# a_4883_413# 0.12fF
C156 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21353_47# 1.17fF
C157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21608_47# 0.15fF
C158 a_37080_47# a_37242_413# 0.04fF
C159 a_30275_413# a_30732_47# 0.01fF
C160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6999_413# 0.26fF
C161 a_41487_21# a_40965_289# 0.03fF
C162 a_41312_47# a_40397_47# 0.29fF
C163 a_41009_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C164 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7109_289# 0.46fF
C165 a_27535_47# a_27956_47# 0.23fF
C166 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# 0.24fF
C167 a_2877_289# a_3224_47# 0.13fF
C168 a_1108_47# a_1217_47# 0.04fF
C169 a_40747_47# a_40843_47# 0.07fF
C170 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25935_47# 0.36fF
C171 a_34399_47# a_34964_47# 0.01fF
C172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15573_289# 0.29fF
C173 a_1108_47# a_1847_47# 0.00fF
C174 a_30167_47# a_30732_47# 0.01fF
C175 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C176 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11028_47# 0.06fF
C177 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C178 a_4775_47# a_5340_47# 0.01fF
C179 a_4425_47# a_4680_47# 0.22fF
C180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23007_47# 0.27fF
C181 a_36515_47# a_36611_47# 0.07fF
C182 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38739_413# 0.26fF
C184 a_3224_47# a_3386_413# 0.04fF
C185 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6541_47# 1.17fF
C186 a_38536_47# a_38631_47# 0.13fF
C187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6796_47# 0.15fF
C188 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28616_47# 0.05fF
C189 a_2877_289# a_3399_21# 0.03fF
C190 a_2309_47# a_3224_47# 0.29fF
C191 a_10311_47# a_10773_47# 0.01fF
C192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26043_413# 0.26fF
C193 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26153_289# 0.46fF
C194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.45fF
C195 a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.36fF
C196 a_30385_289# a_30732_47# 0.13fF
C197 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.71fF
C198 a_30167_47# a_30907_21# 0.02fF
C199 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[10]/D 1.68fF
C200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15005_47# 0.72fF
C201 a_22377_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.45fF
C203 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19237_47# 0.08fF
C204 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12427_47# 0.09fF
C205 a_20891_47# a_21187_47# 0.07fF
C206 a_13804_47# a_13347_413# 0.01fF
C207 a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.71fF
C208 a_4993_289# a_5340_47# 0.13fF
C209 a_4775_47# a_5515_21# 0.02fF
C210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22268_47# 0.39fF
C211 a_2659_47# a_2755_47# 0.07fF
C212 a_2564_47# a_2767_413# 0.02fF
C213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_8195_47# 0.27fF
C214 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40855_413# 0.17fF
C215 a_30275_413# a_30167_47# 0.21fF
C216 a_19587_47# a_19695_413# 0.21fF
C217 a_27535_47# a_28616_47# 0.27fF
C218 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28791_21# 0.22fF
C219 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.11fF
C220 a_2877_289# a_2659_47# 0.50fF
C221 a_2309_47# a_3399_21# 0.10fF
C222 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_27535_47# 0.02fF
C223 a_8912_47# a_9115_413# 0.02fF
C224 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25585_47# 1.17fF
C225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_25840_47# 0.15fF
C226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_29651_47# 0.56fF
C227 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21187_47# 0.99fF
C228 a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.02fF
C229 a_29817_47# a_30732_47# 0.29fF
C230 a_30385_289# a_30907_21# 0.03fF
C231 a_30072_47# a_30275_413# 0.02fF
C232 a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.71fF
C233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11850_413# 0.01fF
C234 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11688_47# 0.68fF
C235 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9572_47# 0.05fF
C236 a_4993_289# a_5515_21# 0.03fF
C237 a_4425_47# a_5340_47# 0.29fF
C238 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.11fF
C239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22443_21# 0.37fF
C240 a_34617_289# a_35139_21# 0.03fF
C241 a_23469_47# a_23007_47# 0.01fF
C242 a_19587_47# a_19492_47# 0.13fF
C243 a_30072_47# a_30167_47# 0.13fF
C244 a_30275_413# a_30385_289# 0.23fF
C245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7456_47# 0.39fF
C246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.19fF
C247 a_19805_289# a_19695_413# 0.23fF
C248 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28051_47# 0.09fF
C249 a_27535_47# a_28791_21# 0.12fF
C250 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.36fF
C251 a_2309_47# a_2659_47# 0.49fF
C252 a_543_47# a_1283_21# 0.02fF
C253 a_40231_47# a_40965_289# 0.16fF
C254 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40397_47# 0.65fF
C255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_27239_47# 0.27fF
C256 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.27fF
C257 a_30385_289# a_30167_47# 0.50fF
C258 a_29817_47# a_30907_21# 0.10fF
C259 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C260 a_38536_47# a_38281_47# 0.22fF
C261 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11863_21# 0.73fF
C262 a_8491_47# a_9572_47# 0.27fF
C263 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9747_21# 0.22fF
C264 a_13804_47# a_14543_47# 0.00fF
C265 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37189_47# 0.01fF
C266 a_20327_21# a_21187_47# 0.02fF
C267 a_13239_47# a_13347_413# 0.21fF
C268 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17579_413# 0.01fF
C269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21703_47# 0.28fF
C270 a_4993_289# a_4775_47# 0.50fF
C271 a_4425_47# a_5515_21# 0.10fF
C272 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_8491_47# 0.02fF
C273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7631_21# 0.37fF
C274 a_3224_47# a_2767_413# 0.01fF
C275 a_30072_47# a_30385_289# 0.00fF
C276 a_30275_413# a_29817_47# 0.12fF
C277 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.11fF
C278 a_19237_47# a_19695_413# 0.12fF
C279 a_19805_289# a_19492_47# 0.00fF
C280 a_27535_47# a_28051_47# 0.42fF
C281 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28269_289# 0.10fF
C282 a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.02fF
C283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26500_47# 0.39fF
C284 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36777_47# 0.01fF
C285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.19fF
C286 a_29817_47# a_30167_47# 0.49fF
C287 a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.71fF
C288 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15463_413# 0.01fF
C289 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.45fF
C291 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11123_47# 0.36fF
C292 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17376_47# 0.53fF
C293 a_13239_47# a_13144_47# 0.13fF
C294 a_13457_289# a_13347_413# 0.23fF
C295 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9007_47# 0.09fF
C296 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19587_47# 0.36fF
C297 a_8491_47# a_9747_21# 0.12fF
C298 a_13979_21# a_14543_47# 0.30fF
C299 a_4425_47# a_4775_47# 0.49fF
C300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21921_289# 0.29fF
C301 a_19587_47# a_20152_47# 0.01fF
C302 a_19237_47# a_19492_47# 0.22fF
C303 a_30072_47# a_29817_47# 0.22fF
C304 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9572_47# 0.02fF
C305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6891_47# 0.28fF
C306 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_27701_47# 0.65fF
C307 a_27535_47# a_28269_289# 0.16fF
C308 a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.27fF
C309 a_41312_47# a_42051_47# 0.00fF
C310 a_40747_47# a_40855_413# 0.21fF
C311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26675_21# 0.37fF
C312 a_25123_47# a_25585_47# 0.01fF
C313 a_29817_47# a_30385_289# 0.41fF
C314 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3578_47# 0.01fF
C315 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15260_47# 0.53fF
C316 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41312_47# 0.68fF
C317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11231_413# 0.26fF
C318 a_13979_21# a_13804_47# 0.62fF
C319 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.68fF
C320 a_13457_289# a_13144_47# 0.00fF
C321 a_12889_47# a_13347_413# 0.12fF
C322 a_16955_47# a_17376_47# 0.23fF
C323 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9225_289# 0.10fF
C324 a_8491_47# a_9007_47# 0.42fF
C325 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19805_289# 0.46fF
C326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21353_47# 0.72fF
C327 a_4425_47# a_4993_289# 0.41fF
C328 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18198_413# 0.01fF
C329 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# 0.27fF
C330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7109_289# 0.29fF
C331 a_3224_47# a_3963_47# 0.00fF
C332 a_2659_47# a_2767_413# 0.21fF
C333 a_19805_289# a_20152_47# 0.13fF
C334 a_19587_47# a_20327_21# 0.02fF
C335 a_27535_47# a_27701_47# 1.60fF
C336 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38536_47# 0.01fF
C337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_25935_47# 0.28fF
C338 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[4]/D 1.68fF
C339 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3333_47# 0.01fF
C340 a_14839_47# a_15260_47# 0.23fF
C341 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# 0.24fF
C342 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37819_47# 0.09fF
C343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11028_47# 0.15fF
C344 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.99fF
C345 a_12889_47# a_13144_47# 0.22fF
C346 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_8657_47# 0.65fF
C347 a_8491_47# a_9225_289# 0.16fF
C348 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19237_47# 1.17fF
C349 a_13239_47# a_13804_47# 0.01fF
C350 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16274_47# 0.01fF
C351 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33010_413# 0.01fF
C352 a_2659_47# a_2564_47# 0.13fF
C353 a_3399_21# a_3963_47# 0.30fF
C354 a_19805_289# a_20327_21# 0.03fF
C355 a_19237_47# a_20152_47# 0.29fF
C356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6541_47# 0.72fF
C357 a_16659_47# a_17121_47# 0.01fF
C358 a_15920_47# a_16082_413# 0.04fF
C359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26153_289# 0.29fF
C360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.45fF
C361 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5502_413# 0.01fF
C362 a_37080_47# a_36623_413# 0.01fF
C363 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15920_47# 0.05fF
C364 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8491_47# 0.99fF
C365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_12427_47# 0.27fF
C366 a_8491_47# a_8657_47# 1.60fF
C367 a_13457_289# a_13804_47# 0.13fF
C368 a_13239_47# a_13979_21# 0.02fF
C369 a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.36fF
C370 a_35073_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C371 a_9734_413# a_9572_47# 0.04fF
C372 a_3399_21# a_3224_47# 0.62fF
C373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40855_413# 0.26fF
C374 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31086_47# 0.01fF
C375 a_19237_47# a_20327_21# 0.10fF
C376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.19fF
C377 a_15355_47# a_15451_47# 0.07fF
C378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_25585_47# 0.72fF
C379 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39371_21# 0.73fF
C380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21187_47# 0.56fF
C381 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3578_47# 0.01fF
C382 a_14839_47# a_15920_47# 0.27fF
C383 a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.21fF
C384 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16095_21# 0.22fF
C385 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_14839_47# 0.02fF
C386 a_40652_47# a_40231_47# 0.23fF
C387 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4680_47# 0.01fF
C388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11688_47# 0.39fF
C389 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.11fF
C390 a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.02fF
C391 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[19]/D 1.30fF
C392 a_13457_289# a_13979_21# 0.03fF
C393 a_12889_47# a_13804_47# 0.29fF
C394 a_40747_47# a_41312_47# 0.01fF
C395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.19fF
C396 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.11fF
C397 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17579_413# 0.17fF
C398 a_2659_47# a_3224_47# 0.01fF
C399 a_9103_47# a_9007_47# 0.07fF
C400 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C401 a_28791_21# a_28970_47# 0.04fF
C402 a_28616_47# a_28725_47# 0.04fF
C403 a_23469_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C404 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[16]/D 1.68fF
C405 a_14839_47# a_16095_21# 0.12fF
C406 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15355_47# 0.09fF
C407 a_34495_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.02fF
C408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11863_21# 0.37fF
C409 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C410 a_13457_289# a_13239_47# 0.50fF
C411 a_12889_47# a_13979_21# 0.10fF
C412 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.27fF
C413 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17376_47# 0.06fF
C414 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33023_21# 0.73fF
C415 a_38536_47# a_38739_413# 0.02fF
C416 a_2659_47# a_3399_21# 0.02fF
C417 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36515_47# 0.36fF
C418 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32391_413# 0.17fF
C419 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# 0.63fF
C420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.19fF
C421 a_4680_47# a_4259_47# 0.23fF
C422 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C423 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13966_413# 0.01fF
C424 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4883_413# 0.17fF
C425 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15573_289# 0.10fF
C426 a_14839_47# a_15355_47# 0.42fF
C427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11123_47# 0.28fF
C428 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34304_47# 0.06fF
C429 a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.02fF
C430 a_12889_47# a_13239_47# 0.49fF
C431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19587_47# 0.28fF
C432 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32283_47# 0.36fF
C433 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38849_289# 0.46fF
C434 a_37255_21# a_37819_47# 0.30fF
C435 a_36515_47# a_36420_47# 0.13fF
C436 a_9115_413# a_9572_47# 0.01fF
C437 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32188_47# 0.06fF
C438 a_39371_21# a_39196_47# 0.62fF
C439 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23915_47# 0.02fF
C440 a_40231_47# a_39935_47# 0.07fF
C441 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12042_47# 0.01fF
C442 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4680_47# 0.06fF
C443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41312_47# 0.39fF
C444 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15005_47# 0.65fF
C445 a_14839_47# a_15573_289# 0.16fF
C446 a_29355_47# a_29817_47# 0.01fF
C447 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.45fF
C448 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11341_289# 0.46fF
C449 a_12889_47# a_13457_289# 0.41fF
C450 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9734_413# 0.01fF
C451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18198_413# 0.01fF
C452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19805_289# 0.29fF
C453 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32501_289# 0.46fF
C454 a_28616_47# a_28778_413# 0.04fF
C455 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30894_413# 0.01fF
C456 a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.09fF
C457 a_41487_21# a_40231_47# 0.12fF
C458 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33587_47# 0.09fF
C459 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31471_47# 0.09fF
C460 a_33023_21# a_33202_47# 0.04fF
C461 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34049_47# 0.65fF
C462 a_5340_47# a_4259_47# 0.27fF
C463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.45fF
C464 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6079_47# 0.09fF
C465 a_14839_47# a_15005_47# 1.60fF
C466 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36165_47# 1.17fF
C467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37819_47# 0.27fF
C468 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10773_47# 1.17fF
C469 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.56fF
C470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19237_47# 0.72fF
C471 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7810_47# 0.01fF
C472 a_28051_47# a_28147_47# 0.07fF
C473 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31933_47# 1.17fF
C474 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_12723_47# 0.02fF
C475 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28970_47# 0.01fF
C476 a_9115_413# a_9007_47# 0.21fF
C477 a_10311_47# a_9572_47# 0.00fF
C478 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32848_47# 0.68fF
C479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33010_413# 0.01fF
C480 a_2143_47# a_1283_21# 0.02fF
C481 a_5515_21# a_4259_47# 0.12fF
C482 a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.71fF
C483 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.11fF
C484 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30732_47# 0.68fF
C485 a_36165_47# a_36420_47# 0.22fF
C486 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5340_47# 0.68fF
C487 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13347_413# 0.17fF
C488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5502_413# 0.01fF
C489 a_34304_47# a_34049_47# 0.22fF
C490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_8491_47# 0.56fF
C491 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35999_47# 0.02fF
C492 a_38849_289# a_39196_47# 0.13fF
C493 a_8912_47# a_9007_47# 0.13fF
C494 a_9115_413# a_9225_289# 0.23fF
C495 a_10311_47# a_9747_21# 0.30fF
C496 a_27956_47# a_28159_413# 0.02fF
C497 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35139_21# 0.73fF
C498 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[11]/D 1.68fF
C499 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30907_21# 0.73fF
C500 a_4775_47# a_4259_47# 0.42fF
C501 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13144_47# 0.06fF
C502 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36623_413# 0.01fF
C503 a_36515_47# a_37255_21# 0.02fF
C504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39371_21# 0.37fF
C505 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5515_21# 0.73fF
C506 a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C507 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4425_47# 0.08fF
C508 a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.36fF
C509 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.08fF
C510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.37fF
C511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.19fF
C512 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9115_413# 0.17fF
C513 a_5515_21# a_5694_47# 0.04fF
C514 a_5340_47# a_5449_47# 0.04fF
C515 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39358_413# 0.01fF
C516 a_33587_47# a_34049_47# 0.01fF
C517 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30275_413# 0.17fF
C518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.19fF
C519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17579_413# 0.26fF
C520 a_8912_47# a_9225_289# 0.00fF
C521 a_9115_413# a_8657_47# 0.12fF
C522 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# 0.27fF
C523 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_1283_21# 0.71fF
C524 a_4993_289# a_4259_47# 0.16fF
C525 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23303_47# 0.99fF
C526 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30167_47# 0.36fF
C527 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23927_413# 0.01fF
C528 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14158_47# 0.01fF
C529 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14543_47# 0.09fF
C530 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38115_47# 0.99fF
C531 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4775_47# 0.36fF
C532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.45fF
C533 a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.02fF
C534 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# 0.63fF
C535 a_34304_47# a_34507_413# 0.02fF
C536 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8912_47# 0.06fF
C537 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6999_413# 0.01fF
C538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33023_21# 0.37fF
C539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17376_47# 0.15fF
C540 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30072_47# 0.06fF
C541 a_8912_47# a_8657_47# 0.22fF
C542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32391_413# 0.26fF
C543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36515_47# 0.28fF
C544 a_28616_47# a_28159_413# 0.01fF
C545 a_761_289# a_1283_21# 0.03fF
C546 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_543_47# 0.30fF
C547 a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C548 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30385_289# 0.46fF
C549 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23724_47# 0.53fF
C550 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28778_413# 0.01fF
C551 a_4425_47# a_4259_47# 1.60fF
C552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13966_413# 0.01fF
C553 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13804_47# 0.68fF
C554 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4883_413# 0.26fF
C555 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4993_289# 0.46fF
C556 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.27fF
C557 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34617_289# 0.46fF
C558 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6796_47# 0.53fF
C559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34304_47# 0.15fF
C560 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10311_47# 0.09fF
C561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32283_47# 0.28fF
C562 a_36165_47# a_37255_21# 0.10fF
C563 a_36733_289# a_36515_47# 0.50fF
C564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38849_289# 0.29fF
C565 a_35139_21# a_34049_47# 0.10fF
C566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32188_47# 0.15fF
C567 a_38281_47# a_38631_47# 0.49fF
C568 a_193_47# a_1283_21# 0.10fF
C569 a_761_289# a_543_47# 0.50fF
C570 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C571 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26854_47# 0.01fF
C572 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_29817_47# 1.17fF
C573 a_23303_47# a_23724_47# 0.23fF
C574 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# 0.24fF
C575 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13979_21# 0.73fF
C576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4680_47# 0.15fF
C577 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4425_47# 1.17fF
C578 a_39358_413# a_39196_47# 0.04fF
C579 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9734_413# 0.01fF
C580 a_6375_47# a_6796_47# 0.23fF
C581 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# 0.24fF
C582 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11341_289# 0.29fF
C583 a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.71fF
C584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32501_289# 0.29fF
C585 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30894_413# 0.01fF
C586 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37080_47# 0.05fF
C587 a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.05fF
C588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33587_47# 0.27fF
C589 a_28616_47# a_29355_47# 0.00fF
C590 a_28051_47# a_28159_413# 0.21fF
C591 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39371_21# 0.22fF
C592 a_38115_47# a_39196_47# 0.27fF
C593 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1283_21# 0.22fF
C594 a_193_47# a_543_47# 0.49fF
C595 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18390_47# 0.01fF
C596 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# 0.63fF
C597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_31471_47# 0.27fF
C598 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20506_47# 0.01fF
C599 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26043_413# 0.01fF
C600 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24384_47# 0.05fF
C601 a_38727_47# a_38631_47# 0.07fF
C602 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13239_47# 0.36fF
C603 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6079_47# 0.27fF
C605 a_18775_47# a_19237_47# 0.01fF
C606 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36165_47# 0.72fF
C607 a_18036_47# a_18198_413# 0.04fF
C608 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.36fF
C609 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7456_47# 0.05fF
C610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_10773_47# 0.72fF
C611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_31933_47# 0.72fF
C612 a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.71fF
C613 a_40855_413# a_40965_289# 0.23fF
C614 a_28791_21# a_29355_47# 0.30fF
C615 a_28051_47# a_27956_47# 0.13fF
C616 a_28269_289# a_28159_413# 0.23fF
C617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32848_47# 0.39fF
C618 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_543_47# 0.09fF
C619 a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.02fF
C620 a_27_47# a_1283_21# 0.12fF
C621 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20261_47# 0.01fF
C622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30732_47# 0.39fF
C623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.19fF
C624 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18145_47# 0.01fF
C625 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.11fF
C626 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_25840_47# 0.53fF
C627 a_23303_47# a_24384_47# 0.27fF
C628 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24559_21# 0.22fF
C629 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_3963_47# 0.01fF
C630 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13457_289# 0.46fF
C631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5340_47# 0.39fF
C632 a_36165_47# a_36733_289# 0.41fF
C633 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13347_413# 0.26fF
C634 a_34617_289# a_34049_47# 0.41fF
C635 a_17471_47# a_17567_47# 0.07fF
C636 a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.02fF
C637 a_6375_47# a_7456_47# 0.27fF
C638 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7631_21# 0.22fF
C639 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_6375_47# 0.02fF
C640 a_37255_21# a_38115_47# 0.02fF
C641 a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.02fF
C642 a_28269_289# a_27956_47# 0.00fF
C643 a_27701_47# a_28159_413# 0.12fF
C644 a_28791_21# a_28616_47# 0.62fF
C645 a_27_47# a_543_47# 0.42fF
C646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35139_21# 0.37fF
C647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.45fF
C648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30907_21# 0.37fF
C649 a_25419_47# a_25840_47# 0.23fF
C650 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# 0.24fF
C651 a_23303_47# a_24559_21# 0.12fF
C652 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23819_47# 0.09fF
C653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13144_47# 0.15fF
C654 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12889_47# 1.17fF
C655 a_15260_47# a_15463_413# 0.02fF
C656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5515_21# 0.37fF
C657 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# 0.63fF
C658 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.27fF
C659 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.17fF
C660 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38849_289# 0.10fF
C661 a_6375_47# a_7631_21# 0.12fF
C662 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6891_47# 0.09fF
C663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39358_413# 0.01fF
C664 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9115_413# 0.26fF
C665 a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.63fF
C666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30275_413# 0.26fF
C667 a_12427_47# a_12723_47# 0.07fF
C668 a_28051_47# a_28616_47# 0.01fF
C669 a_27701_47# a_27956_47# 0.22fF
C670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1283_21# 0.37fF
C671 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21608_47# 0.01fF
C672 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23303_47# 0.56fF
C673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30167_47# 0.28fF
C674 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19492_47# 0.01fF
C675 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24037_289# 0.10fF
C676 a_23303_47# a_23819_47# 0.42fF
C677 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26500_47# 0.05fF
C678 a_35999_47# a_36515_47# 0.42fF
C679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_14543_47# 0.27fF
C680 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38115_47# 0.56fF
C681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4775_47# 0.28fF
C682 a_34399_47# a_33883_47# 0.42fF
C683 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.06fF
C684 a_18036_47# a_17579_413# 0.01fF
C685 a_9747_21# a_9572_47# 0.62fF
C686 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7109_289# 0.10fF
C687 a_6375_47# a_6891_47# 0.42fF
C688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_8912_47# 0.15fF
C689 a_34617_289# a_34507_413# 0.23fF
C690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30072_47# 0.15fF
C691 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41474_413# 0.01fF
C692 a_38893_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C693 a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.01fF
C694 a_28269_289# a_28616_47# 0.13fF
C695 a_28051_47# a_28791_21# 0.02fF
C696 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_543_47# 0.28fF
C697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30385_289# 0.29fF
C698 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38281_47# 0.08fF
C699 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28778_413# 0.01fF
C700 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23469_47# 0.65fF
C701 a_23303_47# a_24037_289# 0.16fF
C702 a_25419_47# a_26500_47# 0.27fF
C703 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26675_21# 0.22fF
C704 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13804_47# 0.39fF
C705 a_15920_47# a_15463_413# 0.01fF
C706 sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.12fF
C707 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20314_413# 0.01fF
C708 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_25419_47# 0.02fF
C709 a_41312_47# a_40965_289# 0.13fF
C710 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4993_289# 0.29fF
C711 a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.09fF
C712 a_20152_47# a_20314_413# 0.04fF
C713 a_9007_47# a_9572_47# 0.01fF
C714 a_35139_21# a_34964_47# 0.62fF
C715 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40397_47# 1.17fF
C716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34617_289# 0.29fF
C717 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6541_47# 0.65fF
C718 a_6375_47# a_7109_289# 0.16fF
C719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_10311_47# 0.27fF
C720 a_11863_21# a_12723_47# 0.02fF
C721 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16274_47# 0.01fF
C722 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[8]/D 1.68fF
C723 a_28269_289# a_28791_21# 0.03fF
C724 a_27701_47# a_28616_47# 0.29fF
C725 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D 0.71fF
C726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_29817_47# 0.72fF
C727 a_25419_47# a_26675_21# 0.12fF
C728 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_25935_47# 0.09fF
C729 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18390_47# 0.01fF
C730 a_23303_47# a_23469_47# 1.60fF
C731 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13979_21# 0.37fF
C732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4425_47# 0.72fF
C733 a_38739_413# a_38631_47# 0.21fF
C734 a_17471_47# a_17579_413# 0.21fF
C735 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.11fF
C736 a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.68fF
C737 a_19492_47# a_19695_413# 0.02fF
C738 a_9225_289# a_9572_47# 0.13fF
C739 a_9007_47# a_9747_21# 0.02fF
C740 a_6375_47# a_6541_47# 1.60fF
C741 a_35999_47# a_36165_47# 1.60fF
C742 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16029_47# 0.01fF
C743 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16955_47# 0.99fF
C744 a_28269_289# a_28051_47# 0.50fF
C745 a_27701_47# a_28791_21# 0.10fF
C746 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# 0.63fF
C747 a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.36fF
C748 a_40652_47# a_40855_413# 0.02fF
C749 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9572_47# 0.68fF
C750 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26153_289# 0.10fF
C751 a_25419_47# a_25935_47# 0.42fF
C752 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.11fF
C753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13239_47# 0.28fF
C754 a_15920_47# a_16659_47# 0.00fF
C755 a_15355_47# a_15463_413# 0.21fF
C756 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.73fF
C757 a_17689_289# a_17579_413# 0.23fF
C758 a_17471_47# a_17376_47# 0.13fF
C759 a_9225_289# a_9747_21# 0.03fF
C760 a_8657_47# a_9572_47# 0.29fF
C761 a_27701_47# a_28051_47# 0.49fF
C762 a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.71fF
C763 a_34617_289# a_34964_47# 0.13fF
C764 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.68fF
C765 a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.71fF
C766 a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.02fF
C767 a_25419_47# a_26153_289# 0.16fF
C768 a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.71fF
C769 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.19fF
C770 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_25585_47# 0.65fF
C771 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19695_413# 0.17fF
C772 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9747_21# 0.73fF
C773 a_15355_47# a_15260_47# 0.13fF
C774 a_16095_21# a_16659_47# 0.30fF
C775 a_15573_289# a_15463_413# 0.23fF
C776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13457_289# 0.29fF
C777 a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.36fF
C778 a_17689_289# a_17376_47# 0.00fF
C779 a_17121_47# a_17579_413# 0.12fF
C780 a_35139_21# a_35999_47# 0.02fF
C781 a_41312_47# a_41421_47# 0.04fF
C782 a_9225_289# a_9007_47# 0.50fF
C783 a_20152_47# a_19695_413# 0.01fF
C784 a_8657_47# a_9747_21# 0.10fF
C785 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40965_289# 0.10fF
C786 a_38536_47# a_38849_289# 0.00fF
C787 a_38739_413# a_38281_47# 0.12fF
C788 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_17376_47# 0.01fF
C789 a_40747_47# a_40397_47# 0.49fF
C790 a_27701_47# a_28269_289# 0.41fF
C791 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37434_47# 0.01fF
C792 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.99fF
C793 a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.27fF
C794 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24546_413# 0.01fF
C795 a_25419_47# a_25585_47# 1.60fF
C796 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9007_47# 0.36fF
C797 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19492_47# 0.06fF
C798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_12889_47# 0.72fF
C799 a_15573_289# a_15260_47# 0.00fF
C800 a_15005_47# a_15463_413# 0.12fF
C801 a_16095_21# a_15920_47# 0.62fF
C802 a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.46fF
C803 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.26fF
C804 a_26662_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.01fF
C805 a_17121_47# a_17376_47# 0.22fF
C806 a_8657_47# a_9007_47# 0.49fF
C807 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.12fF
C808 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.12fF
C809 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4259_47# 0.99fF
C810 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22622_47# 0.01fF
C811 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21353_47# 0.08fF
C812 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7618_413# 0.01fF
C813 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9225_289# 0.46fF
C814 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20891_47# 0.09fF
C815 a_15355_47# a_15920_47# 0.01fF
C816 a_15005_47# a_15260_47# 0.22fF
C817 a_27701_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.17fF
C818 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.15fF
C819 a_8657_47# a_9225_289# 0.41fF
C820 a_20152_47# a_20891_47# 0.00fF
C821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41474_413# 0.01fF
C822 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_42051_47# 0.02fF
C823 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11385_47# 0.01fF
C824 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C825 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.08fF
C826 a_22268_47# a_22430_413# 0.04fF
C827 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8657_47# 1.17fF
C828 a_15355_47# a_16095_21# 0.02fF
C829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20314_413# 0.01fF
C830 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20152_47# 0.68fF
C831 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5694_47# 0.01fF
C832 a_15573_289# a_15920_47# 0.13fF
C833 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13913_47# 0.01fF
C834 a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.27fF
C835 a_20327_21# a_20891_47# 0.30fF
C836 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40397_47# 0.72fF
C838 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.08fF
C839 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C840 a_41421_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C841 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36420_47# 0.06fF
C842 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11219_47# 0.02fF
C843 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41666_47# 0.01fF
C844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.45fF
C845 a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.37fF
C846 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.63fF
C847 a_21703_47# a_21799_47# 0.07fF
C848 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23927_413# 0.17fF
C849 a_21608_47# a_21811_413# 0.02fF
C850 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.63fF
C851 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20327_21# 0.73fF
C852 a_15005_47# a_15920_47# 0.29fF
C853 a_15573_289# a_16095_21# 0.03fF
C854 a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.39fF
C855 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.19fF
C856 a_20327_21# a_20152_47# 0.62fF
C857 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.63fF
C858 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# 0.63fF
C859 a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.63fF
C860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16955_47# 0.56fF
C861 a_193_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.33fF
C862 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# 0.27fF
C863 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23724_47# 0.06fF
C864 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C865 a_24384_47# a_24546_413# 0.04fF
C866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9572_47# 0.39fF
C867 a_15573_289# a_15355_47# 0.50fF
C868 a_15005_47# a_16095_21# 0.10fF
C869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.19fF
C870 a_38536_47# a_38115_47# 0.23fF
C871 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_15260_47# 0.01fF
C872 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.37fF
C873 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33202_47# 0.01fF
C874 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39196_47# 0.68fF
C875 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.12fF
C876 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.53fF
C877 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34049_47# 1.17fF
C878 a_193_47# a_761_289# 0.41fF
C879 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.27fF
C880 a_22268_47# a_21811_413# 0.01fF
C881 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25123_47# 0.09fF
C882 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.45fF
C883 a_41487_21# a_41312_47# 0.62fF
C884 a_23724_47# a_23927_413# 0.02fF
C885 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_19071_47# 0.02fF
C886 a_23819_47# a_23915_47# 0.07fF
C887 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40747_47# 0.36fF
C888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9747_21# 0.37fF
C889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19695_413# 0.26fF
C890 a_15005_47# a_15355_47# 0.49fF
C891 a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C892 a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.28fF
C893 a_6796_47# a_6999_413# 0.02fF
C894 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21965_47# 0.01fF
C895 a_34661_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C896 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.08fF
C897 a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.86fF
C898 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_761_289# 0.10fF
C899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24546_413# 0.01fF
C900 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24384_47# 0.68fF
C901 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.56fF
C902 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19587_47# 0.09fF
C903 a_40397_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C904 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9007_47# 0.28fF
C905 a_15005_47# a_15573_289# 0.41fF
C906 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19492_47# 0.15fF
C907 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37255_21# 0.73fF
C908 a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.29fF
C909 a_14543_47# a_14839_47# 0.07fF
C910 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.12fF
C911 a_26662_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.01fF
C912 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21799_47# 0.02fF
C913 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11231_413# 0.01fF
C914 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4259_47# 0.56fF
C915 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6796_47# 0.01fF
C916 a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.36fF
C917 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34507_413# 0.17fF
C918 a_27_47# a_761_289# 0.16fF
C919 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_193_47# 0.65fF
C920 a_639_47# a_543_47# 0.07fF
C921 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19805_289# 0.10fF
C922 a_19071_47# a_19587_47# 0.42fF
C923 a_22268_47# a_23007_47# 0.00fF
C924 a_21703_47# a_21811_413# 0.21fF
C925 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24559_21# 0.73fF
C926 a_24384_47# a_23927_413# 0.01fF
C927 a_37080_47# a_37819_47# 0.00fF
C928 a_36515_47# a_36623_413# 0.21fF
C929 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9225_289# 0.29fF
C930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20891_47# 0.27fF
C931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7618_413# 0.01fF
C932 a_39371_21# a_39935_47# 0.30fF
C933 a_7456_47# a_6999_413# 0.01fF
C934 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13501_47# 0.01fF
C935 a_27701_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.72fF
C936 a_12723_47# a_13144_47# 0.23fF
C937 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33883_47# 0.02fF
C938 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_39935_47# 0.01fF
C939 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_42051_47# 0.26fF
C940 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11028_47# 0.53fF
C941 a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C942 a_21703_47# a_21608_47# 0.13fF
C943 a_22443_21# a_23007_47# 0.30fF
C944 a_21921_289# a_21811_413# 0.23fF
C945 a_27_47# a_193_47# 1.60fF
C946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 8.78fF
C947 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19237_47# 0.65fF
C948 a_19071_47# a_19805_289# 0.16fF
C949 a_3578_47# a_3399_21# 0.04fF
C950 a_3333_47# a_3224_47# 0.04fF
C951 a_25840_47# a_26043_413# 0.02fF
C952 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23819_47# 0.36fF
C953 a_13979_21# a_14158_47# 0.04fF
C954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_8657_47# 0.72fF
C955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20152_47# 0.39fF
C956 a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.71fF
C957 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C958 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.19fF
C959 a_41312_47# a_40231_47# 0.27fF
C960 a_13979_21# a_14839_47# 0.02fF
C961 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.11fF
C962 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# 0.24fF
C963 a_35139_21# a_35318_47# 0.04fF
C964 a_34964_47# a_35073_47# 0.04fF
C965 a_10607_47# a_11028_47# 0.23fF
C966 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# 0.24fF
C967 a_1283_21# a_1462_47# 0.04fF
C968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36420_47# 0.15fF
C969 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36733_289# 0.46fF
C970 a_27_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.71fF
C971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_761_289# 0.29fF
C972 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_193_47# 0.04fF
C973 a_6079_47# a_6375_47# 0.07fF
C974 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.12fF
C975 a_22443_21# a_22268_47# 0.62fF
C976 a_651_413# a_543_47# 0.21fF
C977 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24037_289# 0.46fF
C978 a_19071_47# a_19237_47# 1.60fF
C979 a_21921_289# a_21608_47# 0.00fF
C980 a_21353_47# a_21811_413# 0.12fF
C981 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23927_413# 0.26fF
C982 a_24384_47# a_25123_47# 0.00fF
C983 a_23819_47# a_23927_413# 0.21fF
C984 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20327_21# 0.37fF
C985 a_7565_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C986 a_7456_47# a_8195_47# 0.00fF
C987 a_6891_47# a_6999_413# 0.21fF
C988 a_12723_47# a_13804_47# 0.27fF
C989 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18036_47# 0.05fF
C990 a_36733_289# a_36420_47# 0.00fF
C991 a_36165_47# a_36623_413# 0.12fF
C992 a_34507_413# a_34049_47# 0.12fF
C993 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11688_47# 0.05fF
C994 a_21353_47# a_21608_47# 0.22fF
C995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_193_47# 0.70fF
C996 a_1847_47# a_1283_21# 0.30fF
C997 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5037_47# 0.01fF
C998 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.04fF
C999 a_448_47# a_543_47# 0.13fF
C1000 a_21703_47# a_22268_47# 0.01fF
C1001 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23469_47# 1.17fF
C1002 a_23819_47# a_23724_47# 0.13fF
C1003 a_24037_289# a_23927_413# 0.23fF
C1004 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23724_47# 0.15fF
C1005 a_26500_47# a_26043_413# 0.01fF
C1006 a_24559_21# a_25123_47# 0.30fF
C1007 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_15005_47# 0.08fF
C1008 a_6891_47# a_6796_47# 0.13fF
C1009 a_7631_21# a_8195_47# 0.30fF
C1010 a_7109_289# a_6999_413# 0.23fF
C1011 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34964_47# 0.68fF
C1012 a_12723_47# a_13979_21# 0.12fF
C1013 a_16955_47# a_18036_47# 0.27fF
C1014 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18211_21# 0.22fF
C1015 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39196_47# 0.39fF
C1016 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21811_413# 0.01fF
C1017 a_36515_47# a_37080_47# 0.01fF
C1018 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16955_47# 0.02fF
C1019 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34049_47# 0.72fF
C1020 a_10607_47# a_11688_47# 0.27fF
C1021 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11863_21# 0.22fF
C1022 a_38631_47# a_39371_21# 0.02fF
C1023 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# 0.44fF
C1024 a_5515_21# a_6375_47# 0.02fF
C1025 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.45fF
C1026 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_25123_47# 0.27fF
C1027 a_1108_47# a_1283_21# 0.62fF
C1028 a_21921_289# a_22268_47# 0.13fF
C1029 a_21703_47# a_22443_21# 0.02fF
C1030 a_18211_21# a_18390_47# 0.04fF
C1031 a_18036_47# a_18145_47# 0.04fF
C1032 a_24037_289# a_23724_47# 0.00fF
C1033 a_23469_47# a_23927_413# 0.12fF
C1034 a_24559_21# a_24384_47# 0.62fF
C1035 a_40231_47# a_39371_21# 0.02fF
C1036 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39196_47# 0.02fF
C1037 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C1038 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C1039 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40747_47# 0.28fF
C1040 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.12fF
C1041 a_7631_21# a_7456_47# 0.62fF
C1042 a_7109_289# a_6796_47# 0.00fF
C1043 a_6541_47# a_6999_413# 0.12fF
C1044 a_37819_47# a_38281_47# 0.01fF
C1045 a_12723_47# a_13239_47# 0.42fF
C1046 a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.71fF
C1047 a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.36fF
C1048 a_16955_47# a_18211_21# 0.12fF
C1049 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17471_47# 0.09fF
C1050 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[18]/D 1.68fF
C1051 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21608_47# 0.53fF
C1052 a_10607_47# a_11863_21# 0.12fF
C1053 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11123_47# 0.09fF
C1054 a_21921_289# a_22443_21# 0.03fF
C1055 a_21353_47# a_22268_47# 0.29fF
C1056 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_27_47# 0.53fF
C1057 a_1108_47# a_543_47# 0.01fF
C1058 a_26500_47# a_27239_47# 0.00fF
C1059 a_25935_47# a_26043_413# 0.21fF
C1060 a_23819_47# a_24384_47# 0.01fF
C1061 a_23469_47# a_23724_47# 0.22fF
C1062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24384_47# 0.39fF
C1063 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# 0.63fF
C1064 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37255_21# 0.37fF
C1065 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32545_47# 0.01fF
C1066 a_6541_47# a_6796_47# 0.22fF
C1067 a_6891_47# a_7456_47# 0.01fF
C1068 a_12723_47# a_13457_289# 0.16fF
C1069 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17689_289# 0.10fF
C1070 a_16955_47# a_17471_47# 0.42fF
C1071 a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.02fF
C1072 a_21187_47# a_21608_47# 0.23fF
C1073 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# 0.24fF
C1074 a_10607_47# a_11123_47# 0.42fF
C1075 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6541_47# 0.08fF
C1076 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/CLK 0.06fF
C1077 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34507_413# 0.26fF
C1078 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.08fF
C1079 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24559_21# 0.37fF
C1080 a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.71fF
C1081 a_21921_289# a_21703_47# 0.50fF
C1082 a_21353_47# a_22443_21# 0.10fF
C1083 a_24037_289# a_24384_47# 0.13fF
C1084 a_23819_47# a_24559_21# 0.02fF
C1085 a_25935_47# a_25840_47# 0.13fF
C1086 a_26675_21# a_27239_47# 0.30fF
C1087 a_26153_289# a_26043_413# 0.23fF
C1088 a_36733_289# a_37255_21# 0.03fF
C1089 a_36165_47# a_37080_47# 0.29fF
C1090 a_34964_47# a_34049_47# 0.29fF
C1091 a_33023_21# a_33883_47# 0.02fF
C1092 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35999_47# 0.99fF
C1093 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32379_47# 0.02fF
C1094 a_38281_47# a_39371_21# 0.10fF
C1095 a_38849_289# a_38631_47# 0.50fF
C1096 a_40397_47# a_40965_289# 0.41fF
C1097 a_7109_289# a_7456_47# 0.13fF
C1098 a_6891_47# a_7631_21# 0.02fF
C1099 a_12723_47# a_12889_47# 1.60fF
C1100 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.27fF
C1101 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17121_47# 0.65fF
C1102 a_16955_47# a_17689_289# 0.16fF
C1103 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_22268_47# 0.05fF
C1104 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.08fF
C1105 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18775_47# 0.09fF
C1106 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# 0.63fF
C1107 a_21353_47# a_21703_47# 0.49fF
C1108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23819_47# 0.28fF
C1109 a_26153_289# a_25840_47# 0.00fF
C1110 a_26675_21# a_26500_47# 0.62fF
C1111 a_25585_47# a_26043_413# 0.12fF
C1112 a_24037_289# a_24559_21# 0.03fF
C1113 a_23469_47# a_24384_47# 0.29fF
C1114 a_35999_47# a_36420_47# 0.23fF
C1115 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26854_47# 0.01fF
C1116 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# 0.24fF
C1117 a_34304_47# a_33883_47# 0.23fF
C1118 a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.24fF
C1119 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39196_47# 0.05fF
C1120 a_7109_289# a_7631_21# 0.03fF
C1121 a_6541_47# a_7456_47# 0.29fF
C1122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.19fF
C1123 a_16955_47# a_17121_47# 1.60fF
C1124 a_21187_47# a_22268_47# 0.27fF
C1125 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_22443_21# 0.22fF
C1126 a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.63fF
C1127 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18036_47# 0.68fF
C1128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36733_289# 0.29fF
C1129 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.12fF
C1130 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.11fF
C1131 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_2143_47# 0.02fF
C1132 a_21353_47# a_21921_289# 0.41fF
C1133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24037_289# 0.29fF
C1134 a_25585_47# a_25840_47# 0.22fF
C1135 a_4425_47# a_3963_47# 0.01fF
C1136 a_23469_47# a_24559_21# 0.10fF
C1137 a_24037_289# a_23819_47# 0.50fF
C1138 a_25935_47# a_26500_47# 0.01fF
C1139 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26609_47# 0.01fF
C1140 a_34964_47# a_34507_413# 0.01fF
C1141 a_7109_289# a_6891_47# 0.50fF
C1142 a_6541_47# a_7631_21# 0.10fF
C1143 a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.36fF
C1144 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32957_47# 0.01fF
C1145 a_11688_47# a_11850_413# 0.04fF
C1146 a_33587_47# a_33883_47# 0.07fF
C1147 a_16095_21# a_16274_47# 0.04fF
C1148 a_15920_47# a_16029_47# 0.04fF
C1149 a_21187_47# a_22443_21# 0.12fF
C1150 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21703_47# 0.09fF
C1151 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.02fF
C1152 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18211_21# 0.73fF
C1153 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2921_47# 0.01fF
C1154 a_38281_47# a_38849_289# 0.41fF
C1155 a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.36fF
C1156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_23469_47# 0.72fF
C1157 a_23469_47# a_23819_47# 0.49fF
C1158 a_26153_289# a_26500_47# 0.13fF
C1159 a_25935_47# a_26675_21# 0.02fF
C1160 a_6541_47# a_6891_47# 0.49fF
C1161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34964_47# 0.39fF
C1162 a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.01fF
C1163 a_11123_47# a_11219_47# 0.07fF
C1164 a_11028_47# a_11231_413# 0.02fF
C1165 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_4259_47# 0.02fF
C1166 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21921_289# 0.10fF
C1167 a_21187_47# a_21703_47# 0.42fF
C1168 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17471_47# 0.36fF
C1169 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C1170 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2755_47# 0.02fF
C1171 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38536_47# 0.06fF
C1172 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_10607_47# 0.02fF
C1173 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.11fF
C1174 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2877_289# 0.10fF
C1175 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33023_21# 0.22fF
C1176 a_25585_47# a_26500_47# 0.29fF
C1177 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C1178 a_23469_47# a_24037_289# 0.41fF
C1179 a_26153_289# a_26675_21# 0.03fF
C1180 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_31767_47# 0.02fF
C1181 a_35703_47# a_36165_47# 0.01fF
C1182 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32391_413# 0.01fF
C1183 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.08fF
C1184 a_6541_47# a_7109_289# 0.41fF
C1185 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21353_47# 0.65fF
C1186 a_21187_47# a_21921_289# 0.16fF
C1187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.45fF
C1188 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36515_47# 0.09fF
C1189 a_35999_47# a_37255_21# 0.12fF
C1190 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37242_413# 0.01fF
C1191 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17689_289# 0.46fF
C1192 a_35139_21# a_33883_47# 0.12fF
C1193 a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.09fF
C1194 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.11fF
C1195 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16082_413# 0.01fF
C1196 a_38115_47# a_38631_47# 0.42fF
C1197 a_2143_47# a_2877_289# 0.16fF
C1198 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_34304_47# 0.01fF
C1199 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2309_47# 0.65fF
C1200 a_26153_289# a_25935_47# 0.50fF
C1201 a_25585_47# a_26675_21# 0.10fF
C1202 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[7]/D 1.68fF
C1203 a_31767_47# a_33023_21# 0.12fF
C1204 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32283_47# 0.09fF
C1205 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.12fF
C1206 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32188_47# 0.53fF
C1207 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C1208 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4871_47# 0.02fF
C1209 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.02fF
C1210 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# 0.63fF
C1211 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12042_47# 0.01fF
C1212 a_11688_47# a_11231_413# 0.01fF
C1213 a_21187_47# a_21353_47# 1.60fF
C1214 a_40652_47# a_40397_47# 0.22fF
C1215 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17121_47# 1.17fF
C1216 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14158_47# 0.01fF
C1217 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_8195_47# 0.01fF
C1218 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11341_289# 0.10fF
C1219 a_34399_47# a_34304_47# 0.13fF
C1220 a_35139_21# a_35703_47# 0.30fF
C1221 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40965_289# 0.46fF
C1222 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14839_47# 0.99fF
C1223 a_2143_47# a_2309_47# 1.60fF
C1224 a_31767_47# a_32283_47# 0.42fF
C1225 a_25585_47# a_25935_47# 0.49fF
C1226 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32501_289# 0.10fF
C1227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35999_47# 0.56fF
C1228 a_31767_47# a_32188_47# 0.23fF
C1229 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# 0.24fF
C1230 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_27239_47# 0.01fF
C1231 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_31471_47# 0.01fF
C1232 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11797_47# 0.01fF
C1233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18775_47# 0.27fF
C1234 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31086_47# 0.01fF
C1235 a_8491_47# a_8195_47# 0.07fF
C1236 a_10607_47# a_11341_289# 0.16fF
C1237 a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.46fF
C1238 sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.12fF
C1239 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_10773_47# 0.65fF
C1240 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D 0.01fF
C1241 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.12fF
C1242 a_25585_47# a_26153_289# 0.41fF
C1243 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_31933_47# 0.65fF
C1244 a_31767_47# a_32501_289# 0.16fF
C1245 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36165_47# 0.65fF
C1246 a_35999_47# a_36733_289# 0.16fF
C1247 a_34617_289# a_33883_47# 0.16fF
C1248 a_13804_47# a_13913_47# 0.04fF
C1249 a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.71fF
C1250 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32848_47# 0.05fF
C1251 a_38115_47# a_38281_47# 1.60fF
C1252 a_27535_47# a_27239_47# 0.07fF
C1253 a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.01fF
C1254 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.12fF
C1255 sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.12fF
C1256 a_11688_47# a_12427_47# 0.00fF
C1257 a_11123_47# a_11231_413# 0.21fF
C1258 a_31767_47# a_31471_47# 0.07fF
C1259 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.12fF
C1260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18036_47# 0.39fF
C1261 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3386_413# 0.01fF
C1262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.19fF
C1263 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2767_413# 0.01fF
C1264 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30841_47# 0.01fF
C1265 a_7153_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C1266 a_10607_47# a_10773_47# 1.60fF
C1267 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.17fF
C1268 a_805_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C1269 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.06fF
C1270 a_1847_47# a_2143_47# 0.07fF
C1271 a_31767_47# a_31933_47# 1.60fF
C1272 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12723_47# 0.99fF
C1273 a_31767_47# a_32848_47# 0.27fF
C1274 a_26197_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C1275 a_9681_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.01fF
C1276 a_11123_47# a_11028_47# 0.13fF
C1277 a_11863_21# a_12427_47# 0.30fF
C1278 a_40397_47# a_39935_47# 0.01fF
C1279 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19849_47# 0.01fF
C1280 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_13144_47# 0.01fF
C1281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.19fF
C1282 a_30429_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C1283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18211_21# 0.37fF
C1284 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_1462_47# 0.01fF
C1285 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2564_47# 0.53fF
C1286 a_8491_47# a_7631_21# 0.02fF
C1287 a_639_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.02fF
C1288 a_651_413# a_761_289# 0.23fF
C1289 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.01fF
C1290 a_6987_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.02fF
C1291 a_40843_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.02fF
C1292 a_38739_413# a_38849_289# 0.23fF
C1293 a_41487_21# a_40397_47# 0.10fF
C1294 a_40747_47# a_40965_289# 0.50fF
C1295 a_34399_47# a_35139_21# 0.02fF
C1296 a_27535_47# a_26675_21# 0.02fF
C1297 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4883_413# 0.01fF
C1298 a_26031_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.02fF
C1299 a_11863_21# a_11688_47# 0.62fF
C1300 a_31767_47# a_30907_21# 0.02fF
C1301 a_30263_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.02fF
C1302 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35318_47# 0.01fF
C1303 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19683_47# 0.02fF
C1304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17471_47# 0.28fF
C1305 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# 0.24fF
C1306 a_2143_47# a_2564_47# 0.23fF
C1307 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_32188_47# 0.01fF
C1308 a_448_47# a_761_289# 0.00fF
C1309 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.09fF
C1310 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.19fF
C1311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38536_47# 0.15fF
C1312 a_651_413# a_193_47# 0.12fF
C1313 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# 0.63fF
C1314 a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.36fF
C1315 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.01fF
C1316 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4680_47# 0.53fF
C1317 a_11123_47# a_11688_47# 0.01fF
C1318 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[3]/D 1.68fF
C1319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37242_413# 0.01fF
C1320 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2767_413# 0.17fF
C1321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17689_289# 0.29fF
C1322 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.19fF
C1323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16082_413# 0.01fF
C1324 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3224_47# 0.05fF
C1325 a_8657_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C1326 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C1327 a_448_47# a_193_47# 0.22fF
C1328 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.08fF
C1329 a_41312_47# a_40855_413# 0.01fF
C1330 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.59fF
C1331 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.01fF
C1332 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24738_47# 0.01fF
C1333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.45fF
C1334 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# 0.24fF
C1335 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40652_47# 0.06fF
C1336 a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.02fF
C1337 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.08fF
C1338 a_39550_47# a_39371_21# 0.04fF
C1339 a_39305_47# a_39196_47# 0.04fF
C1340 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13335_47# 0.02fF
C1341 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# 0.24fF
C1342 a_27701_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C1343 a_31933_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.08fF
C1344 a_11123_47# a_11863_21# 0.02fF
C1345 a_3963_47# a_4259_47# 0.07fF
C1346 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6375_47# 0.99fF
C1347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17121_47# 0.72fF
C1348 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1462_47# 0.01fF
C1349 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2564_47# 0.06fF
C1350 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3399_21# 0.22fF
C1351 a_2143_47# a_3224_47# 0.27fF
C1352 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_38115_47# 0.02fF
C1353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40965_289# 0.29fF
C1354 a_34617_289# a_34399_47# 0.50fF
C1355 a_10311_47# a_10607_47# 0.07fF
C1356 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.53fF
C1357 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[12]/D 1.68fF
C1358 a_1108_47# a_761_289# 0.13fF
C1359 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30732_47# 0.05fF
C1360 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24493_47# 0.01fF
C1361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_14839_47# 0.56fF
C1362 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36623_413# 0.17fF
C1363 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# 0.63fF
C1364 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.27fF
C1365 a_40231_47# a_40397_47# 1.60fF
C1366 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5340_47# 0.05fF
C1367 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23007_47# 0.01fF
C1368 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3963_47# 0.09fF
C1369 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1217_47# 0.01fF
C1370 a_2143_47# a_3399_21# 0.12fF
C1371 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2659_47# 0.09fF
C1372 a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.36fF
C1373 a_1108_47# a_193_47# 0.29fF
C1374 a_1270_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.01fF
C1375 a_448_47# a_27_47# 0.23fF
C1376 a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.29fF
C1377 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.24fF
C1378 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25419_47# 0.99fF
C1379 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30907_21# 0.22fF
C1380 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_29651_47# 0.02fF
C1381 a_36420_47# a_36623_413# 0.02fF
C1382 a_29651_47# a_30732_47# 0.27fF
C1383 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5515_21# 0.22fF
C1384 a_23303_47# a_23007_47# 0.07fF
C1385 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36611_47# 0.02fF
C1386 a_18036_47# a_18775_47# 0.00fF
C1387 a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C1388 a_3399_21# a_4259_47# 0.02fF
C1389 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.53fF
C1390 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19695_413# 0.01fF
C1391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3386_413# 0.01fF
C1392 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3224_47# 0.68fF
C1393 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35126_413# 0.01fF
C1394 a_2143_47# a_2659_47# 0.42fF
C1395 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.72fF
C1396 a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.02fF
C1397 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/CLK 0.01fF
C1398 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.05fF
C1399 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.26fF
C1400 a_19805_289# a_19587_47# 0.50fF
C1401 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39935_47# 0.09fF
C1402 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25840_47# 0.01fF
C1403 a_29651_47# a_30907_21# 0.12fF
C1404 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30167_47# 0.09fF
C1405 a_7810_47# a_7631_21# 0.04fF
C1406 a_7565_47# a_7456_47# 0.04fF
C1407 a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C1408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_12723_47# 0.56fF
C1409 a_14543_47# a_15005_47# 0.01fF
C1410 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4775_47# 0.09fF
C1411 a_41487_21# a_42051_47# 0.30fF
C1412 a_40747_47# a_40652_47# 0.13fF
C1413 a_18211_21# a_18775_47# 0.30fF
C1414 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.53fF
C1415 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12889_47# 0.08fF
C1416 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41487_21# 0.67fF
C1417 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19492_47# 0.53fF
C1418 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3399_21# 0.73fF
C1419 a_11341_289# a_11231_413# 0.23fF
C1420 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2564_47# 0.01fF
C1421 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.15fF
C1422 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.27fF
C1423 a_19237_47# a_19587_47# 0.49fF
C1424 a_1108_47# a_27_47# 0.27fF
C1425 a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C1426 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30385_289# 0.10fF
C1427 a_29651_47# a_30167_47# 0.42fF
C1428 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.12fF
C1429 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13347_413# 0.01fF
C1430 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4993_289# 0.10fF
C1431 a_23303_47# a_22443_21# 0.02fF
C1432 a_41487_21# a_41666_47# 0.04fF
C1433 a_18211_21# a_18036_47# 0.62fF
C1434 a_30072_47# a_29651_47# 0.23fF
C1435 a_11341_289# a_11028_47# 0.00fF
C1436 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37080_47# 0.68fF
C1437 a_19071_47# a_19492_47# 0.23fF
C1438 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# 0.24fF
C1439 a_10773_47# a_11231_413# 0.12fF
C1440 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.71fF
C1441 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2659_47# 0.36fF
C1442 a_19237_47# a_19805_289# 0.41fF
C1443 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.27fF
C1444 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.12fF
C1445 a_25123_47# a_25419_47# 0.07fF
C1446 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_29817_47# 0.65fF
C1447 a_29651_47# a_30385_289# 0.16fF
C1448 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/D 1.68fF
C1449 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13144_47# 0.53fF
C1450 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4425_47# 0.65fF
C1451 a_17471_47# a_18036_47# 0.01fF
C1452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.45fF
C1453 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20152_47# 0.05fF
C1454 a_10773_47# a_11028_47# 0.22fF
C1455 a_39196_47# a_39935_47# 0.00fF
C1456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_2767_413# 0.26fF
C1457 a_6079_47# a_6541_47# 0.01fF
C1458 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.01fF
C1459 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 0.39fF
C1460 a_29651_47# a_29817_47# 1.60fF
C1461 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24081_47# 0.01fF
C1462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40652_47# 0.15fF
C1463 a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.27fF
C1464 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.71fF
C1465 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# 0.24fF
C1466 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19071_47# 0.99fF
C1467 a_17689_289# a_18036_47# 0.13fF
C1468 a_17471_47# a_18211_21# 0.02fF
C1469 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38631_47# 0.36fF
C1470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_6375_47# 0.56fF
C1471 a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.05fF
C1472 a_11341_289# a_11688_47# 0.13fF
C1473 a_19071_47# a_20152_47# 0.27fF
C1474 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20327_21# 0.22fF
C1475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_2564_47# 0.15fF
C1476 a_16659_47# a_16955_47# 0.07fF
C1477 a_40747_47# a_41487_21# 0.02fF
C1478 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40231_47# 0.99fF
C1479 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.12fF
C1480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.45fF
C1481 a_24559_21# a_25419_47# 0.02fF
C1482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36623_413# 0.26fF
C1483 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.11fF
C1484 a_39305_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C1485 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13804_47# 0.05fF
C1486 a_11863_21# a_12042_47# 0.04fF
C1487 a_11688_47# a_11797_47# 0.04fF
C1488 a_17689_289# a_18211_21# 0.03fF
C1489 a_17121_47# a_18036_47# 0.29fF
C1490 sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.12fF
C1491 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33883_47# 0.99fF
C1492 a_19071_47# a_20327_21# 0.12fF
C1493 a_10773_47# a_11688_47# 0.29fF
C1494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3963_47# 0.27fF
C1495 a_11341_289# a_11863_21# 0.03fF
C1496 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15617_47# 0.01fF
C1497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_25419_47# 0.56fF
C1498 a_36733_289# a_36623_413# 0.23fF
C1499 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C1500 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13979_21# 0.22fF
C1501 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.36fF
C1502 a_17689_289# a_17471_47# 0.50fF
C1503 a_17121_47# a_18211_21# 0.10fF
C1504 a_9269_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.01fF
C1505 a_11341_289# a_11123_47# 0.50fF
C1506 a_10773_47# a_11863_21# 0.10fF
C1507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3224_47# 0.39fF
C1508 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35703_47# 0.09fF
C1509 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.27fF
C1510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35126_413# 0.01fF
C1511 a_16095_21# a_16955_47# 0.02fF
C1512 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15451_47# 0.02fF
C1513 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15463_413# 0.17fF
C1514 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38281_47# 1.17fF
C1515 a_37255_21# a_37080_47# 0.62fF
C1516 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25585_47# 0.08fF
C1517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39935_47# 0.27fF
C1518 a_26675_21# a_26854_47# 0.04fF
C1519 a_26500_47# a_26609_47# 0.04fF
C1520 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.63fF
C1521 a_38631_47# a_39196_47# 0.01fF
C1522 a_32283_47# a_32379_47# 0.07fF
C1523 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13239_47# 0.09fF
C1524 a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.02fF
C1525 a_17121_47# a_17471_47# 0.49fF
C1526 a_9103_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.02fF
C1527 a_10607_47# a_9747_21# 0.02fF
C1528 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39935_47# 0.36fF
C1529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41487_21# 0.37fF
C1530 a_10773_47# a_11123_47# 0.49fF
C1531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3399_21# 0.37fF
C1532 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C1533 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15260_47# 0.06fF
C1534 a_40747_47# a_40231_47# 0.42fF
C1535 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13457_289# 0.10fF
C1536 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22430_413# 0.01fF
C1537 a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C1538 a_33883_47# a_34049_47# 1.60fF
C1539 a_17121_47# a_17689_289# 0.41fF
C1540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37080_47# 0.39fF
C1541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_2659_47# 0.28fF
C1542 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_17121_47# 0.08fF
C1543 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28970_47# 0.01fF
C1544 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16659_47# 0.09fF
C1545 a_17376_47# a_17579_413# 0.02fF
C1546 a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.71fF
C1547 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20506_47# 0.01fF
C1548 a_34964_47# a_35126_413# 0.04fF
C1549 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[5]/D 1.68fF
C1550 a_29355_47# a_29651_47# 0.07fF
C1551 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.12fF
C1552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.45fF
C1553 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_12889_47# 0.65fF
C1554 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[15]/D 1.68fF
C1555 a_36733_289# a_37080_47# 0.13fF
C1556 a_10773_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.08fF
C1557 a_38849_289# a_39371_21# 0.03fF
C1558 a_38281_47# a_39196_47# 0.29fF
C1559 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[17]/D 1.68fF
C1560 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15920_47# 0.68fF
C1561 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28725_47# 0.01fF
C1562 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.11fF
C1563 a_34399_47# a_34495_47# 0.07fF
C1564 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10607_47# 0.99fF
C1565 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34399_47# 0.36fF
C1566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19071_47# 0.56fF
C1567 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31767_47# 0.99fF
C1568 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28313_47# 0.01fF
C1569 a_32848_47# a_33010_413# 0.04fF
C1570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38631_47# 0.28fF
C1571 a_20327_21# a_20506_47# 0.04fF
C1572 a_20152_47# a_20261_47# 0.04fF
C1573 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36420_47# 0.53fF
C1574 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.53fF
C1575 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# 0.24fF
C1576 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_8195_47# 0.36fF
C1577 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37434_47# 0.01fF
C1578 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40231_47# 0.56fF
C1579 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16095_21# 0.73fF
C1580 a_32283_47# a_33023_21# 0.02fF
C1581 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.08fF
C1582 a_32283_47# a_32391_413# 0.21fF
C1583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.19fF
C1584 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21811_413# 0.17fF
C1585 a_5340_47# a_5502_413# 0.04fF
C1586 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28147_47# 0.02fF
C1587 a_28791_21# a_29651_47# 0.02fF
C1588 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_27239_47# 0.36fF
C1589 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_40231_47# 0.02fF
C1590 a_32188_47# a_32391_413# 0.02fF
C1591 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.11fF
C1592 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_31471_47# 0.36fF
C1593 a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.01fF
C1594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33883_47# 0.56fF
C1595 a_32957_47# a_32848_47# 0.04fF
C1596 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7456_47# 0.02fF
C1597 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33202_47# 0.01fF
C1598 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24738_47# 0.01fF
C1599 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15355_47# 0.36fF
C1600 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C1601 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0.36fF
C1602 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_30072_47# 0.01fF
C1603 a_32501_289# a_33023_21# 0.03fF
C1604 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.11fF
C1605 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_34049_47# 0.08fF
C1606 a_32283_47# a_32188_47# 0.13fF
C1607 a_33023_21# a_33587_47# 0.30fF
C1608 a_32501_289# a_32391_413# 0.23fF
C1609 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_21187_47# 0.02fF
C1610 a_4680_47# a_4883_413# 0.02fF
C1611 a_4775_47# a_4871_47# 0.07fF
C1612 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26500_47# 0.02fF
C1613 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21608_47# 0.06fF
C1614 a_37819_47# a_38115_47# 0.07fF
C1615 a_12427_47# a_12889_47# 0.01fF
C1616 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1617 a_41421_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1618 sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1619 a_41009_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1620 a_40843_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1621 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1622 a_39305_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1623 a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1624 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1625 a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1626 a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1627 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1628 a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1629 a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1630 a_40397_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1631 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1632 a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1633 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1634 a_38893_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1635 a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1636 a_37189_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1637 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1638 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1639 a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1640 a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.41fF
C1641 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.79fF
C1642 a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.43fF
C1643 a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.44fF
C1644 a_38281_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.47fF
C1645 sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1646 a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.70fF
C1647 sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1648 a_36777_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1649 a_36611_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1650 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1651 a_35073_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1652 a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1653 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1654 a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1655 a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1656 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1657 a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1658 a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1659 a_36165_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1660 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1661 a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1662 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1663 a_34661_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1664 a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1665 a_32957_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1666 a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1667 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1668 a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1669 a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.39fF
C1670 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.75fF
C1671 a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1672 a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.43fF
C1673 a_34049_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.64fF
C1674 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1675 a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.75fF
C1676 sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1677 a_32545_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1678 a_32379_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1679 a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1680 a_30841_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1681 a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1682 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1683 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1684 a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1685 a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1686 a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1687 a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1688 a_31933_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1689 sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1690 a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1691 sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1692 a_30429_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1693 a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1694 a_28725_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1695 a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1696 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1697 a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1698 a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.60fF
C1699 a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.71fF
C1700 a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1701 a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.59fF
C1702 a_29817_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.70fF
C1703 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1704 a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.80fF
C1705 sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1706 a_28313_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1707 a_28147_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1708 a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1709 a_26609_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1710 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1711 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1712 a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1713 a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1714 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1715 a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1716 a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1717 a_27701_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1718 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1719 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1720 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1721 a_26197_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1722 a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1723 a_24493_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1724 a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1725 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1726 a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1727 a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.52fF
C1728 a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.67fF
C1729 a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1730 a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1731 a_25585_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.76fF
C1732 sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.59fF
C1733 a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.96fF
C1734 sky130_fd_sc_hd__dfrbp_1_0[11]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1735 a_24081_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1736 a_23915_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1737 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1738 a_22377_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1739 a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1740 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1741 a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1742 a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1743 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1744 a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1745 a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1746 a_23469_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1747 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1748 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1749 sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1750 a_21965_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1751 a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1752 a_20261_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1753 a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1754 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1755 a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1756 a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.30fF
C1757 a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.63fF
C1758 a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1759 a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1760 a_21353_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.84fF
C1761 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.59fF
C1762 a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.08fF
C1763 sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1764 a_19849_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1765 a_19683_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1766 a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1767 a_18145_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1768 a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1769 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1770 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1771 a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1772 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1773 a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1774 a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1775 a_19237_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1776 sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1777 a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1778 sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1779 a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1780 a_16029_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1781 a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1782 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1783 a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1784 a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.23fF
C1785 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.59fF
C1786 a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1787 a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1788 a_17121_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.88fF
C1789 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.59fF
C1790 a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.15fF
C1791 sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1792 a_15617_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1793 a_15451_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1794 a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1795 a_13913_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1796 a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1797 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1798 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1799 a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1800 a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1801 a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1802 a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1803 a_15005_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1804 sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1805 a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1806 sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1807 a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1808 a_11797_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1809 a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1810 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1811 a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1812 a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.23fF
C1813 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.55fF
C1814 a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1815 a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1816 a_12889_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.91fF
C1817 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.59fF
C1818 a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.19fF
C1819 sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1820 a_11385_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1821 a_11219_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1822 a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1823 a_9681_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1824 a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1825 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1826 a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1827 a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1828 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1829 a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1830 a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1831 a_10773_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1832 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1833 a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1834 sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1835 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1836 a_7565_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1837 a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1838 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1839 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1840 a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.20fF
C1841 a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.51fF
C1842 a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1843 a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1844 a_8657_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.98fF
C1845 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1846 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.19fF
C1847 sky130_fd_sc_hd__dfrbp_1_0[3]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1848 a_7153_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1849 a_6987_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1850 a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1851 a_5449_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1852 a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1853 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1854 a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1855 a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1856 a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1857 a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1858 a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1859 a_6541_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1860 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1861 a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1862 sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1863 a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1864 a_3333_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1865 a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1866 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1867 a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1868 a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.35fF
C1869 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.49fF
C1870 a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1871 a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1872 a_4425_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.98fF
C1873 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1874 a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.19fF
C1875 sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.32fF
C1876 a_2921_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.01fF
C1877 a_2755_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.03fF
C1878 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1879 a_1217_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.01fF
C1880 a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.11fF
C1881 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.23fF
C1882 a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.45fF
C1883 a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.79fF
C1884 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.50fF
C1885 a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.68fF
C1886 a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1887 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.16fF
C1888 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.04fF
C1889 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.42fF
C1890 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.13fF
C1891 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.09fF
C1892 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.08fF
C1893 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.30fF
C1894 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.51fF
C1895 a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB -0.44fF
C1896 a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.46fF
C1897 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.20fF
C1898 a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.40fF
C1899 a_193_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.98fF
C1900 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.58fF
C1901 a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 1.76fF
C1902 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 0.41fF
C1903 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 69.06fF
.end

