* NGSPICE file created from 20bitCounter_flat.ext - technology: sky130A

V1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB GND 1.8
V2 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK GND pulse(0V 1.8V clk_offset clk_risetime clk_falltime {clk_period/2} clk_period 0deg) 
V4 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND pwl(0.0us 1.8V, 0.090us 1.8V, 0.091us 0.0V, 0.100us 0.0V, 0.101us 1.8V)

.param clk_period=1us clk_offset={clk_period/2} clk_risetime=20ns clk_falltime={clk_risetime}
.func data_time(x) {clk_offset/2 + x*(clk_period/2)}

.tran 10ns {32*clk_period}
.save sky130_fd_sc_hd__dfrbp_1_0[0]/CLK sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B
.save sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[2]/Q sky130_fd_sc_hd__dfrbp_1_0[3]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[4]/Q sky130_fd_sc_hd__dfrbp_1_0[5]/Q sky130_fd_sc_hd__dfrbp_1_0[6]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[8]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[11]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[14]/Q sky130_fd_sc_hd__dfrbp_1_[15]/Q
.save sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[17]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/Q

.lib ~/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Top level circuit 20bitCounter_flat

X0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t222 a_41487_21# a_41474_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t104 a_20327_21# a_20314_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_9681_47# a_8491_47# a_9572_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t93 a_22268_47# a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t60 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15617_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_32379_47# a_31933_47# a_32283_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t12 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t59 a_9747_21# a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t11 a_30907_21# a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_24384_47# a_23469_47# a_24037_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_30167_47# a_29651_47# a_30072_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_19237_47# a_19071_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_805_47# a_761_289# a_639_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_38631_47# a_38115_47# a_38536_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t236 a_5515_21# a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t229 a_37255_21# a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_11219_47# a_10773_47# a_11123_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t7 a_28616_47# a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24081_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_19683_47# a_19237_47# a_19587_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 GND a_16095_21# a_16659_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t63 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t66 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 GND sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_17471_47# a_16955_47# a_17376_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t226 a_3399_21# a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t62 a_13979_21# a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t65 a_35139_21# a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t47 a_1283_21# a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 a_28791_21# a_28616_47# a_28970_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t101 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X43 a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1108_47# a_193_47# a_761_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t116 a_11863_21# a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X46 a_15005_47# a_14839_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t200 a_33023_21# a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X48 a_9572_47# a_8657_47# a_9225_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X49 GND sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 a_1283_21# a_1108_47# a_1462_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t34 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_17121_47# a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X53 a_38281_47# a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t8 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X54 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_4425_47# a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t78 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X56 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t33 a_7631_21# a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t153 a_39371_21# a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X58 GND a_37255_21# a_37819_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X59 a_36165_47# a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t94 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X60 a_2309_47# a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t95 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X61 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9269_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X62 a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X63 a_34049_47# a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t89 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X64 a_24384_47# a_23303_47# a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X65 a_41474_413# a_40397_47# a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X66 a_20314_413# a_19237_47# a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X67 a_30841_47# a_29651_47# a_30732_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X68 a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X69 a_26609_47# a_25419_47# a_26500_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X70 a_22268_47# a_21187_47# a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X71 GND a_11863_21# a_11797_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X72 a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X73 a_651_413# a_27_47# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 GND a_37255_21# a_37189_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X75 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 a_28616_47# a_27535_47# a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X77 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X78 a_35073_47# a_33883_47# a_34964_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X79 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X80 a_34617_289# a_34399_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X81 a_26500_47# a_25419_47# a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X82 GND a_16095_21# a_16029_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X83 a_32545_47# a_32501_289# a_32379_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X84 a_13457_289# a_13239_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X85 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t30 a_11341_289# a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 a_38849_289# a_38631_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X88 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t72 a_32501_289# a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X89 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X90 a_11385_47# a_11341_289# a_11219_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X92 a_30732_47# a_29817_47# a_30385_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t31 a_4993_289# a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 GND sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X95 a_26675_21# a_26500_47# a_26854_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t29 a_15573_289# a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t110 a_36733_289# a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t50 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X99 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t131 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t132 a_2877_289# a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X101 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26197_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X102 GND a_18211_21# a_18775_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_19587_47# a_19071_47# a_19492_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X105 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t96 a_13457_289# a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X107 GND sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t82 a_34617_289# a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t21 a_9225_289# a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X111 GND sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_805_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 GND sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 a_28051_47# a_27535_47# a_27956_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X115 a_3399_21# a_3224_47# a_3578_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t41 a_7109_289# a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t53 a_17689_289# a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t55 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t2 a_38849_289# a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X120 a_2755_47# a_2309_47# a_2659_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X121 a_25585_47# a_25419_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X122 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X123 GND a_39371_21# a_39935_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t217 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X125 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30429_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X126 a_32391_413# a_31767_47# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 GND a_3399_21# a_3963_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X128 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X129 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_30275_413# a_29651_47# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X131 a_32957_47# a_31767_47# a_32848_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X132 GND a_26675_21# a_27239_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X133 a_2309_47# a_2143_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t40 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_36623_413# a_35999_47# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 GND a_13979_21# a_13913_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 a_11797_47# a_10607_47# a_11688_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X138 a_37189_47# a_35999_47# a_37080_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X139 a_34507_413# a_33883_47# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 GND a_22443_21# a_22377_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X141 a_9115_413# a_8491_47# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 a_13457_289# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X143 a_34617_289# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X144 a_20261_47# a_19071_47# a_20152_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X145 a_11341_289# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X146 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 a_7109_289# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_32848_47# a_31933_47# a_32501_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X149 a_24037_289# a_23819_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X150 a_17689_289# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X151 a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t81 a_24559_21# a_24546_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_11688_47# a_10773_47# a_11341_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X154 a_15573_289# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X155 a_41421_47# a_40231_47# a_41312_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X156 a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X157 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t52 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 GND a_7631_21# a_7565_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X159 a_25935_47# a_25419_47# a_25840_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X160 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11385_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X162 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X164 a_20152_47# a_19237_47# a_19805_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t69 a_28791_21# a_28778_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 a_9225_289# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t44 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X167 GND a_28791_21# a_29355_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X168 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X169 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t24 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t17 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_16095_21# a_15920_47# a_16274_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_9225_289# a_9007_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X173 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t28 a_26675_21# a_26662_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X175 a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X176 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 a_15451_47# a_15005_47# a_15355_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X178 a_31933_47# a_31767_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X179 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 a_7153_47# a_7109_289# a_6987_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X182 GND sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X183 a_2659_47# a_2143_47# a_2564_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t139 a_16095_21# a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X185 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 a_21703_47# a_21353_47# a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X188 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32545_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t98 a_26500_47# a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X190 a_10773_47# a_10607_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 a_41312_47# a_40397_47# a_40965_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X192 a_10773_47# a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t22 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X193 a_36165_47# a_35999_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 a_40747_47# a_40397_47# a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 a_31933_47# a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t48 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X196 a_5340_47# a_4425_47# a_4993_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X197 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X198 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 a_37255_21# a_37080_47# a_37434_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X200 a_28051_47# a_27701_47# a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X201 a_6541_47# a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X202 a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41009_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X204 a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19849_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X207 a_2921_47# a_2877_289# a_2755_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_36611_47# a_36165_47# a_36515_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X209 a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X210 a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X211 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X212 GND sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_15005_47# a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X214 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 a_23819_47# a_23469_47# a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t122 a_18211_21# a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X217 GND a_1283_21# a_1847_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 a_12889_47# a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X221 GND a_24559_21# a_24493_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 a_22377_47# a_21187_47# a_22268_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X223 a_22430_413# a_21353_47# a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 a_8657_47# a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X226 a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X227 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X228 GND a_33023_21# a_32957_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 a_19237_47# a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X230 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t92 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 a_30385_289# a_30167_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X232 a_26662_413# a_25585_47# a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X233 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X234 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X235 a_19805_289# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t6 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X236 a_40965_289# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t99 a_30732_47# a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X238 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t76 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X239 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X240 a_24546_413# a_23469_47# a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 GND a_9747_21# a_9681_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t64 a_35139_21# a_35126_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 a_7565_47# a_6375_47# a_7456_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X245 a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X246 a_761_289# a_543_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X247 a_41009_47# a_40965_289# a_40843_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t199 a_33023_21# a_33010_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X249 a_22268_47# a_21353_47# a_21921_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X250 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X251 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t150 a_34964_47# a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t49 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X254 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X255 a_28778_413# a_27701_47# a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X256 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t23 a_11688_47# a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t112 a_32848_47# a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X259 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21965_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X260 a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X262 a_17567_47# a_17121_47# a_17471_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t5 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t214 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X265 a_15355_47# a_14839_47# a_15260_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t228 a_37255_21# a_37242_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X267 a_9269_47# a_9225_289# a_9103_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t220 a_41487_21# a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t147 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t91 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X271 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t27 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_12889_47# a_12723_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t26 a_26675_21# a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X274 a_26031_47# a_25585_47# a_25935_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X275 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t43 a_37080_47# a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t149 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X278 a_7456_47# a_6541_47# a_7109_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t119 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t75 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X281 a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t80 a_24559_21# a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X283 a_21353_47# a_21187_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t196 a_19805_289# a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 GND a_35139_21# a_35703_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X286 a_38727_47# a_38281_47# a_38631_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t38 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t202 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X289 a_22443_21# a_22268_47# a_22622_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X290 a_36515_47# a_35999_47# a_36420_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X291 a_40397_47# a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t143 a_22443_21# a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X293 GND a_13979_21# a_14543_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t134 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X295 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t68 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X297 GND a_30907_21# a_30841_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_3224_47# a_2143_47# a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X299 a_11231_413# a_10607_47# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X300 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2921_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 a_6541_47# a_6375_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X302 a_193_47# a_27_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 a_4883_413# a_4259_47# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X304 GND a_35139_21# a_35073_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X305 a_34964_47# a_33883_47# a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X306 a_1108_47# a_27_47# a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 a_7631_21# a_7456_47# a_7810_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 a_32848_47# a_31767_47# a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X309 a_32501_289# a_32283_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X310 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7153_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X311 a_15463_413# a_14839_47# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X312 a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X313 a_2767_413# a_2143_47# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X314 a_30732_47# a_29651_47# a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X315 a_11341_289# a_11123_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X316 a_39196_47# a_38115_47# a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 a_18036_47# a_16955_47# a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 a_13347_413# a_12723_47# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X319 a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X320 a_5340_47# a_4259_47# a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 a_35126_413# a_34049_47# a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X322 a_19695_413# a_19071_47# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_6999_413# a_6375_47# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X324 a_37080_47# a_35999_47# a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X325 a_19805_289# a_19587_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X326 a_17733_47# a_17689_289# a_17567_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X327 a_17579_413# a_16955_47# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 a_38739_413# a_38115_47# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X330 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t238 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t208 a_40965_289# a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X333 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X334 GND sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 a_30429_47# a_30385_289# a_30263_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X336 GND sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 a_38893_47# a_38849_289# a_38727_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 a_40965_289# a_40747_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X339 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X340 a_28147_47# a_27701_47# a_28051_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X341 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t70 a_26153_289# a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X343 a_11863_21# a_11688_47# a_12042_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X344 a_4993_289# a_4775_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X345 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t127 a_24037_289# a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X347 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X348 a_23469_47# a_23303_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X349 a_24559_21# a_24384_47# a_24738_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X350 a_543_47# a_27_47# a_448_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X351 GND a_20327_21# a_20891_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X352 a_15920_47# a_15005_47# a_15573_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X353 a_23915_47# a_23469_47# a_23819_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X354 a_21703_47# a_21187_47# a_21608_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X355 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t204 a_28269_289# a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X357 a_33023_21# a_32848_47# a_33202_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X358 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 GND a_24559_21# a_25123_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 GND sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X361 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 GND sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X363 a_8657_47# a_8491_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X364 a_25935_47# a_25585_47# a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X365 a_9747_21# a_9572_47# a_9926_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X366 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 GND a_20327_21# a_20261_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X368 a_543_47# a_193_47# a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X369 a_6891_47# a_6375_47# a_6796_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X370 a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X371 a_21921_289# a_21703_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X372 a_24037_289# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t87 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X373 a_19849_47# a_19805_289# a_19683_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 GND a_41487_21# a_41421_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X376 a_21921_289# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X377 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X378 GND a_5515_21# a_5449_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 a_3333_47# a_2143_47# a_3224_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t225 a_3399_21# a_3386_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X381 a_28269_289# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X382 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X383 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X384 GND a_28791_21# a_28725_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X385 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t61 a_13979_21# a_13966_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t46 a_1283_21# a_1270_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X388 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X389 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X390 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t54 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X391 a_26153_289# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X392 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t4 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t125 a_3224_47# a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_13979_21# a_13804_47# a_14158_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 a_7109_289# a_6891_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t32 a_7631_21# a_7618_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 a_13335_47# a_12889_47# a_13239_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X398 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X399 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X401 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t10 a_30907_21# a_30894_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t13 a_9572_47# a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X405 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t90 a_13804_47# a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X407 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 GND sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t137 a_1108_47# a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X410 a_5037_47# a_4993_289# a_4871_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t152 a_39371_21# a_39358_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t121 a_18211_21# a_18198_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t234 a_5515_21# a_5502_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X414 GND sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t102 a_20327_21# a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X417 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t19 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t203 a_7456_47# a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 a_28313_47# a_28269_289# a_28147_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X421 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t138 a_16095_21# a_16082_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X423 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38893_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X424 a_34049_47# a_33883_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X425 a_23819_47# a_23303_47# a_23724_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X426 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X427 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X428 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X429 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t108 a_39196_47# a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t109 a_18036_47# a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t117 a_5340_47# a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 a_35139_21# a_34964_47# a_35318_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X434 a_32283_47# a_31933_47# a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t58 a_9747_21# a_9734_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X436 a_34495_47# a_34049_47# a_34399_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X437 GND a_30907_21# a_31471_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X438 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t79 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17733_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X440 a_26500_47# a_25585_47# a_26153_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t20 a_15920_47# a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X442 a_32283_47# a_31767_47# a_32188_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X443 GND sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 GND a_9747_21# a_10311_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 a_30167_47# a_29817_47# a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X446 a_21353_47# a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t73 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X447 a_11123_47# a_10607_47# a_11028_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X448 a_36515_47# a_36165_47# a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X449 a_27701_47# a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X450 a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X452 a_9007_47# a_8491_47# a_8912_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X453 a_34399_47# a_34049_47# a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t67 a_28791_21# a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X456 a_25585_47# a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X457 a_3224_47# a_2309_47# a_2877_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X458 a_1270_413# a_193_47# a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 a_33010_413# a_31933_47# a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X460 a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X461 a_193_47# a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t85 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X462 a_23469_47# a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X463 a_13804_47# a_12723_47# a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X464 a_30894_413# a_29817_47# a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X465 a_29817_47# a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X466 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X467 a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X468 a_11688_47# a_10607_47# a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X469 GND a_18211_21# a_18145_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X470 a_5502_413# a_4425_47# a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X471 a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X472 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X473 a_5449_47# a_4259_47# a_5340_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X474 a_7456_47# a_6375_47# a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X475 a_16082_413# a_15005_47# a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X476 a_37242_413# a_36165_47# a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X477 a_3386_413# a_2309_47# a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X478 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X479 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X480 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X482 a_15920_47# a_14839_47# a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X483 a_28725_47# a_27535_47# a_28616_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X484 a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X486 a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X487 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 GND a_39371_21# a_39305_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X489 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 a_7618_413# a_6541_47# a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X491 a_13239_47# a_12723_47# a_13144_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t74 a_21921_289# a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X493 a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X494 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X495 a_36733_289# a_36515_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X496 a_9572_47# a_8491_47# a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X497 a_39358_413# a_38281_47# a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X498 a_18198_413# a_17121_47# a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 a_34661_47# a_34617_289# a_34495_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X501 a_15573_289# a_15355_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X502 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t106 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X504 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X505 a_41487_21# a_41312_47# a_41666_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_13501_47# a_13457_289# a_13335_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X507 a_40843_47# a_40397_47# a_40747_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X508 GND a_33023_21# a_33587_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t9 a_761_289# a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X510 a_34399_47# a_33883_47# a_34304_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X511 a_28616_47# a_27701_47# a_28269_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t36 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X513 a_20327_21# a_20152_47# a_20506_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X515 GND sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X516 GND a_11863_21# a_12427_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t18 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X518 GND a_41487_21# a_42051_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X519 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28313_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X520 a_37080_47# a_36165_47# a_36733_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X521 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X522 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t51 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X524 a_40397_47# a_40231_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X525 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X526 GND sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 a_21811_413# a_21187_47# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X528 a_5515_21# a_5340_47# a_5694_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X529 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5037_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X530 a_27701_47# a_27535_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X531 a_4871_47# a_4425_47# a_4775_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X532 a_40855_413# a_40231_47# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X533 a_18145_47# a_16955_47# a_18036_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X534 a_17689_289# a_17471_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X535 GND a_5515_21# a_6079_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 a_9103_47# a_8657_47# a_9007_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X537 a_26043_413# a_25419_47# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 a_23927_413# a_23303_47# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 a_41312_47# a_40231_47# a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X540 a_20152_47# a_19071_47# a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X541 a_4425_47# a_4259_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 a_13913_47# a_12723_47# a_13804_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X543 a_39305_47# a_38115_47# a_39196_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X544 a_28159_413# a_27535_47# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X545 a_36777_47# a_36733_289# a_36611_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X546 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X547 a_18036_47# a_17121_47# a_17689_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t216 a_30385_289# a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X549 a_15617_47# a_15573_289# a_15451_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t115 a_11863_21# a_11850_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X551 a_34964_47# a_34049_47# a_34617_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X552 a_26153_289# a_25935_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X553 a_40747_47# a_40231_47# a_40652_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X554 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X555 a_639_47# a_193_47# a_543_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X556 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X557 GND a_1283_21# a_1217_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 a_24081_47# a_24037_289# a_23915_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X559 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X560 a_13804_47# a_12889_47# a_13457_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X561 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_21799_47# a_21353_47# a_21703_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X563 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34661_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X564 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X565 a_39196_47# a_38281_47# a_38849_289# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X566 a_30907_21# a_30732_47# a_31086_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X567 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13501_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 a_39371_21# a_39196_47# a_39550_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X569 a_30263_47# a_29817_47# a_30167_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X570 GND a_22443_21# a_23007_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t88 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_2877_289# a_2659_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X575 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t71 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X576 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X577 a_18211_21# a_18036_47# a_18390_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X578 a_6891_47# a_6541_47# a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X579 a_11123_47# a_10773_47# a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X580 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X583 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X584 a_6987_47# a_6541_47# a_6891_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X585 a_17471_47# a_17121_47# a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 a_38631_47# a_38281_47# a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X587 a_29817_47# a_29651_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 GND sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X589 a_4775_47# a_4425_47# a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X590 a_4775_47# a_4259_47# a_4680_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X591 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t77 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X593 a_15355_47# a_15005_47# a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 a_2659_47# a_2309_47# a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X595 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t14 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_38281_47# a_38115_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 GND a_7631_21# a_8195_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X598 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t15 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 a_9007_47# a_8657_47# a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X600 a_13239_47# a_12889_47# a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X601 GND sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X602 a_17121_47# a_16955_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 GND sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X604 a_11850_413# a_10773_47# a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 a_19587_47# a_19237_47# a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 a_2877_289# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t84 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X607 a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X608 a_16029_47# a_14839_47# a_15920_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X609 a_761_289# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X610 a_32501_289# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t16 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X611 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t35 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X612 GND a_26675_21# a_26609_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X613 a_24493_47# a_23303_47# a_24384_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X614 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X615 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X616 a_30385_289# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t151 a_20152_47# a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X618 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t25 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t83 a_41312_47# a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X620 a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X621 a_13966_413# a_12889_47# a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 a_38849_289# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t56 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X623 a_21965_47# a_21921_289# a_21799_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_4993_289# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t215 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X625 a_9734_413# a_8657_47# a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X626 a_28269_289# a_28051_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X627 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X628 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 a_36733_289# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t141 a_22443_21# a_22430_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t224 a_24384_47# a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 GND a_3399_21# a_3333_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X633 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X634 a_26197_47# a_26153_289# a_26031_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X635 a_1217_47# a_27_47# a_1108_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X636 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 GND sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36777_47# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X638 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X639 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
R0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1612 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t84 225.592
R1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t205 225.592
R2 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n52 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t209 225.592
R3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t56 225.592
R4 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t219 225.592
R5 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n301 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t111 225.592
R6 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n384 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t16 225.592
R7 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t223 225.592
R8 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t42 225.592
R9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n633 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t105 225.592
R10 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t87 225.592
R11 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n799 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t212 225.592
R12 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n882 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t6 225.592
R13 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n965 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t197 225.592
R14 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1048 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t0 225.592
R15 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t39 225.592
R16 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t126 225.592
R17 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t44 225.592
R18 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t86 225.592
R19 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t215 225.592
R20 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t225 119.607
R21 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t46 119.607
R22 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t222 119.607
R23 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t152 119.607
R24 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t228 119.607
R25 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t64 119.607
R26 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t199 119.607
R27 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t10 119.607
R28 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t69 119.607
R29 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t28 119.607
R30 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t81 119.607
R31 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t141 119.607
R32 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t104 119.607
R33 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n951 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t121 119.607
R34 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1034 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t138 119.607
R35 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t61 119.607
R36 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t115 119.607
R37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t58 119.607
R38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t32 119.607
R39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t234 119.607
R40 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t132 93.809
R41 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t9 93.809
R42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n59 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t208 93.809
R43 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t2 93.809
R44 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t110 93.809
R45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t82 93.809
R46 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t72 93.809
R47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t216 93.809
R48 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n557 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t204 93.809
R49 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t70 93.809
R50 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t127 93.809
R51 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t74 93.809
R52 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t196 93.809
R53 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n972 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t53 93.809
R54 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1055 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t29 93.809
R55 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t96 93.809
R56 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t30 93.809
R57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t21 93.809
R58 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t41 93.809
R59 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t31 93.809
R60 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t4 85.217
R61 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t130 85.217
R62 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n76 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t25 85.217
R63 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t237 85.217
R64 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t54 85.217
R65 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n325 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t49 85.217
R66 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t92 85.217
R67 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t76 85.217
R68 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n574 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t100 85.217
R69 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n657 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t52 85.217
R70 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n740 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t107 85.217
R71 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n823 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t35 85.217
R72 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n906 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t19 85.217
R73 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n989 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t37 85.217
R74 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1072 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t133 85.217
R75 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t213 85.217
R76 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t146 85.217
R77 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t118 85.217
R78 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t148 85.217
R79 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t201 85.217
R80 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t117 68.011
R81 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t203 68.011
R82 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t13 68.011
R83 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t23 68.011
R84 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t90 68.011
R85 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1026 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t20 68.011
R86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n943 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t109 68.011
R87 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t151 68.011
R88 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n777 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t93 68.011
R89 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n694 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t224 68.011
R90 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t98 68.011
R91 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t7 68.011
R92 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t99 68.011
R93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t112 68.011
R94 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t150 68.011
R95 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t43 68.011
R96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t108 68.011
R97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n30 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t83 68.011
R98 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t137 68.011
R99 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t125 68.011
R100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t187 63.321
R101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t159 63.321
R102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t156 63.321
R103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t167 63.321
R104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n59 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t176 63.321
R105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t191 63.321
R106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t180 63.321
R107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t164 63.321
R108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t188 63.321
R109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t160 63.321
R110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t185 63.321
R111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t173 63.321
R112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t193 63.321
R113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t175 63.321
R114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t195 63.321
R115 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t174 63.321
R116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n557 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t168 63.321
R117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t179 63.321
R118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t171 63.321
R119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t178 63.321
R120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t170 63.321
R121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t177 63.321
R122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t169 63.321
R123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t192 63.321
R124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t172 63.321
R125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t190 63.321
R126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n972 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t181 63.321
R127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n951 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t163 63.321
R128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1055 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t189 63.321
R129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1034 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t161 63.321
R130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t186 63.321
R131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t157 63.321
R132 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t183 63.321
R133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t165 63.321
R134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t184 63.321
R135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t158 63.321
R136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t182 63.321
R137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t166 63.321
R138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t194 63.321
R139 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t162 63.321
R140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t47 61.575
R141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n16 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t220 61.575
R142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t153 61.575
R143 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t229 61.575
R144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t65 61.575
R145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t200 61.575
R146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t11 61.575
R147 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t67 61.575
R148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n595 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t26 61.575
R149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t80 61.575
R150 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t143 61.575
R151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t102 61.575
R152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n927 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t122 61.575
R153 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1010 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t139 61.575
R154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1093 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t62 61.575
R155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t116 61.575
R156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t59 61.575
R157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t33 61.575
R158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t236 61.575
R159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t226 61.562
R160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1493 50.786
R161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1621 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1620 50.667
R162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1617 50.667
R163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1614 50.667
R164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1610 50.667
R165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1607 50.667
R166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1603 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1602 50.667
R167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1600 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1599 50.667
R168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1596 50.667
R169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1593 50.667
R170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1590 50.667
R171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1586 50.667
R172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1583 50.667
R173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1581 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1580 50.667
R174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1575 50.667
R175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1572 50.667
R176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1569 50.667
R177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1565 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1564 50.667
R178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1562 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1561 50.667
R179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1558 50.667
R180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1555 50.667
R181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1548 50.667
R182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1545 50.667
R183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1540 50.667
R184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1537 50.667
R185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1534 50.667
R186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1531 50.667
R187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1527 50.667
R188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1524 50.667
R189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1519 50.667
R190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1516 50.667
R191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1513 50.667
R192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1510 50.667
R193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1507 50.667
R194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1503 50.667
R195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1500 50.667
R196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1497 50.667
R197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n27 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n26 50.667
R198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n24 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n23 50.667
R199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n34 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n33 50.667
R200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n36 50.667
R201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n41 50.667
R202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n44 50.667
R203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n48 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n47 50.667
R204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n51 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n50 50.667
R205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n55 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n54 50.667
R206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n58 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n57 50.667
R207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n63 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n62 50.667
R208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n66 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n65 50.667
R209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n69 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n68 50.667
R210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n72 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n71 50.667
R211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n75 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n74 50.667
R212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n79 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n78 50.667
R213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n82 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n81 50.667
R214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n85 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n84 50.667
R215 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n90 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n89 50.667
R216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n92 50.667
R217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n95 50.667
R218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n100 50.667
R219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n103 50.667
R220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n106 50.667
R221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n109 50.667
R222 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n116 50.667
R223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n119 50.667
R224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n124 50.667
R225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n127 50.667
R226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n130 50.667
R227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n133 50.667
R228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n137 50.667
R229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n140 50.667
R230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n145 50.667
R231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n148 50.667
R232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n151 50.667
R233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n154 50.667
R234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n157 50.667
R235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n161 50.667
R236 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n164 50.667
R237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n167 50.667
R238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n172 50.667
R239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n175 50.667
R240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n178 50.667
R241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n183 50.667
R242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n186 50.667
R243 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n189 50.667
R244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n192 50.667
R245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n199 50.667
R246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n202 50.667
R247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n207 50.667
R248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n210 50.667
R249 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n213 50.667
R250 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n216 50.667
R251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n220 50.667
R252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n223 50.667
R253 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n228 50.667
R254 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n231 50.667
R255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n234 50.667
R256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n237 50.667
R257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n240 50.667
R258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n244 50.667
R259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n247 50.667
R260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n250 50.667
R261 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n255 50.667
R262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n258 50.667
R263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n261 50.667
R264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n266 50.667
R265 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n269 50.667
R266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n272 50.667
R267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n275 50.667
R268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n282 50.667
R269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n285 50.667
R270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n290 50.667
R271 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n293 50.667
R272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n296 50.667
R273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n299 50.667
R274 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n303 50.667
R275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n306 50.667
R276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n311 50.667
R277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n314 50.667
R278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n317 50.667
R279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n320 50.667
R280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n323 50.667
R281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n327 50.667
R282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n330 50.667
R283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n333 50.667
R284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n338 50.667
R285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n341 50.667
R286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n344 50.667
R287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n349 50.667
R288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n352 50.667
R289 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n355 50.667
R290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n358 50.667
R291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n365 50.667
R292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n368 50.667
R293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n373 50.667
R294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n376 50.667
R295 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n379 50.667
R296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n382 50.667
R297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n386 50.667
R298 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n389 50.667
R299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n394 50.667
R300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n397 50.667
R301 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n400 50.667
R302 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n403 50.667
R303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n406 50.667
R304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n410 50.667
R305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n413 50.667
R306 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n416 50.667
R307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n421 50.667
R308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n424 50.667
R309 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n427 50.667
R310 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n432 50.667
R311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n435 50.667
R312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n438 50.667
R313 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n441 50.667
R314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n448 50.667
R315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n451 50.667
R316 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n456 50.667
R317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n459 50.667
R318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n462 50.667
R319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n465 50.667
R320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n469 50.667
R321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n472 50.667
R322 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n477 50.667
R323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n480 50.667
R324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n483 50.667
R325 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n486 50.667
R326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n489 50.667
R327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n493 50.667
R328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n496 50.667
R329 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n499 50.667
R330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n504 50.667
R331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n507 50.667
R332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n510 50.667
R333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n515 50.667
R334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n518 50.667
R335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n521 50.667
R336 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n524 50.667
R337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n531 50.667
R338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n534 50.667
R339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n539 50.667
R340 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n542 50.667
R341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n545 50.667
R342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n548 50.667
R343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n552 50.667
R344 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n555 50.667
R345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n560 50.667
R346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n563 50.667
R347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n566 50.667
R348 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n569 50.667
R349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n572 50.667
R350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n576 50.667
R351 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n579 50.667
R352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n582 50.667
R353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n587 50.667
R354 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n590 50.667
R355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n593 50.667
R356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n598 50.667
R357 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n601 50.667
R358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n604 50.667
R359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n607 50.667
R360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n614 50.667
R361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n617 50.667
R362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n622 50.667
R363 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n625 50.667
R364 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n628 50.667
R365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n631 50.667
R366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n636 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n635 50.667
R367 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n638 50.667
R368 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n643 50.667
R369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n646 50.667
R370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n649 50.667
R371 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n652 50.667
R372 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n655 50.667
R373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n660 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n659 50.667
R374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n662 50.667
R375 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n665 50.667
R376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n670 50.667
R377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n673 50.667
R378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n676 50.667
R379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n681 50.667
R380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n684 50.667
R381 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n687 50.667
R382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n690 50.667
R383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n697 50.667
R384 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n700 50.667
R385 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n705 50.667
R386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n708 50.667
R387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n711 50.667
R388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n714 50.667
R389 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n718 50.667
R390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n721 50.667
R391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n726 50.667
R392 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n729 50.667
R393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n732 50.667
R394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n735 50.667
R395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n738 50.667
R396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n742 50.667
R397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n745 50.667
R398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n748 50.667
R399 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n753 50.667
R400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n756 50.667
R401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n759 50.667
R402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n764 50.667
R403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n767 50.667
R404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n770 50.667
R405 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n773 50.667
R406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n780 50.667
R407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n783 50.667
R408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n788 50.667
R409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n791 50.667
R410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n794 50.667
R411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n797 50.667
R412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n801 50.667
R413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n804 50.667
R414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n809 50.667
R415 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n812 50.667
R416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n815 50.667
R417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n818 50.667
R418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n821 50.667
R419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n825 50.667
R420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n828 50.667
R421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n831 50.667
R422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n836 50.667
R423 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n839 50.667
R424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n842 50.667
R425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n847 50.667
R426 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n850 50.667
R427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n853 50.667
R428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n856 50.667
R429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n863 50.667
R430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n866 50.667
R431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n871 50.667
R432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n874 50.667
R433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n877 50.667
R434 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n880 50.667
R435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n884 50.667
R436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n887 50.667
R437 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n892 50.667
R438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n896 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n895 50.667
R439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n898 50.667
R440 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n902 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n901 50.667
R441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n905 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n904 50.667
R442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n909 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n908 50.667
R443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n912 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n911 50.667
R444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n915 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n914 50.667
R445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n920 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n919 50.667
R446 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n923 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n922 50.667
R447 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n926 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n925 50.667
R448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n930 50.667
R449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n934 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n933 50.667
R450 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n937 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n936 50.667
R451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n940 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n939 50.667
R452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n947 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n946 50.667
R453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n950 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n949 50.667
R454 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n954 50.667
R455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n958 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n957 50.667
R456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n961 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n960 50.667
R457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n964 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n963 50.667
R458 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n967 50.667
R459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n970 50.667
R460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n976 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n975 50.667
R461 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n979 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n978 50.667
R462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n982 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n981 50.667
R463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n985 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n984 50.667
R464 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n988 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n987 50.667
R465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n992 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n991 50.667
R466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n994 50.667
R467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n998 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n997 50.667
R468 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1003 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1002 50.667
R469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1006 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1005 50.667
R470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1009 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1008 50.667
R471 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1014 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1013 50.667
R472 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1017 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1016 50.667
R473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1020 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1019 50.667
R474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1023 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1022 50.667
R475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1030 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1029 50.667
R476 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1033 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1032 50.667
R477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1038 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1037 50.667
R478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1041 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1040 50.667
R479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1044 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1043 50.667
R480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1047 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1046 50.667
R481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1051 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1050 50.667
R482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1054 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1053 50.667
R483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1059 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1058 50.667
R484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1061 50.667
R485 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1065 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1064 50.667
R486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1068 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1067 50.667
R487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1071 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1070 50.667
R488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1075 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1074 50.667
R489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1078 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1077 50.667
R490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1081 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1080 50.667
R491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1086 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1085 50.667
R492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1089 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1088 50.667
R493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1092 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1091 50.667
R494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1097 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1096 50.667
R495 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1099 50.667
R496 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1102 50.667
R497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1105 50.667
R498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1112 50.667
R499 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1115 50.667
R500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1120 50.667
R501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1123 50.667
R502 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1126 50.667
R503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1129 50.667
R504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1133 50.667
R505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1136 50.667
R506 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1141 50.667
R507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1144 50.667
R508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1147 50.667
R509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1150 50.667
R510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1153 50.667
R511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1157 50.667
R512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1160 50.667
R513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1163 50.667
R514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1168 50.667
R515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1171 50.667
R516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1174 50.667
R517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1179 50.667
R518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1182 50.667
R519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1185 50.667
R520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1188 50.667
R521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1195 50.667
R522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1198 50.667
R523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1203 50.667
R524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1206 50.667
R525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1209 50.667
R526 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1212 50.667
R527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1216 50.667
R528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1219 50.667
R529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1224 50.667
R530 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1227 50.667
R531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1230 50.667
R532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1233 50.667
R533 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1236 50.667
R534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1240 50.667
R535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1243 50.667
R536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1246 50.667
R537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1251 50.667
R538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1254 50.667
R539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1257 50.667
R540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1262 50.667
R541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1265 50.667
R542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1268 50.667
R543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1271 50.667
R544 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1278 50.667
R545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1281 50.667
R546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1286 50.667
R547 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1289 50.667
R548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1292 50.667
R549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1295 50.667
R550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1299 50.667
R551 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1302 50.667
R552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1307 50.667
R553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1310 50.667
R554 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1313 50.667
R555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1316 50.667
R556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1319 50.667
R557 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1323 50.667
R558 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1326 50.667
R559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1329 50.667
R560 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1334 50.667
R561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1337 50.667
R562 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1340 50.667
R563 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1345 50.667
R564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1348 50.667
R565 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1351 50.667
R566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1354 50.667
R567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1361 50.667
R568 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1364 50.667
R569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1369 50.667
R570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1372 50.667
R571 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1375 50.667
R572 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1378 50.667
R573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1382 50.667
R574 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1385 50.667
R575 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1390 50.667
R576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1393 50.667
R577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1396 50.667
R578 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1399 50.667
R579 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1402 50.667
R580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1406 50.667
R581 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1409 50.667
R582 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1412 50.667
R583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1417 50.667
R584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1420 50.667
R585 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1423 50.667
R586 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1428 50.667
R587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1431 50.667
R588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1434 50.667
R589 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1437 50.667
R590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1444 50.667
R591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1447 50.667
R592 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1452 50.667
R593 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1455 50.667
R594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1458 50.667
R595 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1461 50.667
R596 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1465 50.667
R597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1468 50.667
R598 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1473 50.667
R599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1476 50.667
R600 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1479 50.667
R601 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1482 50.667
R602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1485 50.667
R603 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1629 50.667
R604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t95 41.554
R605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t131 41.554
R606 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t85 41.554
R607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t217 41.554
R608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t1 41.554
R609 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t238 41.554
R610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t8 41.554
R611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t55 41.554
R612 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t94 41.554
R613 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t50 41.554
R614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t89 41.554
R615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t91 41.554
R616 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t48 41.554
R617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t75 41.554
R618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t232 41.554
R619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t101 41.554
R620 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t136 41.554
R621 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t51 41.554
R622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t97 41.554
R623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t106 41.554
R624 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t145 41.554
R625 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t36 41.554
R626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t73 41.554
R627 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t18 41.554
R628 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n916 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t231 41.554
R629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n916 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t38 41.554
R630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n999 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t135 41.554
R631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n999 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t134 41.554
R632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1082 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t144 41.554
R633 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1082 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t214 41.554
R634 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t239 41.554
R635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t147 41.554
R636 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t22 41.554
R637 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t119 41.554
R638 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t233 41.554
R639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t149 41.554
R640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t210 41.554
R641 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t202 41.554
R642 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t78 41.554
R643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t5 41.554
R644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1655 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1654 40.334
R645 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t211 30.569
R646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n16 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t24 30.569
R647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t129 30.569
R648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t15 30.569
R649 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t71 30.569
R650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t113 30.569
R651 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t57 30.569
R652 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t155 30.569
R653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n595 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t218 30.569
R654 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t206 30.569
R655 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t120 30.569
R656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t17 30.569
R657 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n927 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t124 30.569
R658 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1010 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t40 30.569
R659 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1093 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t88 30.569
R660 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t207 30.569
R661 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t128 30.569
R662 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t77 30.569
R663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t14 30.569
R664 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t235 29.315
R665 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t34 29.315
R666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t60 29.315
R667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t114 29.315
R668 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t63 29.315
R669 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1024 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t140 29.315
R670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n941 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t123 29.315
R671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n858 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t103 29.315
R672 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n775 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t142 29.315
R673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n692 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t79 29.315
R674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n609 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t27 29.315
R675 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n526 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t68 29.315
R676 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t12 29.315
R677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t198 29.315
R678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t66 29.315
R679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t230 29.315
R680 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t154 29.315
R681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n28 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t221 29.315
R682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t45 29.315
R683 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t227 29.315
R684 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1652 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t3 29.055
R685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n21 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n20 28.517
R686 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1566 27.22
R687 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n19 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n16 27.22
R688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n98 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n97 27.22
R689 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n180 27.22
R690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n263 27.22
R691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n346 27.22
R692 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n429 27.22
R693 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n512 27.22
R694 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n596 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n595 27.22
R695 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n678 27.22
R696 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n762 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n761 27.22
R697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n845 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n844 27.22
R698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n928 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n927 27.22
R699 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1011 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1010 27.22
R700 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1094 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1093 27.22
R701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1176 27.22
R702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1259 27.22
R703 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1342 27.22
R704 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1426 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1425 27.22
R705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1654 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1651 25.815
R706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1578 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1577 22.842
R707 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1495 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1494 22.842
R708 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n87 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n86 22.842
R709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n169 22.842
R710 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n253 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n252 22.842
R711 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n336 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n335 22.842
R712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n418 22.842
R713 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n502 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n501 22.842
R714 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n585 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n584 22.842
R715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n668 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n667 22.842
R716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n751 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n750 22.842
R717 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n834 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n833 22.842
R718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n917 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n916 22.842
R719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1000 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n999 22.842
R720 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1083 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1082 22.842
R721 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1165 22.842
R722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1249 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1248 22.842
R723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1331 22.842
R724 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1415 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1414 22.842
R725 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n10 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n0 22.842
R726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1632 21.896
R727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1542 21.896
R728 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n38 21.896
R729 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n121 21.896
R730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n204 21.896
R731 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n287 21.896
R732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n371 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n370 21.896
R733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n454 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n453 21.896
R734 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n536 21.896
R735 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n620 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n619 21.896
R736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n703 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n702 21.896
R737 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n786 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n785 21.896
R738 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n868 21.896
R739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n952 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n951 21.896
R740 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1035 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1034 21.896
R741 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1117 21.896
R742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1200 21.896
R743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1283 21.896
R744 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1367 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1366 21.896
R745 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1450 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1449 21.896
R746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1604 20.254
R747 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1521 20.254
R748 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n60 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n59 20.254
R749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n143 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n142 20.254
R750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n225 20.254
R751 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n309 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n308 20.254
R752 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n392 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n391 20.254
R753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n474 20.254
R754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n558 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n557 20.254
R755 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n641 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n640 20.254
R756 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n724 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n723 20.254
R757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n807 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n806 20.254
R758 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n890 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n889 20.254
R759 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n973 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n972 20.254
R760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1056 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1055 20.254
R761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1139 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1138 20.254
R762 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1222 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1221 20.254
R763 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1304 20.254
R764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1387 20.254
R765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1471 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1470 20.254
R766 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1637 15.167
R767 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n7 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n5 15.167
R768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n7 15.167
R769 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n14 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n12 15.167
R770 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n14 15.167
R771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1648 15.167
R772 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1646 15.167
R773 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n12 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n10 14.837
R774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n19 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n18 13.683
R775 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1651 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1650 13.683
R776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1634 13.024
R777 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n3 12.035
R778 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1631 7.5
R779 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1643 7.5
R780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1552 7.5
R781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1551 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1550 7.5
R782 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n31 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n30 7.5
R783 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n29 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n28 7.5
R784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n113 7.5
R785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n111 7.5
R786 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n196 7.5
R787 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n194 7.5
R788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n279 7.5
R789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n277 7.5
R790 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n363 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n362 7.5
R791 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n360 7.5
R792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n446 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n445 7.5
R793 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n443 7.5
R794 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n528 7.5
R795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n526 7.5
R796 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n612 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n611 7.5
R797 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n609 7.5
R798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n695 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n694 7.5
R799 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n693 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n692 7.5
R800 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n778 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n777 7.5
R801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n775 7.5
R802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n861 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n860 7.5
R803 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n859 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n858 7.5
R804 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n944 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n943 7.5
R805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n942 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n941 7.5
R806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1027 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1026 7.5
R807 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1025 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1024 7.5
R808 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1109 7.5
R809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1107 7.5
R810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1192 7.5
R811 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1190 7.5
R812 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1275 7.5
R813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1274 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1273 7.5
R814 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1358 7.5
R815 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1357 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1356 7.5
R816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1441 7.5
R817 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1440 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1439 7.5
R818 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1496 7.147
R819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1499 7.147
R820 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1502 7.147
R821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1506 7.147
R822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1509 7.147
R823 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1512 7.147
R824 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1515 7.147
R825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1518 7.147
R826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1523 7.147
R827 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1526 7.147
R828 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1530 7.147
R829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1533 7.147
R830 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1536 7.147
R831 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1539 7.147
R832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1544 7.147
R833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1547 7.147
R834 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1554 7.147
R835 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1558 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1557 7.147
R836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1560 7.147
R837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1563 7.147
R838 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1568 7.147
R839 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1572 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1571 7.147
R840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1575 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1574 7.147
R841 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1579 7.147
R842 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1582 7.147
R843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1586 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1585 7.147
R844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1589 7.147
R845 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1593 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1592 7.147
R846 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1596 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1595 7.147
R847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1598 7.147
R848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1601 7.147
R849 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1606 7.147
R850 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1609 7.147
R851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1613 7.147
R852 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1616 7.147
R853 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1620 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1619 7.147
R854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1634 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1633 7.147
R855 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1637 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1636 7.147
R856 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1638 7.147
R857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1642 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1641 7.147
R858 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n26 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n25 7.147
R859 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n23 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n22 7.147
R860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n18 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n17 7.147
R861 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n33 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n32 7.147
R862 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n108 7.147
R863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n105 7.147
R864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n102 7.147
R865 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n99 7.147
R866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n95 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n94 7.147
R867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n92 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n91 7.147
R868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n89 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n88 7.147
R869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n84 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n83 7.147
R870 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n81 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n80 7.147
R871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n78 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n77 7.147
R872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n74 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n73 7.147
R873 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n71 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n70 7.147
R874 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n68 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n67 7.147
R875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n65 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n64 7.147
R876 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n62 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n61 7.147
R877 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n56 7.147
R878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n54 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n53 7.147
R879 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n50 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n49 7.147
R880 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n46 7.147
R881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n44 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n43 7.147
R882 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n41 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n40 7.147
R883 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n36 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n35 7.147
R884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n115 7.147
R885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n191 7.147
R886 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n188 7.147
R887 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n185 7.147
R888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n182 7.147
R889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n177 7.147
R890 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n174 7.147
R891 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n171 7.147
R892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n166 7.147
R893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n163 7.147
R894 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n160 7.147
R895 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n156 7.147
R896 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n153 7.147
R897 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n150 7.147
R898 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n147 7.147
R899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n144 7.147
R900 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n139 7.147
R901 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n136 7.147
R902 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n132 7.147
R903 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n129 7.147
R904 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n126 7.147
R905 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n123 7.147
R906 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n118 7.147
R907 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n198 7.147
R908 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n274 7.147
R909 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n271 7.147
R910 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n268 7.147
R911 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n265 7.147
R912 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n261 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n260 7.147
R913 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n257 7.147
R914 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n254 7.147
R915 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n250 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n249 7.147
R916 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n246 7.147
R917 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n243 7.147
R918 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n239 7.147
R919 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n236 7.147
R920 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n233 7.147
R921 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n230 7.147
R922 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n227 7.147
R923 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n222 7.147
R924 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n219 7.147
R925 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n215 7.147
R926 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n212 7.147
R927 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n209 7.147
R928 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n206 7.147
R929 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n201 7.147
R930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n281 7.147
R931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n357 7.147
R932 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n354 7.147
R933 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n351 7.147
R934 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n348 7.147
R935 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n344 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n343 7.147
R936 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n340 7.147
R937 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n337 7.147
R938 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n332 7.147
R939 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n329 7.147
R940 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n326 7.147
R941 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n322 7.147
R942 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n319 7.147
R943 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n316 7.147
R944 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n313 7.147
R945 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n310 7.147
R946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n306 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n305 7.147
R947 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n302 7.147
R948 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n298 7.147
R949 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n295 7.147
R950 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n292 7.147
R951 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n289 7.147
R952 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n284 7.147
R953 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n364 7.147
R954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n440 7.147
R955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n437 7.147
R956 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n434 7.147
R957 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n431 7.147
R958 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n426 7.147
R959 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n423 7.147
R960 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n420 7.147
R961 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n415 7.147
R962 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n412 7.147
R963 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n409 7.147
R964 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n405 7.147
R965 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n402 7.147
R966 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n399 7.147
R967 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n396 7.147
R968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n393 7.147
R969 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n389 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n388 7.147
R970 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n385 7.147
R971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n381 7.147
R972 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n378 7.147
R973 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n375 7.147
R974 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n372 7.147
R975 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n368 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n367 7.147
R976 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n447 7.147
R977 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n523 7.147
R978 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n520 7.147
R979 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n517 7.147
R980 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n514 7.147
R981 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n509 7.147
R982 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n506 7.147
R983 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n503 7.147
R984 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n499 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n498 7.147
R985 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n496 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n495 7.147
R986 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n492 7.147
R987 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n488 7.147
R988 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n485 7.147
R989 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n482 7.147
R990 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n479 7.147
R991 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n476 7.147
R992 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n472 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n471 7.147
R993 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n468 7.147
R994 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n464 7.147
R995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n461 7.147
R996 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n458 7.147
R997 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n455 7.147
R998 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n450 7.147
R999 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n530 7.147
R1000 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n606 7.147
R1001 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n603 7.147
R1002 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n601 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n600 7.147
R1003 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n598 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n597 7.147
R1004 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n593 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n592 7.147
R1005 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n589 7.147
R1006 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n586 7.147
R1007 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n582 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n581 7.147
R1008 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n579 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n578 7.147
R1009 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n575 7.147
R1010 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n572 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n571 7.147
R1011 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n568 7.147
R1012 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n565 7.147
R1013 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n563 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n562 7.147
R1014 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n560 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n559 7.147
R1015 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n554 7.147
R1016 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n551 7.147
R1017 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n547 7.147
R1018 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n544 7.147
R1019 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n541 7.147
R1020 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n538 7.147
R1021 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n533 7.147
R1022 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n613 7.147
R1023 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n689 7.147
R1024 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n687 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n686 7.147
R1025 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n684 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n683 7.147
R1026 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n680 7.147
R1027 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n676 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n675 7.147
R1028 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n672 7.147
R1029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n669 7.147
R1030 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n665 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n664 7.147
R1031 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n662 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n661 7.147
R1032 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n659 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n658 7.147
R1033 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n655 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n654 7.147
R1034 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n652 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n651 7.147
R1035 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n649 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n648 7.147
R1036 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n645 7.147
R1037 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n642 7.147
R1038 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n638 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n637 7.147
R1039 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n634 7.147
R1040 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n630 7.147
R1041 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n628 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n627 7.147
R1042 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n625 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n624 7.147
R1043 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n621 7.147
R1044 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n616 7.147
R1045 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n696 7.147
R1046 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n773 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n772 7.147
R1047 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n770 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n769 7.147
R1048 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n767 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n766 7.147
R1049 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n763 7.147
R1050 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n759 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n758 7.147
R1051 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n756 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n755 7.147
R1052 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n752 7.147
R1053 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n748 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n747 7.147
R1054 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n745 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n744 7.147
R1055 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n741 7.147
R1056 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n738 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n737 7.147
R1057 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n735 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n734 7.147
R1058 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n731 7.147
R1059 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n729 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n728 7.147
R1060 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n725 7.147
R1061 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n721 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n720 7.147
R1062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n717 7.147
R1063 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n714 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n713 7.147
R1064 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n711 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n710 7.147
R1065 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n708 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n707 7.147
R1066 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n704 7.147
R1067 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n700 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n699 7.147
R1068 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n779 7.147
R1069 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n856 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n855 7.147
R1070 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n853 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n852 7.147
R1071 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n850 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n849 7.147
R1072 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n846 7.147
R1073 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n842 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n841 7.147
R1074 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n839 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n838 7.147
R1075 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n835 7.147
R1076 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n831 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n830 7.147
R1077 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n828 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n827 7.147
R1078 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n824 7.147
R1079 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n820 7.147
R1080 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n818 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n817 7.147
R1081 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n815 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n814 7.147
R1082 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n812 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n811 7.147
R1083 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n808 7.147
R1084 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n804 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n803 7.147
R1085 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n800 7.147
R1086 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n797 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n796 7.147
R1087 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n794 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n793 7.147
R1088 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n791 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n790 7.147
R1089 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n787 7.147
R1090 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n783 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n782 7.147
R1091 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n862 7.147
R1092 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n939 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n938 7.147
R1093 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n936 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n935 7.147
R1094 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n933 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n932 7.147
R1095 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n929 7.147
R1096 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n925 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n924 7.147
R1097 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n922 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n921 7.147
R1098 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n919 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n918 7.147
R1099 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n914 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n913 7.147
R1100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n911 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n910 7.147
R1101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n908 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n907 7.147
R1102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n904 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n903 7.147
R1103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n901 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n900 7.147
R1104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n898 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n897 7.147
R1105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n895 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n894 7.147
R1106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n891 7.147
R1107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n887 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n886 7.147
R1108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n883 7.147
R1109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n880 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n879 7.147
R1110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n877 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n876 7.147
R1111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n874 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n873 7.147
R1112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n870 7.147
R1113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n865 7.147
R1114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n945 7.147
R1115 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1022 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1021 7.147
R1116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1019 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1018 7.147
R1117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1016 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1015 7.147
R1118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1013 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1012 7.147
R1119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1008 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1007 7.147
R1120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1005 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1004 7.147
R1121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1002 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1001 7.147
R1122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n997 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n996 7.147
R1123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n994 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n993 7.147
R1124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n991 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n990 7.147
R1125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n987 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n986 7.147
R1126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n984 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n983 7.147
R1127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n981 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n980 7.147
R1128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n978 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n977 7.147
R1129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n975 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n974 7.147
R1130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n970 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n969 7.147
R1131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n967 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n966 7.147
R1132 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n963 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n962 7.147
R1133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n960 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n959 7.147
R1134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n957 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n956 7.147
R1135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n953 7.147
R1136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n949 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n948 7.147
R1137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1028 7.147
R1138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1104 7.147
R1139 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1101 7.147
R1140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1099 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1098 7.147
R1141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1096 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1095 7.147
R1142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1091 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1090 7.147
R1143 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1088 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1087 7.147
R1144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1085 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1084 7.147
R1145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1080 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1079 7.147
R1146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1077 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1076 7.147
R1147 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1074 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1073 7.147
R1148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1070 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1069 7.147
R1149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1067 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1066 7.147
R1150 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1064 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1063 7.147
R1151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1061 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1060 7.147
R1152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1058 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1057 7.147
R1153 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1053 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1052 7.147
R1154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1050 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1049 7.147
R1155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1046 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1045 7.147
R1156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1043 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1042 7.147
R1157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1040 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1039 7.147
R1158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1037 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1036 7.147
R1159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1032 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1031 7.147
R1160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1111 7.147
R1161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1187 7.147
R1162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1184 7.147
R1163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1181 7.147
R1164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1178 7.147
R1165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1173 7.147
R1166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1170 7.147
R1167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1167 7.147
R1168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1162 7.147
R1169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1159 7.147
R1170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1156 7.147
R1171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1153 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1152 7.147
R1172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1150 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1149 7.147
R1173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1147 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1146 7.147
R1174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1143 7.147
R1175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1140 7.147
R1176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1135 7.147
R1177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1132 7.147
R1178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1128 7.147
R1179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1125 7.147
R1180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1122 7.147
R1181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1119 7.147
R1182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1115 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1114 7.147
R1183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1194 7.147
R1184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1271 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1270 7.147
R1185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1267 7.147
R1186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1265 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1264 7.147
R1187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1261 7.147
R1188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1256 7.147
R1189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1254 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1253 7.147
R1190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1250 7.147
R1191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1245 7.147
R1192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1243 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1242 7.147
R1193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1239 7.147
R1194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1236 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1235 7.147
R1195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1232 7.147
R1196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1229 7.147
R1197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1226 7.147
R1198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1223 7.147
R1199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1218 7.147
R1200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1215 7.147
R1201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1211 7.147
R1202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1208 7.147
R1203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1205 7.147
R1204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1202 7.147
R1205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1197 7.147
R1206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1277 7.147
R1207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1354 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1353 7.147
R1208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1351 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1350 7.147
R1209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1348 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1347 7.147
R1210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1344 7.147
R1211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1340 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1339 7.147
R1212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1336 7.147
R1213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1333 7.147
R1214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1329 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1328 7.147
R1215 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1325 7.147
R1216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1322 7.147
R1217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1318 7.147
R1218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1316 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1315 7.147
R1219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1313 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1312 7.147
R1220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1310 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1309 7.147
R1221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1306 7.147
R1222 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1302 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1301 7.147
R1223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1298 7.147
R1224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1295 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1294 7.147
R1225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1291 7.147
R1226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1289 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1288 7.147
R1227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1285 7.147
R1228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1280 7.147
R1229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1360 7.147
R1230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1437 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1436 7.147
R1231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1434 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1433 7.147
R1232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1430 7.147
R1233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1427 7.147
R1234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1423 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1422 7.147
R1235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1419 7.147
R1236 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1416 7.147
R1237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1411 7.147
R1238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1408 7.147
R1239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1405 7.147
R1240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1401 7.147
R1241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1399 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1398 7.147
R1242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1395 7.147
R1243 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1392 7.147
R1244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1389 7.147
R1245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1385 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1384 7.147
R1246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1381 7.147
R1247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1377 7.147
R1248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1375 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1374 7.147
R1249 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1372 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1371 7.147
R1250 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1368 7.147
R1251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1364 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1363 7.147
R1252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1443 7.147
R1253 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1645 7.147
R1254 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1647 7.147
R1255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1649 7.147
R1256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n15 7.147
R1257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n14 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n13 7.147
R1258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n12 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n11 7.147
R1259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n8 7.147
R1260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n7 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n6 7.147
R1261 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n5 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n4 7.147
R1262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n2 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1 7.147
R1263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1485 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1484 7.147
R1264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1481 7.147
R1265 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1478 7.147
R1266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1476 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1475 7.147
R1267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1472 7.147
R1268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1468 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1467 7.147
R1269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1464 7.147
R1270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1461 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1460 7.147
R1271 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1458 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1457 7.147
R1272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1454 7.147
R1273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1451 7.147
R1274 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1447 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1446 7.147
R1275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1605 7.089
R1276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1522 7.089
R1277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n62 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n60 7.089
R1278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n143 7.089
R1279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n226 7.089
R1280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n309 7.089
R1281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n392 7.089
R1282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n475 7.089
R1283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n560 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n558 7.089
R1284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n641 7.089
R1285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n724 7.089
R1286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n807 7.089
R1287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n890 7.089
R1288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n975 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n973 7.089
R1289 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1058 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1056 7.089
R1290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1139 7.089
R1291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1222 7.089
R1292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1305 7.089
R1293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1388 7.089
R1294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1471 7.089
R1295 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1639 6.64
R1296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1644 5.321
R1297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1612 4.945
R1298 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1529 4.945
R1299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n54 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n52 4.945
R1300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n135 4.945
R1301 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n218 4.945
R1302 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n301 4.945
R1303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n384 4.945
R1304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n467 4.945
R1305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n550 4.945
R1306 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n633 4.945
R1307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n716 4.945
R1308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n799 4.945
R1309 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n882 4.945
R1310 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n967 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n965 4.945
R1311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1050 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1048 4.945
R1312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1131 4.945
R1313 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1214 4.945
R1314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1297 4.945
R1315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1380 4.945
R1316 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1463 4.945
R1317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1642 3.497
R1318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1551 3.497
R1319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n33 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n29 3.497
R1320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n112 3.497
R1321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n195 3.497
R1322 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n278 3.497
R1323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n361 3.497
R1324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n444 3.497
R1325 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n527 3.497
R1326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n610 3.497
R1327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n693 3.497
R1328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n776 3.497
R1329 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n859 3.497
R1330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n942 3.497
R1331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1025 3.497
R1332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1108 3.497
R1333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1191 3.497
R1334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1274 3.497
R1335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1357 3.497
R1336 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1440 3.497
R1337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1588 3.132
R1338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1505 3.132
R1339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n78 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n76 3.132
R1340 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n159 3.132
R1341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n242 3.132
R1342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n325 3.132
R1343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n408 3.132
R1344 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n491 3.132
R1345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n574 3.132
R1346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n659 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n657 3.132
R1347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n740 3.132
R1348 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n823 3.132
R1349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n908 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n906 3.132
R1350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n991 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n989 3.132
R1351 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1074 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1072 3.132
R1352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1155 3.132
R1353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1238 3.132
R1354 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1321 3.132
R1355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1404 3.132
R1356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n2 3.132
R1357 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1642 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1640 2.846
R1358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1553 2.846
R1359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n33 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n31 2.846
R1360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n114 2.846
R1361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n197 2.846
R1362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n280 2.846
R1363 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n363 2.846
R1364 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n446 2.846
R1365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n529 2.846
R1366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n612 2.846
R1367 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n695 2.846
R1368 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n778 2.846
R1369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n861 2.846
R1370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n944 2.846
R1371 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1027 2.846
R1372 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1110 2.846
R1373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1193 2.846
R1374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1276 2.846
R1375 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1359 2.846
R1376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1442 2.846
R1377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1637 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1635 2.143
R1378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1543 2.143
R1379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n41 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n39 2.143
R1380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n122 2.143
R1381 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n205 2.143
R1382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n288 2.143
R1383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n371 2.143
R1384 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n454 2.143
R1385 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n537 2.143
R1386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n620 2.143
R1387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n703 2.143
R1388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n786 2.143
R1389 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n869 2.143
R1390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n952 2.143
R1391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1037 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1035 2.143
R1392 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1118 2.143
R1393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1201 2.143
R1394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1284 2.143
R1395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1367 2.143
R1396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1450 2.143
R1397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n20 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n19 1.618
R1398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1652 1.539
R1399 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1567 1.483
R1400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n98 1.483
R1401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n181 1.483
R1402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n264 1.483
R1403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n347 1.483
R1404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n430 1.483
R1405 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n513 1.483
R1406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n598 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n596 1.483
R1407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n679 1.483
R1408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n762 1.483
R1409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n845 1.483
R1410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n928 1.483
R1411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1013 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1011 1.483
R1412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1096 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1094 1.483
R1413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1177 1.483
R1414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1260 1.483
R1415 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1343 1.483
R1416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1426 1.483
R1417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1651 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1630 1.483
R1418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1654 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1653 1.428
R1419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1578 0.329
R1420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1495 0.329
R1421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n89 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n87 0.329
R1422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n170 0.329
R1423 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n253 0.329
R1424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n336 0.329
R1425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n419 0.329
R1426 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n502 0.329
R1427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n585 0.329
R1428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n668 0.329
R1429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n751 0.329
R1430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n834 0.329
R1431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n919 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n917 0.329
R1432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1002 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1000 0.329
R1433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1085 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1083 0.329
R1434 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1166 0.329
R1435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1249 0.329
R1436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1332 0.329
R1437 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1415 0.329
R1438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n10 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n9 0.329
R1439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n24 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n21 0.119
R1440 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n27 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n24 0.119
R1441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n34 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n27 0.119
R1442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n34 0.119
R1443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n37 0.119
R1444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n42 0.119
R1445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n48 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n45 0.119
R1446 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n51 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n48 0.119
R1447 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n55 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n51 0.119
R1448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n58 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n55 0.119
R1449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n63 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n58 0.119
R1450 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n66 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n63 0.119
R1451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n69 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n66 0.119
R1452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n72 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n69 0.119
R1453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n75 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n72 0.119
R1454 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n79 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n75 0.119
R1455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n82 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n79 0.119
R1456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n85 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n82 0.119
R1457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n90 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n85 0.119
R1458 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n90 0.119
R1459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n93 0.119
R1460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n96 0.119
R1461 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n101 0.119
R1462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n104 0.119
R1463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n107 0.119
R1464 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n110 0.119
R1465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n117 0.119
R1466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n120 0.119
R1467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n125 0.119
R1468 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n128 0.119
R1469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n131 0.119
R1470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n134 0.119
R1471 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n138 0.119
R1472 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n141 0.119
R1473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n146 0.119
R1474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n149 0.119
R1475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n152 0.119
R1476 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n155 0.119
R1477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n158 0.119
R1478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n162 0.119
R1479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n165 0.119
R1480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n168 0.119
R1481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n173 0.119
R1482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n176 0.119
R1483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n179 0.119
R1484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n184 0.119
R1485 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n187 0.119
R1486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n190 0.119
R1487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n193 0.119
R1488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n200 0.119
R1489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n203 0.119
R1490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n208 0.119
R1491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n211 0.119
R1492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n214 0.119
R1493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n217 0.119
R1494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n221 0.119
R1495 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n224 0.119
R1496 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n229 0.119
R1497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n232 0.119
R1498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n235 0.119
R1499 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n238 0.119
R1500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n241 0.119
R1501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n245 0.119
R1502 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n248 0.119
R1503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n251 0.119
R1504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n256 0.119
R1505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n259 0.119
R1506 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n262 0.119
R1507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n267 0.119
R1508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n270 0.119
R1509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n273 0.119
R1510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n276 0.119
R1511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n283 0.119
R1512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n286 0.119
R1513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n291 0.119
R1514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n294 0.119
R1515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n297 0.119
R1516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n300 0.119
R1517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n304 0.119
R1518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n307 0.119
R1519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n312 0.119
R1520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n315 0.119
R1521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n318 0.119
R1522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n321 0.119
R1523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n324 0.119
R1524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n328 0.119
R1525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n331 0.119
R1526 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n334 0.119
R1527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n339 0.119
R1528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n342 0.119
R1529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n345 0.119
R1530 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n350 0.119
R1531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n353 0.119
R1532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n356 0.119
R1533 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n359 0.119
R1534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n366 0.119
R1535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n369 0.119
R1536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n374 0.119
R1537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n377 0.119
R1538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n380 0.119
R1539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n383 0.119
R1540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n387 0.119
R1541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n390 0.119
R1542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n395 0.119
R1543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n398 0.119
R1544 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n401 0.119
R1545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n404 0.119
R1546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n407 0.119
R1547 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n411 0.119
R1548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n414 0.119
R1549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n417 0.119
R1550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n422 0.119
R1551 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n425 0.119
R1552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n428 0.119
R1553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n433 0.119
R1554 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n436 0.119
R1555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n439 0.119
R1556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n442 0.119
R1557 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n449 0.119
R1558 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n452 0.119
R1559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n457 0.119
R1560 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n460 0.119
R1561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n463 0.119
R1562 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n466 0.119
R1563 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n470 0.119
R1564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n473 0.119
R1565 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n478 0.119
R1566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n481 0.119
R1567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n484 0.119
R1568 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n487 0.119
R1569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n490 0.119
R1570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n494 0.119
R1571 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n497 0.119
R1572 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n500 0.119
R1573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n505 0.119
R1574 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n508 0.119
R1575 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n511 0.119
R1576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n516 0.119
R1577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n519 0.119
R1578 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n522 0.119
R1579 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n525 0.119
R1580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n532 0.119
R1581 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n535 0.119
R1582 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n540 0.119
R1583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n543 0.119
R1584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n546 0.119
R1585 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n549 0.119
R1586 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n553 0.119
R1587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n556 0.119
R1588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n561 0.119
R1589 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n564 0.119
R1590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n567 0.119
R1591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n570 0.119
R1592 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n573 0.119
R1593 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n577 0.119
R1594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n580 0.119
R1595 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n583 0.119
R1596 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n588 0.119
R1597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n591 0.119
R1598 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n594 0.119
R1599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n599 0.119
R1600 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n602 0.119
R1601 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n605 0.119
R1602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n608 0.119
R1603 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n615 0.119
R1604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n618 0.119
R1605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n623 0.119
R1606 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n626 0.119
R1607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n629 0.119
R1608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n636 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n632 0.119
R1609 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n636 0.119
R1610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n639 0.119
R1611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n644 0.119
R1612 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n647 0.119
R1613 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n650 0.119
R1614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n653 0.119
R1615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n660 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n656 0.119
R1616 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n660 0.119
R1617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n663 0.119
R1618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n666 0.119
R1619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n671 0.119
R1620 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n674 0.119
R1621 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n677 0.119
R1622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n682 0.119
R1623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n685 0.119
R1624 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n688 0.119
R1625 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n691 0.119
R1626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n698 0.119
R1627 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n701 0.119
R1628 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n706 0.119
R1629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n709 0.119
R1630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n712 0.119
R1631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n715 0.119
R1632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n719 0.119
R1633 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n722 0.119
R1634 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n727 0.119
R1635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n730 0.119
R1636 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n733 0.119
R1637 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n736 0.119
R1638 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n739 0.119
R1639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n743 0.119
R1640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n746 0.119
R1641 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n749 0.119
R1642 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n754 0.119
R1643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n757 0.119
R1644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n760 0.119
R1645 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n765 0.119
R1646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n768 0.119
R1647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n771 0.119
R1648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n774 0.119
R1649 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n781 0.119
R1650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n784 0.119
R1651 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n789 0.119
R1652 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n792 0.119
R1653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n795 0.119
R1654 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n798 0.119
R1655 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n802 0.119
R1656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n805 0.119
R1657 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n810 0.119
R1658 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n813 0.119
R1659 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n816 0.119
R1660 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n819 0.119
R1661 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n822 0.119
R1662 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n826 0.119
R1663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n829 0.119
R1664 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n832 0.119
R1665 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n837 0.119
R1666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n840 0.119
R1667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n843 0.119
R1668 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n848 0.119
R1669 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n851 0.119
R1670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n854 0.119
R1671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n857 0.119
R1672 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n864 0.119
R1673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n867 0.119
R1674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n872 0.119
R1675 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n875 0.119
R1676 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n878 0.119
R1677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n881 0.119
R1678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n885 0.119
R1679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n888 0.119
R1680 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n896 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n893 0.119
R1681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n896 0.119
R1682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n902 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n899 0.119
R1683 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n905 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n902 0.119
R1684 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n909 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n905 0.119
R1685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n912 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n909 0.119
R1686 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n915 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n912 0.119
R1687 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n920 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n915 0.119
R1688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n923 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n920 0.119
R1689 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n926 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n923 0.119
R1690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n926 0.119
R1691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n934 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n931 0.119
R1692 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n937 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n934 0.119
R1693 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n940 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n937 0.119
R1694 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n947 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n940 0.119
R1695 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n950 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n947 0.119
R1696 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n950 0.119
R1697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n958 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n955 0.119
R1698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n961 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n958 0.119
R1699 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n964 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n961 0.119
R1700 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n964 0.119
R1701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n968 0.119
R1702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n976 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n971 0.119
R1703 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n979 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n976 0.119
R1704 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n982 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n979 0.119
R1705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n985 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n982 0.119
R1706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n988 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n985 0.119
R1707 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n992 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n988 0.119
R1708 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n992 0.119
R1709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n998 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n995 0.119
R1710 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1003 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n998 0.119
R1711 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1006 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1003 0.119
R1712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1009 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1006 0.119
R1713 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1014 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1009 0.119
R1714 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1017 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1014 0.119
R1715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1020 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1017 0.119
R1716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1023 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1020 0.119
R1717 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1030 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1023 0.119
R1718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1033 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1030 0.119
R1719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1038 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1033 0.119
R1720 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1041 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1038 0.119
R1721 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1044 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1041 0.119
R1722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1047 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1044 0.119
R1723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1051 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1047 0.119
R1724 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1054 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1051 0.119
R1725 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1059 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1054 0.119
R1726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1059 0.119
R1727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1065 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1062 0.119
R1728 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1068 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1065 0.119
R1729 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1071 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1068 0.119
R1730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1075 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1071 0.119
R1731 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1078 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1075 0.119
R1732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1081 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1078 0.119
R1733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1086 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1081 0.119
R1734 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1089 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1086 0.119
R1735 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1092 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1089 0.119
R1736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1097 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1092 0.119
R1737 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1097 0.119
R1738 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1100 0.119
R1739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1103 0.119
R1740 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1106 0.119
R1741 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1113 0.119
R1742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1116 0.119
R1743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1121 0.119
R1744 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1124 0.119
R1745 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1127 0.119
R1746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1130 0.119
R1747 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1134 0.119
R1748 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1137 0.119
R1749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1142 0.119
R1750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1145 0.119
R1751 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1148 0.119
R1752 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1151 0.119
R1753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1154 0.119
R1754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1158 0.119
R1755 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1161 0.119
R1756 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1164 0.119
R1757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1169 0.119
R1758 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1172 0.119
R1759 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1175 0.119
R1760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1180 0.119
R1761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1183 0.119
R1762 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1186 0.119
R1763 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1189 0.119
R1764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1196 0.119
R1765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1199 0.119
R1766 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1204 0.119
R1767 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1207 0.119
R1768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1210 0.119
R1769 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1213 0.119
R1770 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1217 0.119
R1771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1220 0.119
R1772 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1225 0.119
R1773 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1228 0.119
R1774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1231 0.119
R1775 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1234 0.119
R1776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1237 0.119
R1777 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1241 0.119
R1778 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1244 0.119
R1779 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1247 0.119
R1780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1252 0.119
R1781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1255 0.119
R1782 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1258 0.119
R1783 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1263 0.119
R1784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1266 0.119
R1785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1269 0.119
R1786 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1272 0.119
R1787 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1279 0.119
R1788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1282 0.119
R1789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1287 0.119
R1790 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1290 0.119
R1791 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1293 0.119
R1792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1296 0.119
R1793 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1300 0.119
R1794 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1303 0.119
R1795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1308 0.119
R1796 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1311 0.119
R1797 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1314 0.119
R1798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1317 0.119
R1799 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1320 0.119
R1800 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1324 0.119
R1801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1327 0.119
R1802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1330 0.119
R1803 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1335 0.119
R1804 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1338 0.119
R1805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1341 0.119
R1806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1346 0.119
R1807 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1349 0.119
R1808 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1352 0.119
R1809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1355 0.119
R1810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1362 0.119
R1811 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1365 0.119
R1812 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1370 0.119
R1813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1373 0.119
R1814 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1376 0.119
R1815 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1379 0.119
R1816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1383 0.119
R1817 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1386 0.119
R1818 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1391 0.119
R1819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1394 0.119
R1820 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1397 0.119
R1821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1400 0.119
R1822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1403 0.119
R1823 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1407 0.119
R1824 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1410 0.119
R1825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1413 0.119
R1826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1418 0.119
R1827 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1421 0.119
R1828 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1424 0.119
R1829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1429 0.119
R1830 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1432 0.119
R1831 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1435 0.119
R1832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1438 0.119
R1833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1445 0.119
R1834 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1448 0.119
R1835 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1453 0.119
R1836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1456 0.119
R1837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1459 0.119
R1838 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1462 0.119
R1839 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1466 0.119
R1840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1469 0.119
R1841 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1474 0.119
R1842 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1477 0.119
R1843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1480 0.119
R1844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1483 0.119
R1845 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1486 0.119
R1846 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1487 0.119
R1847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1488 0.119
R1848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1489 0.119
R1849 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1490 0.119
R1850 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1491 0.119
R1851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1492 0.119
R1852 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1628 0.119
R1853 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1628 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1627 0.119
R1854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1627 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1626 0.119
R1855 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1625 0.119
R1856 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1625 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1624 0.119
R1857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1624 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1623 0.119
R1858 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1622 0.119
R1859 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1621 0.119
R1860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1621 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1618 0.119
R1861 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1615 0.119
R1862 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1611 0.119
R1863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1608 0.119
R1864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1603 0.119
R1865 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1603 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1600 0.119
R1866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1600 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1597 0.119
R1867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1594 0.119
R1868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1591 0.119
R1869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1587 0.119
R1870 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1584 0.119
R1871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1581 0.119
R1872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1581 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1576 0.119
R1873 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1573 0.119
R1874 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1570 0.119
R1875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1565 0.119
R1876 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1565 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1562 0.119
R1877 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1562 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1559 0.119
R1878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1556 0.119
R1879 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1549 0.119
R1880 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1546 0.119
R1881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1541 0.119
R1882 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1538 0.119
R1883 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1535 0.119
R1884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1532 0.119
R1885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1528 0.119
R1886 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1525 0.119
R1887 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1520 0.119
R1888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1517 0.119
R1889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1514 0.119
R1890 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1511 0.119
R1891 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1508 0.119
R1892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1504 0.119
R1893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1501 0.119
R1894 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1498 0.119
C0 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6541_47# 0.08fF
C1 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1283_21# 0.22fF
C2 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11231_413# 0.17fF
C3 a_1108_47# a_1283_21# 0.62fF
C4 a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C5 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8491_47# 0.99fF
C6 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32283_47# 0.36fF
C7 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C8 a_8491_47# a_8912_47# 0.23fF
C9 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# 0.24fF
C10 a_16955_47# a_17376_47# 0.23fF
C11 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# 0.24fF
C12 a_39371_21# a_39935_47# 0.30fF
C13 a_19492_47# a_19071_47# 0.23fF
C14 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.24fF
C15 a_21187_47# a_21608_47# 0.23fF
C16 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# 0.24fF
C17 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2921_47# 0.01fF
C18 a_40965_289# a_40855_413# 0.23fF
C19 a_29817_47# a_30072_47# 0.22fF
C20 a_9572_47# a_9681_47# 0.04fF
C21 a_23819_47# a_24384_47# 0.01fF
C22 a_37080_47# a_36623_413# 0.01fF
C23 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.12fF
C24 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38849_289# 0.46fF
C25 a_7109_289# a_7456_47# 0.13fF
C26 a_6891_47# a_7631_21# 0.02fF
C27 a_29651_47# a_30907_21# 0.12fF
C28 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30167_47# 0.09fF
C29 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9926_47# 0.01fF
C30 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23927_413# 0.01fF
C31 a_36733_289# a_37080_47# 0.13fF
C32 a_31471_47# a_31933_47# 0.01fF
C33 a_13979_21# a_14839_47# 0.02fF
C34 a_19805_289# a_19587_47# 0.50fF
C35 a_27239_47# a_26500_47# 0.00fF
C36 a_26031_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.02fF
C37 a_26043_413# a_25935_47# 0.21fF
C38 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_38115_47# 0.02fF
C39 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.11fF
C40 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.27fF
C41 a_35999_47# a_36515_47# 0.42fF
C42 a_543_47# a_1283_21# 0.02fF
C43 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6796_47# 0.53fF
C44 a_38739_413# a_38849_289# 0.23fF
C45 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4425_47# 0.08fF
C46 a_32848_47# a_32957_47# 0.04fF
C47 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23007_47# 0.01fF
C48 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13501_47# 0.01fF
C49 a_8657_47# a_9225_289# 0.41fF
C50 a_25123_47# a_25585_47# 0.01fF
C51 a_13913_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.01fF
C52 a_39371_21# a_39550_47# 0.04fF
C53 a_39196_47# a_39305_47# 0.04fF
C54 a_32501_289# a_33023_21# 0.03fF
C55 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28616_47# 0.02fF
C56 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.68fF
C57 a_4993_289# a_5515_21# 0.03fF
C58 a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.05fF
C59 a_10607_47# a_11863_21# 0.12fF
C60 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11123_47# 0.09fF
C61 a_28051_47# a_28616_47# 0.01fF
C62 a_3399_21# a_3963_47# 0.30fF
C63 a_2659_47# a_2564_47# 0.13fF
C64 a_2877_289# a_2767_413# 0.23fF
C65 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25585_47# 0.08fF
C66 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26043_413# 0.17fF
C67 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.27fF
C68 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12042_47# 0.01fF
C69 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16659_47# 0.09fF
C70 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11688_47# 0.68fF
C71 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20891_47# 0.09fF
C72 a_26153_289# a_26675_21# 0.03fF
C73 a_25585_47# a_26500_47# 0.29fF
C74 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_10607_47# 0.02fF
C75 a_38849_289# a_38631_47# 0.50fF
C76 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# 0.27fF
C77 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[7]/D 1.68fF
C78 a_8491_47# a_9747_21# 0.12fF
C79 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9007_47# 0.09fF
C80 a_16955_47# a_18211_21# 0.12fF
C81 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17471_47# 0.09fF
C82 a_24037_289# a_24559_21# 0.03fF
C83 a_23469_47# a_24384_47# 0.29fF
C84 a_20327_21# a_19071_47# 0.12fF
C85 a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.09fF
C86 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21703_47# 0.09fF
C87 a_21187_47# a_22443_21# 0.12fF
C88 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_27956_47# 0.06fF
C89 a_34399_47# a_35139_21# 0.02fF
C90 a_13804_47# a_14543_47# 0.00fF
C91 a_13239_47# a_13347_413# 0.21fF
C92 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16955_47# 0.02fF
C93 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8195_47# 0.09fF
C94 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_21187_47# 0.02fF
C95 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_15005_47# 0.08fF
C96 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_27701_47# 1.17fF
C97 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28159_413# 0.01fF
C98 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.11fF
C99 a_11688_47# a_11850_413# 0.04fF
C100 a_6541_47# a_6891_47# 0.49fF
C101 a_16095_21# a_15920_47# 0.62fF
C102 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4680_47# 0.53fF
C103 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28269_289# 0.10fF
C104 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30894_413# 0.01fF
C105 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.01fF
C106 a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.01fF
C107 a_39305_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C108 a_32391_413# a_32283_47# 0.21fF
C109 a_32379_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.02fF
C110 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34304_47# 0.53fF
C111 a_10607_47# a_11341_289# 0.16fF
C112 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_10773_47# 0.65fF
C113 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.02fF
C114 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.63fF
C115 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40652_47# 0.53fF
C116 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30732_47# 0.68fF
C117 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13347_413# 0.17fF
C118 a_6375_47# a_7456_47# 0.27fF
C119 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7631_21# 0.22fF
C120 a_11123_47# a_11219_47# 0.07fF
C121 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34049_47# 0.65fF
C122 a_33883_47# a_34617_289# 0.16fF
C123 a_23303_47# a_22443_21# 0.02fF
C124 a_40231_47# a_40965_289# 0.16fF
C125 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40397_47# 0.65fF
C126 a_16955_47# a_17689_289# 0.16fF
C127 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17121_47# 0.65fF
C128 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_29355_47# 0.01fF
C129 a_36515_47# a_36611_47# 0.07fF
C130 a_19805_289# a_19071_47# 0.16fF
C131 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21353_47# 0.65fF
C132 a_21187_47# a_21921_289# 0.16fF
C133 a_2877_289# a_3224_47# 0.13fF
C134 a_2659_47# a_3399_21# 0.02fF
C135 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33023_21# 0.73fF
C136 a_13457_289# a_13144_47# 0.00fF
C137 a_12889_47# a_13347_413# 0.12fF
C138 a_41421_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C139 a_39196_47# a_39935_47# 0.00fF
C140 a_30072_47# a_30275_413# 0.02fF
C141 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19587_47# 0.36fF
C142 a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.09fF
C143 a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.02fF
C144 a_8491_47# a_8657_47# 1.60fF
C145 a_35999_47# a_35703_47# 0.07fF
C146 a_30385_289# a_30072_47# 0.00fF
C147 a_29817_47# a_30275_413# 0.12fF
C148 a_15573_289# a_15920_47# 0.13fF
C149 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35999_47# 0.99fF
C150 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_6375_47# 0.02fF
C151 a_4425_47# a_4775_47# 0.49fF
C152 a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.02fF
C153 a_13239_47# a_13804_47# 0.01fF
C154 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2564_47# 0.53fF
C155 a_23724_47# a_23927_413# 0.02fF
C156 a_20261_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C157 a_29817_47# a_30385_289# 0.41fF
C158 a_29651_47# a_30732_47# 0.27fF
C159 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30907_21# 0.22fF
C160 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6891_47# 0.36fF
C161 a_1217_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C162 a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.71fF
C163 a_32848_47# a_33010_413# 0.04fF
C164 a_15463_413# a_15920_47# 0.01fF
C165 a_1108_47# a_1217_47# 0.04fF
C166 a_23303_47# a_24559_21# 0.12fF
C167 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.01fF
C168 a_36165_47# a_36420_47# 0.22fF
C169 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23819_47# 0.09fF
C170 a_4259_47# a_5340_47# 0.27fF
C171 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5515_21# 0.22fF
C172 a_26197_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C173 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.01fF
C174 a_23469_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C175 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36515_47# 0.09fF
C176 a_35999_47# a_37255_21# 0.12fF
C177 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_23303_47# 0.02fF
C178 a_30907_21# a_31767_47# 0.02fF
C179 a_11863_21# a_12723_47# 0.02fF
C180 a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.63fF
C181 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C182 a_37819_47# a_38281_47# 0.01fF
C183 a_18775_47# a_19237_47# 0.01fF
C184 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13804_47# 0.68fF
C185 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_29355_47# 0.36fF
C186 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11385_47# 0.01fF
C187 a_6375_47# a_7109_289# 0.16fF
C188 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6541_47# 0.65fF
C189 a_38536_47# a_38115_47# 0.23fF
C190 a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.24fF
C191 a_10311_47# a_10773_47# 0.01fF
C192 a_28791_21# a_28616_47# 0.62fF
C193 a_31767_47# a_32283_47# 0.42fF
C194 a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.36fF
C195 a_41009_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C196 a_26153_289# a_26500_47# 0.13fF
C197 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.27fF
C198 a_2309_47# a_2659_47# 0.49fF
C199 a_13457_289# a_13979_21# 0.03fF
C200 a_12889_47# a_13804_47# 0.29fF
C201 a_15451_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.02fF
C202 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_34964_47# 0.02fF
C203 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C204 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28159_413# 0.17fF
C205 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[5]/D 1.68fF
C206 a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.36fF
C207 a_34399_47# a_34964_47# 0.01fF
C208 a_25419_47# a_25935_47# 0.42fF
C209 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23469_47# 0.65fF
C210 a_23303_47# a_24037_289# 0.16fF
C211 a_15005_47# a_15355_47# 0.49fF
C212 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28269_289# 0.46fF
C213 a_9572_47# a_9734_413# 0.04fF
C214 a_2143_47# a_3224_47# 0.27fF
C215 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3399_21# 0.22fF
C216 a_12723_47# a_13144_47# 0.23fF
C217 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# 0.24fF
C218 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12889_47# 0.08fF
C219 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19071_47# 0.99fF
C220 a_11028_47# a_11231_413# 0.02fF
C221 a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.02fF
C222 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25419_47# 0.99fF
C223 a_8657_47# a_8195_47# 0.01fF
C224 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37434_47# 0.01fF
C225 a_15260_47# a_15355_47# 0.13fF
C226 a_16659_47# a_16095_21# 0.30fF
C227 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C228 a_32545_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C229 a_14839_47# a_15920_47# 0.27fF
C230 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16095_21# 0.22fF
C231 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34507_413# 0.01fF
C232 a_4259_47# a_4993_289# 0.16fF
C233 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40855_413# 0.01fF
C234 sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C235 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39371_21# 0.73fF
C236 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31471_47# 0.09fF
C237 a_17376_47# a_17579_413# 0.02fF
C238 a_21608_47# a_21811_413# 0.02fF
C239 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[3]/D 1.68fF
C240 a_32848_47# a_31933_47# 0.29fF
C241 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C242 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34617_289# 0.10fF
C243 a_20152_47# a_20314_413# 0.04fF
C244 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_2143_47# 0.02fF
C245 a_40747_47# a_41487_21# 0.02fF
C246 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40965_289# 0.10fF
C247 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.01fF
C248 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.01fF
C249 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C250 a_37434_47# a_37255_21# 0.04fF
C251 a_37189_47# a_37080_47# 0.04fF
C252 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.08fF
C253 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0.36fF
C254 a_29817_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.08fF
C255 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C256 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17376_47# 0.06fF
C257 a_6079_47# a_6541_47# 0.01fF
C258 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21608_47# 0.06fF
C259 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3578_47# 0.01fF
C260 a_19587_47# a_19683_47# 0.07fF
C261 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_35703_47# 0.01fF
C262 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[17]/D 1.68fF
C263 a_30385_289# a_30275_413# 0.23fF
C264 a_15260_47# a_15005_47# 0.22fF
C265 a_23819_47# a_23724_47# 0.13fF
C266 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.12fF
C267 a_36420_47# a_36623_413# 0.02fF
C268 sky130_fd_sc_hd__dfrbp_1_0[9]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.12fF
C269 a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.37fF
C270 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15573_289# 0.10fF
C271 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30732_47# 0.05fF
C272 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10311_47# 0.09fF
C273 a_39371_21# a_38631_47# 0.02fF
C274 a_22622_47# a_22443_21# 0.04fF
C275 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2309_47# 0.65fF
C276 a_2143_47# a_2877_289# 0.16fF
C277 a_12723_47# a_13979_21# 0.12fF
C278 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13239_47# 0.09fF
C279 a_9572_47# a_9115_413# 0.01fF
C280 a_36733_289# a_36420_47# 0.00fF
C281 a_36165_47# a_36623_413# 0.12fF
C282 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38115_47# 0.99fF
C283 a_5340_47# a_5502_413# 0.04fF
C284 a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.36fF
C285 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.68fF
C286 a_26043_413# a_26500_47# 0.01fF
C287 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_12723_47# 0.02fF
C288 a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C289 sky130_fd_sc_hd__dfrbp_1_0[12]/Q sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.12fF
C290 a_32848_47# a_33587_47# 0.00fF
C291 a_36165_47# a_36733_289# 0.41fF
C292 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37255_21# 0.22fF
C293 a_35999_47# a_37080_47# 0.27fF
C294 sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.08fF
C295 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# 0.27fF
C296 a_28616_47# a_28778_413# 0.04fF
C297 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.01fF
C298 a_651_413# a_761_289# 0.23fF
C299 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9269_47# 0.01fF
C300 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31086_47# 0.01fF
C301 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9926_47# 0.01fF
C302 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.53fF
C303 a_28791_21# a_29355_47# 0.30fF
C304 a_28051_47# a_27956_47# 0.13fF
C305 a_31767_47# a_33023_21# 0.12fF
C306 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32283_47# 0.09fF
C307 a_37255_21# a_38115_47# 0.02fF
C308 sky130_fd_sc_hd__dfrbp_1_0[19]/Q sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.12fF
C309 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[6]/D 1.68fF
C310 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6079_47# 0.09fF
C311 a_20327_21# a_21187_47# 0.02fF
C312 a_639_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.02fF
C313 a_27701_47# a_28051_47# 0.49fF
C314 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35703_47# 0.36fF
C315 a_448_47# a_651_413# 0.02fF
C316 a_23469_47# a_23724_47# 0.22fF
C317 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18211_21# 0.73fF
C318 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22443_21# 0.73fF
C319 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[16]/Q 0.11fF
C320 a_35139_21# a_34964_47# 0.62fF
C321 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.04fF
C322 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4680_47# 0.01fF
C323 a_25419_47# a_26675_21# 0.12fF
C324 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_25935_47# 0.09fF
C325 a_38115_47# a_38631_47# 0.42fF
C326 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_12889_47# 0.65fF
C327 a_12723_47# a_13457_289# 0.16fF
C328 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34399_47# 0.36fF
C329 a_28970_47# a_28791_21# 0.04fF
C330 a_28725_47# a_28616_47# 0.04fF
C331 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.11fF
C332 a_11341_289# a_11231_413# 0.23fF
C333 a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.71fF
C334 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.11fF
C335 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10773_47# 0.08fF
C336 a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.71fF
C337 sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.12fF
C338 a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.02fF
C339 a_30841_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C340 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9007_47# 0.36fF
C341 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[12]/D 1.68fF
C342 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39358_413# 0.01fF
C343 a_9007_47# a_8912_47# 0.13fF
C344 a_9747_21# a_10311_47# 0.30fF
C345 a_9225_289# a_9115_413# 0.23fF
C346 a_17689_289# a_17579_413# 0.23fF
C347 a_11863_21# a_12042_47# 0.04fF
C348 a_11688_47# a_11797_47# 0.04fF
C349 a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.27fF
C350 sky130_fd_sc_hd__dfrbp_1_0[15]/Q sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.12fF
C351 a_21921_289# a_21811_413# 0.23fF
C352 a_5340_47# a_4883_413# 0.01fF
C353 a_11863_21# a_11688_47# 0.62fF
C354 a_20152_47# a_20891_47# 0.00fF
C355 a_19587_47# a_19695_413# 0.21fF
C356 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39196_47# 0.68fF
C357 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30072_47# 0.06fF
C358 a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.71fF
C359 a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.71fF
C360 a_32848_47# a_32501_289# 0.13fF
C361 a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.86fF
C362 a_639_47# a_543_47# 0.07fF
C363 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_761_289# 0.10fF
C364 a_1108_47# a_761_289# 0.13fF
C365 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24559_21# 0.73fF
C366 a_40747_47# a_41312_47# 0.01fF
C367 a_18211_21# a_18036_47# 0.62fF
C368 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_29817_47# 1.17fF
C369 a_22443_21# a_22268_47# 0.62fF
C370 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17689_289# 0.46fF
C371 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21921_289# 0.46fF
C372 a_9747_21# a_9926_47# 0.04fF
C373 a_8657_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C374 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.08fF
C375 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[10]/Q 0.11fF
C376 a_1847_47# a_2143_47# 0.07fF
C377 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23915_47# 0.02fF
C378 a_39196_47# a_38739_413# 0.01fF
C379 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4775_47# 0.36fF
C380 a_14543_47# a_15005_47# 0.01fF
C381 a_26031_47# a_25935_47# 0.07fF
C382 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.53fF
C383 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C384 a_7456_47# a_8195_47# 0.00fF
C385 a_6891_47# a_6999_413# 0.21fF
C386 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.12fF
C387 a_36165_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C388 a_23819_47# a_23927_413# 0.21fF
C389 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# 0.63fF
C390 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_40231_47# 0.02fF
C391 a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.63fF
C392 a_29651_47# a_30072_47# 0.23fF
C393 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# 0.24fF
C394 a_11341_289# a_11688_47# 0.13fF
C395 a_39196_47# a_38631_47# 0.01fF
C396 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.11fF
C397 a_19805_289# a_19492_47# 0.00fF
C398 a_36733_289# a_36623_413# 0.23fF
C399 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[18]/D 1.68fF
C400 a_761_289# a_543_47# 0.50fF
C401 a_29651_47# a_29817_47# 1.60fF
C402 a_193_47# a_1283_21# 0.10fF
C403 a_3963_47# a_4259_47# 0.07fF
C404 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40747_47# 0.36fF
C405 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24037_289# 0.46fF
C406 a_9225_289# a_9572_47# 0.13fF
C407 a_9007_47# a_9747_21# 0.02fF
C408 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_27535_47# 0.02fF
C409 a_17689_289# a_18036_47# 0.13fF
C410 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37080_47# 0.05fF
C411 a_31471_47# a_31767_47# 0.07fF
C412 a_21921_289# a_22268_47# 0.13fF
C413 a_4775_47# a_4680_47# 0.13fF
C414 a_5515_21# a_6079_47# 0.30fF
C415 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11028_47# 0.53fF
C416 a_2143_47# a_1283_21# 0.02fF
C417 a_4993_289# a_4883_413# 0.23fF
C418 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22268_47# 0.02fF
C419 a_19587_47# a_20152_47# 0.01fF
C420 a_25840_47# a_25585_47# 0.22fF
C421 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33010_413# 0.01fF
C422 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C423 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28147_47# 0.02fF
C424 a_1847_47# a_1283_21# 0.30fF
C425 a_28051_47# a_28159_413# 0.21fF
C426 a_448_47# a_543_47# 0.13fF
C427 a_28616_47# a_29355_47# 0.00fF
C428 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[4]/D 1.68fF
C429 a_25123_47# a_25419_47# 0.07fF
C430 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_8912_47# 0.53fF
C431 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33023_21# 0.22fF
C432 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15355_47# 0.36fF
C433 a_31933_47# a_32501_289# 0.41fF
C434 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17376_47# 0.53fF
C435 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32848_47# 0.68fF
C436 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.53fF
C437 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21608_47# 0.53fF
C438 a_34964_47# a_35126_413# 0.04fF
C439 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.12fF
C440 a_13144_47# a_13347_413# 0.02fF
C441 a_28269_289# a_28051_47# 0.50fF
C442 a_27701_47# a_28791_21# 0.10fF
C443 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33202_47# 0.01fF
C444 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# 0.63fF
C445 a_23469_47# a_23927_413# 0.12fF
C446 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5694_47# 0.01fF
C447 a_32379_47# a_32283_47# 0.07fF
C448 a_27_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.71fF
C449 a_25585_47# a_26153_289# 0.41fF
C450 a_25419_47# a_26500_47# 0.27fF
C451 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26675_21# 0.22fF
C452 a_34399_47# a_34304_47# 0.13fF
C453 a_35139_21# a_35703_47# 0.30fF
C454 a_1108_47# a_27_47# 0.27fF
C455 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38631_47# 0.09fF
C456 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35139_21# 0.73fF
C457 a_24559_21# a_24384_47# 0.62fF
C458 a_6891_47# a_7456_47# 0.01fF
C459 a_6541_47# a_6796_47# 0.22fF
C460 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16955_47# 0.99fF
C461 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21187_47# 0.99fF
C462 a_34049_47# a_34399_47# 0.49fF
C463 a_23469_47# a_23007_47# 0.01fF
C464 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.11fF
C465 a_4425_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.17fF
C466 a_10773_47# a_11123_47# 0.49fF
C467 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_27535_47# 0.99fF
C468 a_19805_289# a_20327_21# 0.03fF
C469 a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C470 a_35318_47# a_35139_21# 0.04fF
C471 a_35073_47# a_34964_47# 0.04fF
C472 a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.02fF
C473 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6999_413# 0.01fF
C474 a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.02fF
C475 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.12fF
C476 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39935_47# 0.09fF
C477 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15005_47# 1.17fF
C478 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30275_413# 0.17fF
C479 a_8657_47# a_9007_47# 0.49fF
C480 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11797_47# 0.01fF
C481 a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.01fF
C482 a_17121_47# a_17471_47# 0.49fF
C483 a_19587_47# a_19237_47# 0.49fF
C484 a_21353_47# a_21703_47# 0.49fF
C485 a_32188_47# a_31933_47# 0.22fF
C486 a_10607_47# a_11688_47# 0.27fF
C487 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11863_21# 0.22fF
C488 a_3224_47# a_3963_47# 0.00fF
C489 a_2659_47# a_2767_413# 0.21fF
C490 a_4993_289# a_5340_47# 0.13fF
C491 a_4775_47# a_5515_21# 0.02fF
C492 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# 0.27fF
C493 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30385_289# 0.46fF
C494 a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.02fF
C495 a_41487_21# a_41312_47# 0.62fF
C496 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13966_413# 0.01fF
C497 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.27fF
C498 a_18390_47# a_18211_21# 0.04fF
C499 a_18145_47# a_18036_47# 0.04fF
C500 a_30167_47# a_30907_21# 0.02fF
C501 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12427_47# 0.09fF
C502 a_20327_21# a_20506_47# 0.04fF
C503 a_27_47# a_543_47# 0.42fF
C504 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.01fF
C505 a_20152_47# a_20261_47# 0.04fF
C506 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15260_47# 0.06fF
C507 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19492_47# 0.06fF
C508 a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.71fF
C509 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23303_47# 0.99fF
C510 a_8491_47# a_9572_47# 0.27fF
C511 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9747_21# 0.22fF
C512 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24081_47# 0.01fF
C513 a_16955_47# a_18036_47# 0.27fF
C514 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18211_21# 0.22fF
C515 a_24037_289# a_24384_47# 0.13fF
C516 a_20152_47# a_19071_47# 0.27fF
C517 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.22fF
C518 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_22443_21# 0.22fF
C519 a_21187_47# a_22268_47# 0.27fF
C520 a_4425_47# a_4680_47# 0.22fF
C521 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31933_47# 1.17fF
C522 a_12427_47# a_12889_47# 0.01fF
C523 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6796_47# 0.06fF
C524 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# 0.63fF
C525 a_7810_47# a_7631_21# 0.04fF
C526 a_7565_47# a_7456_47# 0.04fF
C527 a_7109_289# a_6891_47# 0.50fF
C528 a_6541_47# a_7631_21# 0.10fF
C529 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30072_47# 0.53fF
C530 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4883_413# 0.01fF
C531 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_39550_47# 0.01fF
C532 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_13144_47# 0.01fF
C533 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_29817_47# 0.65fF
C534 a_29651_47# a_30385_289# 0.16fF
C535 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41487_21# 0.67fF
C536 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11341_289# 0.10fF
C537 a_16082_413# a_15920_47# 0.04fF
C538 a_32848_47# a_32391_413# 0.01fF
C539 a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C540 a_35999_47# a_36420_47# 0.23fF
C541 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# 0.24fF
C542 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7456_47# 0.05fF
C543 a_25840_47# a_26153_289# 0.00fF
C544 a_26043_413# a_25585_47# 0.12fF
C545 a_27239_47# a_27701_47# 0.01fF
C546 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17689_289# 0.10fF
C547 a_35999_47# a_36165_47# 1.60fF
C548 a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.10fF
C549 a_5515_21# a_5694_47# 0.04fF
C550 a_5340_47# a_5449_47# 0.04fF
C551 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21921_289# 0.10fF
C552 a_13457_289# a_13347_413# 0.23fF
C553 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33883_47# 0.02fF
C554 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28313_47# 0.01fF
C555 a_2659_47# a_3224_47# 0.01fF
C556 a_2309_47# a_2564_47# 0.22fF
C557 a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C558 sky130_fd_sc_hd__dfrbp_1_0[10]/Q sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.12fF
C559 a_15451_47# a_15355_47# 0.07fF
C560 a_37819_47# a_38115_47# 0.07fF
C561 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33587_47# 0.09fF
C562 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.06fF
C563 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11123_47# 0.36fF
C564 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20327_21# 0.73fF
C565 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# 0.63fF
C566 a_26609_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C567 a_19071_47# a_19237_47# 1.60fF
C568 a_28269_289# a_28791_21# 0.03fF
C569 a_27701_47# a_28616_47# 0.29fF
C570 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_8657_47# 0.65fF
C571 a_8491_47# a_9225_289# 0.16fF
C572 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35126_413# 0.01fF
C573 a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.36fF
C574 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C575 a_24738_47# a_24559_21# 0.04fF
C576 a_23469_47# a_23819_47# 0.49fF
C577 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34495_47# 0.02fF
C578 a_4425_47# a_5515_21# 0.10fF
C579 a_34399_47# a_34507_413# 0.21fF
C580 a_34964_47# a_35703_47# 0.00fF
C581 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.36fF
C582 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26500_47# 0.05fF
C583 a_13979_21# a_13804_47# 0.62fF
C584 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2767_413# 0.01fF
C585 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40843_47# 0.02fF
C586 a_38281_47# a_38849_289# 0.41fF
C587 a_27535_47# a_26675_21# 0.02fF
C588 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34964_47# 0.68fF
C589 a_24559_21# a_25123_47# 0.30fF
C590 a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C591 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7631_21# 0.73fF
C592 a_34617_289# a_34399_47# 0.50fF
C593 a_34049_47# a_35139_21# 0.10fF
C594 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C595 a_22377_47# a_22268_47# 0.04fF
C596 a_23303_47# a_24384_47# 0.27fF
C597 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24559_21# 0.22fF
C598 a_15355_47# a_16095_21# 0.02fF
C599 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5340_47# 0.05fF
C600 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[13]/D 1.68fF
C601 a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.36fF
C602 a_3399_21# a_3578_47# 0.04fF
C603 a_3224_47# a_3333_47# 0.04fF
C604 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9681_47# 0.01fF
C605 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# 0.63fF
C606 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38536_47# 0.06fF
C607 a_41312_47# a_41474_413# 0.04fF
C608 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14543_47# 0.09fF
C609 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.12fF
C610 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7109_289# 0.10fF
C611 a_6375_47# a_6891_47# 0.42fF
C612 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C613 a_32188_47# a_32501_289# 0.00fF
C614 a_32391_413# a_31933_47# 0.12fF
C615 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36515_47# 0.36fF
C616 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10773_47# 1.17fF
C617 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19805_289# 0.46fF
C618 a_16955_47# a_16095_21# 0.02fF
C619 a_40747_47# a_40652_47# 0.13fF
C620 a_41487_21# a_42051_47# 0.30fF
C621 a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.36fF
C622 a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.02fF
C623 a_30167_47# a_30732_47# 0.01fF
C624 a_40397_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C625 a_32848_47# a_31767_47# 0.27fF
C626 a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.02fF
C627 a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.71fF
C628 a_2309_47# a_3399_21# 0.10fF
C629 a_15617_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C630 a_2877_289# a_2659_47# 0.50fF
C631 a_13457_289# a_13804_47# 0.13fF
C632 a_40397_47# a_40747_47# 0.49fF
C633 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[11]/Q 0.12fF
C634 a_32957_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C635 a_38536_47# a_38739_413# 0.02fF
C636 a_18145_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.01fF
C637 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.73fF
C638 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32501_289# 0.46fF
C639 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24037_289# 0.10fF
C640 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16274_47# 0.01fF
C641 a_36515_47# a_37255_21# 0.02fF
C642 a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.63fF
C643 a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.71fF
C644 a_33883_47# a_33023_21# 0.02fF
C645 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20506_47# 0.01fF
C646 a_15573_289# a_15355_47# 0.50fF
C647 a_15005_47# a_16095_21# 0.10fF
C648 a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.71fF
C649 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7810_47# 0.01fF
C650 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3224_47# 0.05fF
C651 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13144_47# 0.53fF
C652 a_25840_47# a_26043_413# 0.02fF
C653 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/D 1.68fF
C654 a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.36fF
C655 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30275_413# 0.01fF
C656 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6541_47# 1.17fF
C657 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C658 a_38536_47# a_38631_47# 0.13fF
C659 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41474_413# 0.01fF
C660 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_11028_47# 0.01fF
C661 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[12]/Q 0.11fF
C662 a_16659_47# a_15920_47# 0.00fF
C663 a_15463_413# a_15355_47# 0.21fF
C664 a_16659_47# a_17121_47# 0.01fF
C665 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15920_47# 0.05fF
C666 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30385_289# 0.10fF
C667 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4993_289# 0.10fF
C668 a_4259_47# a_4775_47# 0.42fF
C669 a_20891_47# a_21353_47# 0.01fF
C670 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22622_47# 0.01fF
C671 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41312_47# 0.68fF
C672 a_17121_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.08fF
C673 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36420_47# 0.53fF
C674 a_39371_21# a_40231_47# 0.02fF
C675 a_26043_413# a_26153_289# 0.23fF
C676 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13239_47# 0.36fF
C677 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31933_47# 0.08fF
C678 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36165_47# 0.65fF
C679 a_35999_47# a_36733_289# 0.16fF
C680 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_3578_47# 0.01fF
C681 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.01fF
C682 a_28616_47# a_28159_413# 0.01fF
C683 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.63fF
C684 a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C685 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32188_47# 0.06fF
C686 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17579_413# 0.17fF
C687 a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.27fF
C688 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21811_413# 0.17fF
C689 a_15005_47# a_15573_289# 0.41fF
C690 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25935_47# 0.36fF
C691 a_28269_289# a_28616_47# 0.13fF
C692 a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C693 a_12889_47# a_13239_47# 0.49fF
C694 a_18775_47# a_19071_47# 0.07fF
C695 a_33587_47# a_34049_47# 0.01fF
C696 a_31767_47# a_31933_47# 1.60fF
C697 a_39935_47# a_40397_47# 0.01fF
C698 a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.71fF
C699 a_10311_47# a_10607_47# 0.07fF
C700 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.17fF
C701 a_27535_47# a_28051_47# 0.42fF
C702 a_15463_413# a_15005_47# 0.12fF
C703 a_15260_47# a_15573_289# 0.00fF
C704 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35703_47# 0.09fF
C705 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8912_47# 0.06fF
C706 a_34617_289# a_35139_21# 0.03fF
C707 a_34049_47# a_34964_47# 0.29fF
C708 a_25419_47# a_25585_47# 1.60fF
C709 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2877_289# 0.10fF
C710 a_2143_47# a_2659_47# 0.42fF
C711 a_12723_47# a_13804_47# 0.27fF
C712 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13979_21# 0.22fF
C713 a_15260_47# a_15463_413# 0.02fF
C714 a_11688_47# a_11231_413# 0.01fF
C715 a_19492_47# a_19695_413# 0.02fF
C716 a_22377_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C717 a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.71fF
C718 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12889_47# 1.17fF
C719 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_35318_47# 0.01fF
C720 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5449_47# 0.01fF
C721 a_14839_47# a_15355_47# 0.42fF
C722 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.12fF
C723 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.06fF
C724 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38739_413# 0.17fF
C725 a_18036_47# a_17579_413# 0.01fF
C726 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# 0.63fF
C727 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11850_413# 0.01fF
C728 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37255_21# 0.73fF
C729 a_22268_47# a_21811_413# 0.01fF
C730 a_32391_413# a_32501_289# 0.23fF
C731 a_8491_47# a_8195_47# 0.07fF
C732 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_193_47# 0.04fF
C733 a_41312_47# a_42051_47# 0.00fF
C734 a_40747_47# a_40855_413# 0.21fF
C735 a_23819_47# a_23915_47# 0.07fF
C736 a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[17]/Q 0.36fF
C737 a_4259_47# a_4425_47# 1.60fF
C738 a_30907_21# a_30732_47# 0.62fF
C739 a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.05fF
C740 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4680_47# 0.06fF
C741 a_805_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C742 a_40397_47# a_41487_21# 0.10fF
C743 a_40965_289# a_40747_47# 0.50fF
C744 a_24037_289# a_23724_47# 0.00fF
C745 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_29651_47# 0.99fF
C746 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38631_47# 0.36fF
C747 a_6891_47# a_6987_47# 0.07fF
C748 a_6796_47# a_6999_413# 0.02fF
C749 a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C750 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18036_47# 0.68fF
C751 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22268_47# 0.68fF
C752 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# 0.27fF
C753 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13457_289# 0.10fF
C754 a_36515_47# a_37080_47# 0.01fF
C755 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.08fF
C756 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17567_47# 0.02fF
C757 a_19683_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.02fF
C758 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21799_47# 0.02fF
C759 a_6079_47# a_6375_47# 0.07fF
C760 a_38739_413# a_38631_47# 0.21fF
C761 a_38727_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.02fF
C762 a_14839_47# a_15005_47# 1.60fF
C763 a_193_47# a_761_289# 0.41fF
C764 a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.36fF
C765 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9747_21# 0.73fF
C766 a_28051_47# a_28147_47# 0.07fF
C767 a_9572_47# a_10311_47# 0.00fF
C768 a_9007_47# a_9115_413# 0.21fF
C769 a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.63fF
C770 a_32283_47# a_33023_21# 0.02fF
C771 a_11123_47# a_11028_47# 0.13fF
C772 a_11863_21# a_12427_47# 0.30fF
C773 a_39371_21# a_38281_47# 0.10fF
C774 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.27fF
C775 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_42051_47# 0.02fF
C776 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24546_413# 0.01fF
C777 a_2309_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.08fF
C778 a_15260_47# a_14839_47# 0.23fF
C779 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.24fF
C780 a_32188_47# a_32391_413# 0.02fF
C781 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36623_413# 0.01fF
C782 sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 1.27fF
C783 a_25935_47# a_26675_21# 0.02fF
C784 a_16274_47# a_16095_21# 0.04fF
C785 a_16029_47# a_15920_47# 0.04fF
C786 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24384_47# 0.68fF
C787 a_448_47# a_193_47# 0.22fF
C788 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D 0.71fF
C789 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.59fF
C790 a_17471_47# a_17376_47# 0.13fF
C791 a_18211_21# a_18775_47# 0.30fF
C792 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36733_289# 0.10fF
C793 a_21703_47# a_21608_47# 0.13fF
C794 a_22443_21# a_23007_47# 0.30fF
C795 a_25840_47# a_25419_47# 0.23fF
C796 a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.24fF
C797 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D 0.01fF
C798 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32391_413# 0.17fF
C799 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.11fF
C800 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26675_21# 0.73fF
C801 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5515_21# 0.73fF
C802 a_27701_47# a_27956_47# 0.22fF
C803 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.01fF
C804 a_1108_47# a_651_413# 0.01fF
C805 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38281_47# 0.08fF
C806 a_31767_47# a_32501_289# 0.16fF
C807 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_31933_47# 0.65fF
C808 sky130_fd_sc_hd__dfrbp_1_0[13]/Q sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.12fF
C809 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# 0.27fF
C810 a_34964_47# a_34507_413# 0.01fF
C811 a_27535_47# a_28791_21# 0.12fF
C812 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28051_47# 0.09fF
C813 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34304_47# 0.06fF
C814 sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.08fF
C815 sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.08fF
C816 a_34617_289# a_34964_47# 0.13fF
C817 a_10773_47# a_11028_47# 0.22fF
C818 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_25585_47# 0.65fF
C819 a_25419_47# a_26153_289# 0.16fF
C820 a_19805_289# a_19695_413# 0.23fF
C821 a_38115_47# a_38281_47# 1.60fF
C822 a_34661_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C823 a_23303_47# a_23724_47# 0.23fF
C824 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34049_47# 1.17fF
C825 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6987_47# 0.02fF
C826 a_761_289# a_1283_21# 0.03fF
C827 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_543_47# 0.30fF
C828 a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.63fF
C829 a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.01fF
C830 a_33883_47# a_34399_47# 0.42fF
C831 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C832 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_8657_47# 1.17fF
C833 a_9007_47# a_9572_47# 0.01fF
C834 a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.71fF
C835 a_8657_47# a_8912_47# 0.22fF
C836 a_40231_47# a_40747_47# 0.42fF
C837 a_17121_47# a_17376_47# 0.22fF
C838 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.27fF
C839 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37242_413# 0.01fF
C840 a_19492_47# a_19237_47# 0.22fF
C841 a_21353_47# a_21608_47# 0.22fF
C842 a_11123_47# a_11863_21# 0.02fF
C843 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11231_413# 0.01fF
C844 a_4775_47# a_4883_413# 0.21fF
C845 a_5340_47# a_6079_47# 0.00fF
C846 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.01fF
C847 a_2564_47# a_2767_413# 0.02fF
C848 a_2659_47# a_2755_47# 0.07fF
C849 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# 0.63fF
C850 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_23007_47# 0.36fF
C851 a_20327_21# a_20152_47# 0.62fF
C852 a_30732_47# a_30894_413# 0.04fF
C853 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37080_47# 0.68fF
C854 sky130_fd_sc_hd__dfrbp_1_0[1]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.11fF
C855 a_651_413# a_543_47# 0.21fF
C856 a_27_47# a_193_47# 1.60fF
C857 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9115_413# 0.01fF
C858 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16095_21# 0.73fF
C859 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17579_413# 0.01fF
C860 a_17471_47# a_18211_21# 0.02fF
C861 a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C862 a_30167_47# a_30072_47# 0.13fF
C863 a_30907_21# a_31471_47# 0.30fF
C864 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.24fF
C865 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21811_413# 0.01fF
C866 a_32188_47# a_31767_47# 0.23fF
C867 a_21703_47# a_22443_21# 0.02fF
C868 a_40965_289# a_41487_21# 0.03fF
C869 a_40397_47# a_41312_47# 0.29fF
C870 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.11fF
C871 a_24037_289# a_23927_413# 0.23fF
C872 a_24493_47# a_24384_47# 0.04fF
C873 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[14]/D 1.68fF
C874 a_24384_47# a_24546_413# 0.04fF
C875 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7618_413# 0.01fF
C876 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14158_47# 0.01fF
C877 a_29817_47# a_30167_47# 0.49fF
C878 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18390_47# 0.01fF
C879 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26500_47# 0.02fF
C880 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.05fF
C881 a_37255_21# a_37080_47# 0.62fF
C882 a_41666_47# a_41487_21# 0.04fF
C883 a_41421_47# a_41312_47# 0.04fF
C884 a_7631_21# a_7456_47# 0.62fF
C885 a_7109_289# a_6796_47# 0.00fF
C886 a_6541_47# a_6999_413# 0.12fF
C887 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4871_47# 0.02fF
C888 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[8]/D 1.68fF
C889 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[10]/D 1.68fF
C890 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.63fF
C891 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_31767_47# 0.99fF
C892 a_38893_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.01fF
C893 a_11341_289# a_11123_47# 0.50fF
C894 a_10773_47# a_11863_21# 0.10fF
C895 a_14543_47# a_14839_47# 0.07fF
C896 a_19805_289# a_20152_47# 0.13fF
C897 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.08fF
C898 a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.36fF
C899 a_3399_21# a_4259_47# 0.02fF
C900 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40652_47# 0.06fF
C901 a_39196_47# a_38281_47# 0.29fF
C902 a_39371_21# a_38849_289# 0.03fF
C903 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24738_47# 0.01fF
C904 a_9225_289# a_9007_47# 0.50fF
C905 a_8657_47# a_9747_21# 0.10fF
C906 a_17689_289# a_17471_47# 0.50fF
C907 a_17121_47# a_18211_21# 0.10fF
C908 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15573_289# 0.46fF
C909 a_39935_47# a_40231_47# 0.07fF
C910 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12042_47# 0.01fF
C911 a_20327_21# a_19237_47# 0.10fF
C912 a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D 0.71fF
C913 a_34399_47# a_34495_47# 0.07fF
C914 a_21921_289# a_21703_47# 0.50fF
C915 a_21353_47# a_22443_21# 0.10fF
C916 a_4775_47# a_5340_47# 0.01fF
C917 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11688_47# 0.05fF
C918 a_25935_47# a_26500_47# 0.01fF
C919 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_15920_47# 0.02fF
C920 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40397_47# 1.17fF
C921 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25123_47# 0.09fF
C922 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11028_47# 0.06fF
C923 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15463_413# 0.17fF
C924 a_27_47# a_1283_21# 0.12fF
C925 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_543_47# 0.09fF
C926 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19695_413# 0.17fF
C927 a_3386_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.01fF
C928 a_27956_47# a_28159_413# 0.02fF
C929 a_16029_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C930 a_1108_47# a_543_47# 0.01fF
C931 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[11]/D 1.68fF
C932 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9572_47# 0.05fF
C933 a_27239_47# a_27535_47# 0.07fF
C934 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[13]/Q 0.11fF
C935 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.53fF
C936 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18036_47# 0.05fF
C937 a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.05fF
C938 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_22268_47# 0.05fF
C939 a_4425_47# a_4883_413# 0.12fF
C940 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26500_47# 0.68fF
C941 a_31086_47# a_30907_21# 0.04fF
C942 a_13804_47# a_13347_413# 0.01fF
C943 a_30841_47# a_30732_47# 0.04fF
C944 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2755_47# 0.02fF
C945 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28051_47# 0.36fF
C946 a_28269_289# a_27956_47# 0.00fF
C947 a_27701_47# a_28159_413# 0.12fF
C948 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_32501_289# 0.10fF
C949 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# 0.27fF
C950 sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C951 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6999_413# 0.17fF
C952 a_10773_47# a_11341_289# 0.41fF
C953 a_27701_47# a_28269_289# 0.41fF
C954 a_27535_47# a_28616_47# 0.27fF
C955 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28791_21# 0.22fF
C956 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34507_413# 0.17fF
C957 a_23819_47# a_24559_21# 0.02fF
C958 a_7109_289# a_7631_21# 0.03fF
C959 a_6541_47# a_7456_47# 0.29fF
C960 a_34049_47# a_34304_47# 0.22fF
C961 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_26153_289# 0.10fF
C962 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38281_47# 0.65fF
C963 a_38115_47# a_38849_289# 0.16fF
C964 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_19071_47# 0.02fF
C965 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34617_289# 0.46fF
C966 sky130_fd_sc_hd__dfrbp_1_0[16]/Q sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.12fF
C967 a_17121_47# a_17689_289# 0.41fF
C968 a_19805_289# a_19237_47# 0.41fF
C969 a_21353_47# a_21921_289# 0.41fF
C970 sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C971 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34399_47# 0.09fF
C972 a_33883_47# a_35139_21# 0.12fF
C973 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_40747_47# 0.09fF
C974 a_40231_47# a_41487_21# 0.12fF
C975 a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.02fF
C976 a_29817_47# a_29355_47# 0.01fF
C977 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# 0.24fF
C978 a_6375_47# a_6796_47# 0.23fF
C979 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_29651_47# 0.02fF
C980 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13335_47# 0.02fF
C981 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C982 a_23303_47# a_23007_47# 0.07fF
C983 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_37819_47# 0.09fF
C984 a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.99fF
C985 a_10607_47# a_11123_47# 0.42fF
C986 a_3399_21# a_3224_47# 0.62fF
C987 a_2877_289# a_2564_47# 0.00fF
C988 a_2309_47# a_2767_413# 0.12fF
C989 a_4993_289# a_4775_47# 0.50fF
C990 a_41312_47# a_40855_413# 0.01fF
C991 a_30732_47# a_31471_47# 0.00fF
C992 a_30167_47# a_30275_413# 0.21fF
C993 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30263_47# 0.02fF
C994 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11863_21# 0.73fF
C995 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.53fF
C996 sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[2]/D 0.08fF
C997 a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.17fF
C998 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20152_47# 0.68fF
C999 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_19237_47# 0.65fF
C1000 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9225_289# 0.10fF
C1001 a_8491_47# a_9007_47# 0.42fF
C1002 a_40965_289# a_41312_47# 0.13fF
C1003 a_37080_47# a_37242_413# 0.04fF
C1004 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_14839_47# 0.99fF
C1005 a_24037_289# a_23819_47# 0.50fF
C1006 a_23469_47# a_24559_21# 0.10fF
C1007 a_16955_47# a_17471_47# 0.42fF
C1008 a_19587_47# a_19071_47# 0.42fF
C1009 a_4425_47# a_5340_47# 0.29fF
C1010 a_21187_47# a_21703_47# 0.42fF
C1011 a_30385_289# a_30167_47# 0.50fF
C1012 a_29817_47# a_30907_21# 0.10fF
C1013 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.11fF
C1014 a_13979_21# a_14543_47# 0.30fF
C1015 a_13239_47# a_13144_47# 0.13fF
C1016 a_24384_47# a_25123_47# 0.00fF
C1017 a_36515_47# a_36420_47# 0.13fF
C1018 a_37255_21# a_37819_47# 0.30fF
C1019 a_24493_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.01fF
C1020 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7456_47# 0.68fF
C1021 a_37189_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.01fF
C1022 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[15]/D 1.68fF
C1023 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_24384_47# 0.05fF
C1024 a_6541_47# a_7109_289# 0.41fF
C1025 a_36165_47# a_36515_47# 0.49fF
C1026 a_15355_47# a_15920_47# 0.01fF
C1027 a_4259_47# a_4680_47# 0.23fF
C1028 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# 0.24fF
C1029 sky130_fd_sc_hd__dfrbp_1_0[18]/Q sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.12fF
C1030 a_12427_47# a_12723_47# 0.07fF
C1031 a_39196_47# a_38849_289# 0.13fF
C1032 sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.08fF
C1033 a_10607_47# a_10773_47# 1.60fF
C1034 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40855_413# 0.17fF
C1035 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26662_413# 0.01fF
C1036 a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D 0.01fF
C1037 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13144_47# 0.06fF
C1038 a_6375_47# a_7631_21# 0.12fF
C1039 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_6891_47# 0.09fF
C1040 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11341_289# 0.46fF
C1041 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.11fF
C1042 a_26675_21# a_26500_47# 0.62fF
C1043 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40965_289# 0.46fF
C1044 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23724_47# 0.06fF
C1045 a_23469_47# a_24037_289# 0.41fF
C1046 a_16955_47# a_17121_47# 1.60fF
C1047 a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[7]/Q 0.36fF
C1048 a_21187_47# a_21353_47# 1.60fF
C1049 a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/Q 0.36fF
C1050 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26854_47# 0.01fF
C1051 a_2877_289# a_3399_21# 0.03fF
C1052 a_2309_47# a_3224_47# 0.29fF
C1053 a_12889_47# a_13144_47# 0.22fF
C1054 sky130_fd_sc_hd__dfrbp_1_0[7]/Q sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.12fF
C1055 a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C1056 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41666_47# 0.01fF
C1057 a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.01fF
C1058 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19237_47# 1.17fF
C1059 a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.71fF
C1060 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# 0.63fF
C1061 a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D 0.01fF
C1062 a_1462_47# a_1283_21# 0.04fF
C1063 a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.68fF
C1064 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28791_21# 0.73fF
C1065 a_28269_289# a_28159_413# 0.23fF
C1066 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[8]/Q 0.27fF
C1067 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41312_47# 0.02fF
C1068 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18198_413# 0.01fF
C1069 a_15573_289# a_16095_21# 0.03fF
C1070 a_15005_47# a_15920_47# 0.29fF
C1071 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_22430_413# 0.01fF
C1072 a_34304_47# a_34507_413# 0.02fF
C1073 a_4425_47# a_4993_289# 0.41fF
C1074 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.01fF
C1075 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9734_413# 0.01fF
C1076 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.11fF
C1077 a_2143_47# a_2564_47# 0.23fF
C1078 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# 0.24fF
C1079 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_28616_47# 0.05fF
C1080 a_33587_47# a_33883_47# 0.07fF
C1081 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13347_413# 0.01fF
C1082 a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[4]/Q 0.27fF
C1083 a_13239_47# a_13979_21# 0.02fF
C1084 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7109_289# 0.46fF
C1085 a_34617_289# a_34304_47# 0.00fF
C1086 a_34049_47# a_34507_413# 0.12fF
C1087 a_40747_47# a_40843_47# 0.07fF
C1088 a_27701_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.08fF
C1089 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_38849_289# 0.10fF
C1090 a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D 0.71fF
C1091 a_23303_47# a_23819_47# 0.42fF
C1092 a_32848_47# a_32283_47# 0.01fF
C1093 a_34049_47# a_34617_289# 0.41fF
C1094 a_4259_47# a_5515_21# 0.12fF
C1095 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4775_47# 0.09fF
C1096 a_33883_47# a_34964_47# 0.27fF
C1097 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35139_21# 0.22fF
C1098 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.11fF
C1099 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_41487_21# 0.19fF
C1100 a_40231_47# a_41312_47# 0.27fF
C1101 a_28725_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.01fF
C1102 a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.36fF
C1103 a_7565_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C1104 a_29651_47# a_28791_21# 0.02fF
C1105 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13979_21# 0.73fF
C1106 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_11219_47# 0.02fF
C1107 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36420_47# 0.06fF
C1108 a_6375_47# a_6541_47# 1.60fF
C1109 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5502_413# 0.01fF
C1110 sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.08fF
C1111 a_18036_47# a_18198_413# 0.04fF
C1112 a_36165_47# a_35703_47# 0.01fF
C1113 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[19]/Q 0.02fF
C1114 a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[3]/Q 0.02fF
C1115 a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[12]/Q 0.36fF
C1116 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[5]/Q 0.11fF
C1117 a_22268_47# a_22430_413# 0.04fF
C1118 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35999_47# 0.02fF
C1119 a_38727_47# a_38631_47# 0.07fF
C1120 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_30429_47# 0.01fF
C1121 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36165_47# 1.17fF
C1122 a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C1123 a_12889_47# a_13979_21# 0.10fF
C1124 a_13457_289# a_13239_47# 0.50fF
C1125 a_2309_47# a_2877_289# 0.41fF
C1126 a_40397_47# a_40652_47# 0.22fF
C1127 a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C1128 a_30385_289# a_30907_21# 0.03fF
C1129 a_29817_47# a_30732_47# 0.29fF
C1130 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_10607_47# 0.99fF
C1131 a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.46fF
C1132 a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.01fF
C1133 a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.02fF
C1134 a_15463_413# a_15573_289# 0.23fF
C1135 a_17471_47# a_17567_47# 0.07fF
C1136 a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D 0.01fF
C1137 a_36515_47# a_36623_413# 0.21fF
C1138 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36611_47# 0.02fF
C1139 a_23303_47# a_23469_47# 1.60fF
C1140 a_37080_47# a_37819_47# 0.00fF
C1141 a_21703_47# a_21799_47# 0.07fF
C1142 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.01fF
C1143 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_4259_47# 0.02fF
C1144 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9115_413# 0.17fF
C1145 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_13804_47# 0.05fF
C1146 a_9007_47# a_9103_47# 0.07fF
C1147 a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D 0.01fF
C1148 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_40231_47# 0.99fF
C1149 a_2143_47# a_3399_21# 0.12fF
C1150 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_2659_47# 0.09fF
C1151 a_8912_47# a_9115_413# 0.02fF
C1152 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# 0.24fF
C1153 a_36165_47# a_37255_21# 0.10fF
C1154 a_36733_289# a_36515_47# 0.50fF
C1155 a_34049_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.08fF
C1156 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[2]/Q 0.27fF
C1157 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13457_289# 0.46fF
C1158 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5694_47# 0.01fF
C1159 a_14839_47# a_16095_21# 0.12fF
C1160 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15355_47# 0.09fF
C1161 a_38536_47# a_38281_47# 0.22fF
C1162 a_26854_47# a_26675_21# 0.04fF
C1163 a_26609_47# a_26500_47# 0.04fF
C1164 a_31933_47# a_32283_47# 0.49fF
C1165 sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[6]/D 0.08fF
C1166 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_14839_47# 0.02fF
C1167 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_6375_47# 0.99fF
C1168 a_39371_21# a_38115_47# 0.12fF
C1169 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_8195_47# 0.01fF
C1170 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_27239_47# 0.09fF
C1171 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23927_413# 0.17fF
C1172 a_12889_47# a_13457_289# 0.41fF
C1173 a_16659_47# a_16955_47# 0.07fF
C1174 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4883_413# 0.17fF
C1175 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_4425_47# 0.65fF
C1176 a_25585_47# a_25935_47# 0.49fF
C1177 a_20891_47# a_21187_47# 0.07fF
C1178 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28778_413# 0.01fF
C1179 sky130_fd_sc_hd__dfrbp_1_0[0]/Q sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.12fF
C1180 a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.63fF
C1181 a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[0]/Q 0.02fF
C1182 a_7456_47# a_7618_413# 0.04fF
C1183 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.08fF
C1184 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_18775_47# 0.09fF
C1185 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23007_47# 0.09fF
C1186 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3333_47# 0.01fF
C1187 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28616_47# 0.68fF
C1188 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/CLK 0.01fF
C1189 a_18211_21# a_19071_47# 0.02fF
C1190 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_42051_47# 0.36fF
C1191 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25585_47# 1.17fF
C1192 a_9747_21# a_10607_47# 0.02fF
C1193 a_27535_47# a_27956_47# 0.23fF
C1194 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# 0.24fF
C1195 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C1196 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_17733_47# 0.01fF
C1197 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# 0.63fF
C1198 a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D 0.71fF
C1199 a_19849_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.01fF
C1200 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_21965_47# 0.01fF
C1201 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_15005_47# 0.65fF
C1202 a_14839_47# a_15573_289# 0.16fF
C1203 a_193_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.33fF
C1204 a_34617_289# a_34507_413# 0.23fF
C1205 a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.01fF
C1206 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9572_47# 0.68fF
C1207 a_2143_47# a_2309_47# 1.60fF
C1208 a_12723_47# a_13239_47# 0.42fF
C1209 a_27535_47# a_27701_47# 1.60fF
C1210 a_4680_47# a_4883_413# 0.02fF
C1211 a_4775_47# a_4871_47# 0.07fF
C1212 a_32848_47# a_33023_21# 0.62fF
C1213 a_11123_47# a_11231_413# 0.21fF
C1214 a_11688_47# a_12427_47# 0.00fF
C1215 a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[1]/Q 0.02fF
C1216 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_34964_47# 0.05fF
C1217 a_20152_47# a_19695_413# 0.01fF
C1218 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.99fF
C1219 a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D 0.71fF
C1220 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_41312_47# 0.05fF
C1221 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30167_47# 0.36fF
C1222 a_1847_47# a_2309_47# 0.01fF
C1223 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.53fF
C1224 a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D 0.01fF
C1225 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_33883_47# 0.99fF
C1226 a_33202_47# a_33023_21# 0.04fF
C1227 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6796_47# 0.01fF
C1228 a_448_47# a_761_289# 0.00fF
C1229 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D 0.01fF
C1230 a_651_413# a_193_47# 0.12fF
C1231 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B 0.09fF
C1232 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_9103_47# 0.02fF
C1233 a_17471_47# a_17579_413# 0.21fF
C1234 a_18036_47# a_18775_47# 0.00fF
C1235 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36623_413# 0.17fF
C1236 a_22268_47# a_23007_47# 0.00fF
C1237 a_21703_47# a_21811_413# 0.21fF
C1238 a_8491_47# a_7631_21# 0.02fF
C1239 a_24559_21# a_25419_47# 0.02fF
C1240 a_40652_47# a_40855_413# 0.02fF
C1241 a_35073_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D 0.01fF
C1242 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19237_47# 0.08fF
C1243 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_12723_47# 0.99fF
C1244 a_21353_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D 0.08fF
C1245 a_39371_21# a_39196_47# 0.62fF
C1246 a_30732_47# a_30275_413# 0.01fF
C1247 sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[14]/Q 0.12fF
C1248 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36733_289# 0.46fF
C1249 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5340_47# 0.68fF
C1250 a_40965_289# a_40652_47# 0.00fF
C1251 a_40397_47# a_40855_413# 0.12fF
C1252 a_35999_47# a_35139_21# 0.02fF
C1253 a_1108_47# a_1270_413# 0.04fF
C1254 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17471_47# 0.36fF
C1255 a_7456_47# a_6999_413# 0.01fF
C1256 a_30385_289# a_30732_47# 0.13fF
C1257 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21703_47# 0.36fF
C1258 a_3963_47# a_4425_47# 0.01fF
C1259 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# 0.44fF
C1260 a_12723_47# a_12889_47# 1.60fF
C1261 a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[15]/Q 0.36fF
C1262 a_40397_47# a_40965_289# 0.41fF
C1263 a_24384_47# a_23927_413# 0.01fF
C1264 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_36777_47# 0.01fF
C1265 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_31767_47# 0.02fF
C1266 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38281_47# 1.17fF
C1267 a_29651_47# a_30167_47# 0.42fF
C1268 a_11341_289# a_11028_47# 0.00fF
C1269 a_10773_47# a_11231_413# 0.12fF
C1270 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[19]/D 1.30fF
C1271 a_26662_413# a_26500_47# 0.04fF
C1272 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_23724_47# 0.53fF
C1273 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_7153_47# 0.01fF
C1274 a_36733_289# a_37255_21# 0.03fF
C1275 a_36165_47# a_37080_47# 0.29fF
C1276 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_1283_21# 0.71fF
C1277 a_5515_21# a_6375_47# 0.02fF
C1278 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[6]/Q 0.27fF
C1279 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9225_289# 0.46fF
C1280 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_25419_47# 0.02fF
C1281 a_9225_289# a_8912_47# 0.00fF
C1282 a_8657_47# a_9115_413# 0.12fF
C1283 a_25840_47# a_25935_47# 0.13fF
C1284 a_27239_47# a_26675_21# 0.30fF
C1285 a_9747_21# a_9572_47# 0.62fF
C1286 a_14158_47# a_13979_21# 0.04fF
C1287 a_13913_47# a_13804_47# 0.04fF
C1288 a_17689_289# a_17376_47# 0.00fF
C1289 a_17121_47# a_17579_413# 0.12fF
C1290 a_19695_413# a_19237_47# 0.12fF
C1291 a_21921_289# a_21608_47# 0.00fF
C1292 a_21353_47# a_21811_413# 0.12fF
C1293 a_11123_47# a_11688_47# 0.01fF
C1294 a_3224_47# a_3386_413# 0.04fF
C1295 a_38739_413# a_38281_47# 0.12fF
C1296 a_38536_47# a_38849_289# 0.00fF
C1297 a_19587_47# a_19492_47# 0.13fF
C1298 a_20327_21# a_20891_47# 0.30fF
C1299 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[5]/D 0.08fF
C1300 a_32501_289# a_32283_47# 0.50fF
C1301 a_31933_47# a_33023_21# 0.10fF
C1302 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# 0.27fF
C1303 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_193_47# 0.65fF
C1304 a_27_47# a_761_289# 0.16fF
C1305 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.22fF
C1306 a_39196_47# a_38115_47# 0.27fF
C1307 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23819_47# 0.36fF
C1308 a_28051_47# a_28791_21# 0.02fF
C1309 a_1108_47# a_193_47# 0.29fF
C1310 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_25840_47# 0.06fF
C1311 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15920_47# 0.68fF
C1312 a_17471_47# a_18036_47# 0.01fF
C1313 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17121_47# 1.17fF
C1314 a_21703_47# a_22268_47# 0.01fF
C1315 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21353_47# 1.17fF
C1316 a_26153_289# a_25935_47# 0.50fF
C1317 a_25585_47# a_26675_21# 0.10fF
C1318 a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.63fF
C1319 a_38281_47# a_38631_47# 0.49fF
C1320 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_16082_413# 0.01fF
C1321 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_20314_413# 0.01fF
C1322 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_29355_47# 0.09fF
C1323 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_4993_289# 0.46fF
C1324 a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D 0.24fF
C1325 a_448_47# a_27_47# 0.23fF
C1326 a_1108_47# a_1847_47# 0.00fF
C1327 a_6891_47# a_6796_47# 0.13fF
C1328 a_7109_289# a_6999_413# 0.23fF
C1329 a_7631_21# a_8195_47# 0.30fF
C1330 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_5037_47# 0.01fF
C1331 sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[3]/D 0.08fF
C1332 a_13804_47# a_13966_413# 0.04fF
C1333 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26153_289# 0.46fF
C1334 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[18]/Q 0.11fF
C1335 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_27956_47# 0.53fF
C1336 sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.08fF
C1337 a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D 0.01fF
C1338 a_11341_289# a_11863_21# 0.03fF
C1339 a_10773_47# a_11688_47# 0.29fF
C1340 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28970_47# 0.01fF
C1341 a_27535_47# a_28269_289# 0.16fF
C1342 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_27701_47# 0.65fF
C1343 a_30167_47# a_30263_47# 0.07fF
C1344 a_32188_47# a_32283_47# 0.13fF
C1345 a_33587_47# a_33023_21# 0.30fF
C1346 a_193_47# a_543_47# 0.49fF
C1347 a_13239_47# a_13335_47# 0.07fF
C1348 a_33883_47# a_34304_47# 0.23fF
C1349 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# 0.24fF
C1350 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_23469_47# 1.17fF
C1351 a_9225_289# a_9747_21# 0.03fF
C1352 a_8657_47# a_9572_47# 0.29fF
C1353 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30907_21# 0.73fF
C1354 a_40231_47# a_40652_47# 0.23fF
C1355 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# 0.21fF
C1356 a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D 0.71fF
C1357 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[16]/D 1.68fF
C1358 a_17689_289# a_18211_21# 0.03fF
C1359 a_17121_47# a_18036_47# 0.29fF
C1360 a_20152_47# a_19237_47# 0.29fF
C1361 a_21921_289# a_22443_21# 0.03fF
C1362 a_21353_47# a_22268_47# 0.29fF
C1363 a_10607_47# a_11028_47# 0.23fF
C1364 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# 0.24fF
C1365 a_3224_47# a_2767_413# 0.01fF
C1366 a_33883_47# a_34049_47# 1.60fF
C1367 a_4993_289# a_4680_47# 0.00fF
C1368 a_5515_21# a_5340_47# 0.62fF
C1369 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# 0.27fF
C1370 a_19587_47# a_20327_21# 0.02fF
C1371 a_29651_47# a_29355_47# 0.07fF
C1372 a_40231_47# a_40397_47# 1.60fF
C1373 a_39196_47# a_39358_413# 0.04fF
C1374 a_41666_47# GND 0.01fF
C1375 a_41421_47# GND 0.01fF
C1376 sky130_fd_sc_hd__dfrbp_1_0[19]/Q GND 0.32fF
C1377 a_41009_47# GND 0.01fF
C1378 a_40843_47# GND 0.03fF
C1379 a_39550_47# GND -0.01fF
C1380 a_39305_47# GND -0.01fF
C1381 a_40855_413# GND 0.11fF
C1382 a_40652_47# GND 0.23fF
C1383 a_42051_47# GND 0.45fF
C1384 a_41312_47# GND 0.79fF
C1385 a_41487_21# GND 1.50fF
C1386 a_40747_47# GND 0.68fF
C1387 a_40965_289# GND 0.58fF
C1388 a_40397_47# GND 0.16fF
C1389 sky130_fd_sc_hd__dfrbp_1_0[19]/D GND 0.04fF
C1390 a_40231_47# GND 0.42fF
C1391 sky130_fd_sc_hd__dfrbp_1_0[18]/Q GND 0.13fF
C1392 a_38893_47# GND -0.01fF
C1393 a_37434_47# GND 0.01fF
C1394 a_37189_47# GND 0.01fF
C1395 a_38739_413# GND 0.09fF
C1396 a_38536_47# GND 0.08fF
C1397 a_39935_47# GND 0.30fF
C1398 a_39196_47# GND -0.41fF
C1399 a_39371_21# GND -0.79fF
C1400 a_38631_47# GND 0.43fF
C1401 a_38849_289# GND -0.44fF
C1402 a_38281_47# GND 0.47fF
C1403 sky130_fd_sc_hd__dfrbp_1_0[18]/D GND 0.58fF
C1404 a_38115_47# GND 0.70fF
C1405 sky130_fd_sc_hd__dfrbp_1_0[17]/Q GND 0.32fF
C1406 a_36777_47# GND 0.01fF
C1407 a_36611_47# GND 0.03fF
C1408 a_35318_47# GND -0.01fF
C1409 a_35073_47# GND -0.01fF
C1410 a_36623_413# GND 0.11fF
C1411 a_36420_47# GND 0.23fF
C1412 a_37819_47# GND 0.45fF
C1413 a_37080_47# GND 0.79fF
C1414 a_37255_21# GND 1.50fF
C1415 a_36515_47# GND 0.68fF
C1416 a_36733_289# GND 0.58fF
C1417 a_36165_47# GND 0.16fF
C1418 sky130_fd_sc_hd__dfrbp_1_0[17]/D GND 0.04fF
C1419 a_35999_47# GND 0.42fF
C1420 sky130_fd_sc_hd__dfrbp_1_0[16]/Q GND 0.13fF
C1421 a_34661_47# GND -0.01fF
C1422 a_33202_47# GND 0.01fF
C1423 a_32957_47# GND 0.01fF
C1424 a_34507_413# GND 0.09fF
C1425 a_34304_47# GND 0.08fF
C1426 a_35703_47# GND 0.30fF
C1427 a_34964_47# GND -0.39fF
C1428 a_35139_21# GND -0.75fF
C1429 a_34399_47# GND 0.46fF
C1430 a_34617_289# GND -0.43fF
C1431 a_34049_47# GND 0.64fF
C1432 sky130_fd_sc_hd__dfrbp_1_0[16]/D GND 0.58fF
C1433 a_33883_47# GND 0.75fF
C1434 sky130_fd_sc_hd__dfrbp_1_0[15]/Q GND 0.32fF
C1435 a_32545_47# GND 0.01fF
C1436 a_32379_47# GND 0.03fF
C1437 a_31086_47# GND -0.01fF
C1438 a_30841_47# GND -0.01fF
C1439 a_32391_413# GND 0.11fF
C1440 a_32188_47# GND 0.23fF
C1441 a_33587_47# GND 0.45fF
C1442 a_32848_47# GND 0.79fF
C1443 a_33023_21# GND 1.50fF
C1444 a_32283_47# GND 0.68fF
C1445 a_32501_289# GND 0.58fF
C1446 a_31933_47# GND 0.16fF
C1447 sky130_fd_sc_hd__dfrbp_1_0[15]/D GND 0.04fF
C1448 a_31767_47# GND 0.42fF
C1449 sky130_fd_sc_hd__dfrbp_1_0[14]/Q GND 0.13fF
C1450 a_30429_47# GND -0.01fF
C1451 a_28970_47# GND 0.01fF
C1452 a_28725_47# GND 0.01fF
C1453 a_30275_413# GND 0.09fF
C1454 a_30072_47# GND 0.08fF
C1455 a_31471_47# GND 0.30fF
C1456 a_30732_47# GND -0.60fF
C1457 a_30907_21# GND -0.71fF
C1458 a_30167_47# GND 0.46fF
C1459 a_30385_289# GND -0.59fF
C1460 a_29817_47# GND 0.70fF
C1461 sky130_fd_sc_hd__dfrbp_1_0[14]/D GND 0.58fF
C1462 a_29651_47# GND 0.80fF
C1463 sky130_fd_sc_hd__dfrbp_1_0[13]/Q GND 0.32fF
C1464 a_28313_47# GND 0.01fF
C1465 a_28147_47# GND 0.03fF
C1466 a_26854_47# GND -0.01fF
C1467 a_26609_47# GND -0.01fF
C1468 a_28159_413# GND 0.11fF
C1469 a_27956_47# GND 0.23fF
C1470 a_29355_47# GND 0.45fF
C1471 a_28616_47# GND 0.79fF
C1472 a_28791_21# GND 1.50fF
C1473 a_28051_47# GND 0.68fF
C1474 a_28269_289# GND 0.58fF
C1475 a_27701_47# GND 0.16fF
C1476 sky130_fd_sc_hd__dfrbp_1_0[13]/D GND 0.04fF
C1477 a_27535_47# GND 0.42fF
C1478 sky130_fd_sc_hd__dfrbp_1_0[12]/Q GND 0.13fF
C1479 a_26197_47# GND -0.01fF
C1480 a_24738_47# GND 0.01fF
C1481 a_24493_47# GND 0.01fF
C1482 a_26043_413# GND 0.09fF
C1483 a_25840_47# GND 0.08fF
C1484 a_27239_47# GND 0.30fF
C1485 a_26500_47# GND -0.52fF
C1486 a_26675_21# GND -0.67fF
C1487 a_25935_47# GND 0.46fF
C1488 a_26153_289# GND 0.40fF
C1489 a_25585_47# GND 0.76fF
C1490 sky130_fd_sc_hd__dfrbp_1_0[12]/D GND 0.59fF
C1491 a_25419_47# GND 0.96fF
C1492 sky130_fd_sc_hd__dfrbp_1_0[11]/Q GND 0.32fF
C1493 a_24081_47# GND 0.01fF
C1494 a_23915_47# GND 0.03fF
C1495 a_22622_47# GND -0.01fF
C1496 a_22377_47# GND -0.01fF
C1497 a_23927_413# GND 0.11fF
C1498 a_23724_47# GND 0.23fF
C1499 a_25123_47# GND 0.45fF
C1500 a_24384_47# GND 0.79fF
C1501 a_24559_21# GND 1.50fF
C1502 a_23819_47# GND 0.68fF
C1503 a_24037_289# GND 0.58fF
C1504 a_23469_47# GND 0.16fF
C1505 sky130_fd_sc_hd__dfrbp_1_0[11]/D GND 0.04fF
C1506 a_23303_47# GND 0.42fF
C1507 sky130_fd_sc_hd__dfrbp_1_0[10]/Q GND 0.13fF
C1508 a_21965_47# GND -0.01fF
C1509 a_20506_47# GND 0.01fF
C1510 a_20261_47# GND 0.01fF
C1511 a_21811_413# GND 0.09fF
C1512 a_21608_47# GND 0.08fF
C1513 a_23007_47# GND 0.30fF
C1514 a_22268_47# GND -0.30fF
C1515 a_22443_21# GND -0.63fF
C1516 a_21703_47# GND 0.46fF
C1517 a_21921_289# GND 0.40fF
C1518 a_21353_47# GND 0.84fF
C1519 sky130_fd_sc_hd__dfrbp_1_0[10]/D GND 0.59fF
C1520 a_21187_47# GND 1.08fF
C1521 sky130_fd_sc_hd__dfrbp_1_0[9]/Q GND 0.32fF
C1522 a_19849_47# GND 0.01fF
C1523 a_19683_47# GND 0.03fF
C1524 a_18390_47# GND -0.01fF
C1525 a_18145_47# GND -0.01fF
C1526 a_19695_413# GND 0.11fF
C1527 a_19492_47# GND 0.23fF
C1528 a_20891_47# GND 0.45fF
C1529 a_20152_47# GND 0.79fF
C1530 a_20327_21# GND 1.50fF
C1531 a_19587_47# GND 0.68fF
C1532 a_19805_289# GND 0.58fF
C1533 a_19237_47# GND 0.16fF
C1534 sky130_fd_sc_hd__dfrbp_1_0[9]/D GND 0.04fF
C1535 a_19071_47# GND 0.42fF
C1536 sky130_fd_sc_hd__dfrbp_1_0[8]/Q GND 0.13fF
C1537 a_16274_47# GND 0.01fF
C1538 a_16029_47# GND 0.01fF
C1539 a_17579_413# GND 0.09fF
C1540 a_17376_47# GND 0.08fF
C1541 a_18775_47# GND 0.30fF
C1542 a_18036_47# GND -0.23fF
C1543 a_18211_21# GND -0.59fF
C1544 a_17471_47# GND 0.46fF
C1545 a_17689_289# GND 0.40fF
C1546 a_17121_47# GND 0.88fF
C1547 sky130_fd_sc_hd__dfrbp_1_0[8]/D GND 0.59fF
C1548 a_16955_47# GND 1.15fF
C1549 sky130_fd_sc_hd__dfrbp_1_0[7]/Q GND 0.32fF
C1550 a_15617_47# GND 0.01fF
C1551 a_15451_47# GND 0.03fF
C1552 a_14158_47# GND -0.01fF
C1553 a_13913_47# GND -0.01fF
C1554 a_15463_413# GND 0.11fF
C1555 a_15260_47# GND 0.23fF
C1556 a_16659_47# GND 0.45fF
C1557 a_15920_47# GND 0.79fF
C1558 a_16095_21# GND 1.50fF
C1559 a_15355_47# GND 0.68fF
C1560 a_15573_289# GND 0.58fF
C1561 a_15005_47# GND 0.16fF
C1562 sky130_fd_sc_hd__dfrbp_1_0[7]/D GND 0.04fF
C1563 a_14839_47# GND 0.42fF
C1564 sky130_fd_sc_hd__dfrbp_1_0[6]/Q GND 0.13fF
C1565 a_12042_47# GND 0.01fF
C1566 a_11797_47# GND 0.01fF
C1567 a_13347_413# GND 0.09fF
C1568 a_13144_47# GND 0.08fF
C1569 a_14543_47# GND 0.30fF
C1570 a_13804_47# GND -0.23fF
C1571 a_13979_21# GND -0.55fF
C1572 a_13239_47# GND 0.46fF
C1573 a_13457_289# GND 0.40fF
C1574 a_12889_47# GND 0.91fF
C1575 sky130_fd_sc_hd__dfrbp_1_0[6]/D GND 0.59fF
C1576 a_12723_47# GND 1.19fF
C1577 sky130_fd_sc_hd__dfrbp_1_0[5]/Q GND 0.32fF
C1578 a_11385_47# GND 0.01fF
C1579 a_11219_47# GND 0.03fF
C1580 a_9926_47# GND -0.01fF
C1581 a_9681_47# GND -0.01fF
C1582 a_11231_413# GND 0.11fF
C1583 a_11028_47# GND 0.23fF
C1584 a_12427_47# GND 0.45fF
C1585 a_11688_47# GND 0.79fF
C1586 a_11863_21# GND 1.50fF
C1587 a_11123_47# GND 0.68fF
C1588 a_11341_289# GND 0.58fF
C1589 a_10773_47# GND 0.16fF
C1590 sky130_fd_sc_hd__dfrbp_1_0[5]/D GND 0.04fF
C1591 a_10607_47# GND 0.42fF
C1592 sky130_fd_sc_hd__dfrbp_1_0[4]/Q GND 0.13fF
C1593 a_7810_47# GND 0.01fF
C1594 a_7565_47# GND 0.01fF
C1595 a_9115_413# GND 0.09fF
C1596 a_8912_47# GND 0.08fF
C1597 a_10311_47# GND 0.30fF
C1598 a_9572_47# GND -0.20fF
C1599 a_9747_21# GND -0.51fF
C1600 a_9007_47# GND 0.46fF
C1601 a_9225_289# GND 0.40fF
C1602 a_8657_47# GND 0.98fF
C1603 sky130_fd_sc_hd__dfrbp_1_0[4]/D GND 0.58fF
C1604 a_8491_47# GND 1.19fF
C1605 sky130_fd_sc_hd__dfrbp_1_0[3]/Q GND 0.32fF
C1606 a_7153_47# GND 0.01fF
C1607 a_6987_47# GND 0.03fF
C1608 a_5694_47# GND -0.01fF
C1609 a_5449_47# GND -0.01fF
C1610 a_6999_413# GND 0.11fF
C1611 a_6796_47# GND 0.23fF
C1612 a_8195_47# GND 0.45fF
C1613 a_7456_47# GND 0.79fF
C1614 a_7631_21# GND 1.50fF
C1615 a_6891_47# GND 0.68fF
C1616 a_7109_289# GND 0.58fF
C1617 a_6541_47# GND 0.16fF
C1618 sky130_fd_sc_hd__dfrbp_1_0[3]/D GND 0.04fF
C1619 a_6375_47# GND 0.42fF
C1620 sky130_fd_sc_hd__dfrbp_1_0[2]/Q GND 0.13fF
C1621 a_3578_47# GND 0.01fF
C1622 a_3333_47# GND 0.01fF
C1623 a_4883_413# GND 0.09fF
C1624 a_4680_47# GND 0.08fF
C1625 a_6079_47# GND 0.30fF
C1626 a_5340_47# GND -0.35fF
C1627 a_5515_21# GND -0.49fF
C1628 a_4775_47# GND 0.46fF
C1629 a_4993_289# GND 0.40fF
C1630 a_4425_47# GND 0.98fF
C1631 sky130_fd_sc_hd__dfrbp_1_0[2]/D GND 0.58fF
C1632 a_4259_47# GND 1.19fF
C1633 sky130_fd_sc_hd__dfrbp_1_0[1]/Q GND 0.32fF
C1634 a_2921_47# GND 0.01fF
C1635 a_2755_47# GND 0.03fF
C1636 a_1462_47# GND -0.01fF
C1637 a_1217_47# GND -0.01fF
C1638 a_2767_413# GND 0.11fF
C1639 a_2564_47# GND 0.23fF
C1640 a_3963_47# GND 0.45fF
C1641 a_3224_47# GND 0.79fF
C1642 a_3399_21# GND 1.50fF
C1643 a_2659_47# GND 0.68fF
C1644 a_2877_289# GND 0.58fF
C1645 a_2309_47# GND 0.16fF
C1646 sky130_fd_sc_hd__dfrbp_1_0[1]/D GND 0.04fF
C1647 a_2143_47# GND 0.42fF
C1648 sky130_fd_sc_hd__dfrbp_1_0[0]/Q GND 0.13fF
C1649 a_651_413# GND 0.09fF
C1650 a_448_47# GND 0.08fF
C1651 a_1847_47# GND 0.30fF
C1652 a_1108_47# GND -0.51fF
C1653 a_1283_21# GND -0.44fF
C1654 a_543_47# GND 0.46fF
C1655 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B GND 0.20fF
C1656 a_761_289# GND 0.40fF
C1657 a_193_47# GND 0.98fF
C1658 sky130_fd_sc_hd__dfrbp_1_0[0]/D GND 0.58fF
C1659 a_27_47# GND 1.76fF
C1660 sky130_fd_sc_hd__dfrbp_1_0[0]/CLK GND 0.41fF
C1661 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t78 GND 0.01fF
C1662 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t5 GND 0.01fF
C1663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n0 GND 0.04fF $ **FLOATING
C1664 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t201 GND 0.02fF
C1665 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1 GND 0.02fF $ **FLOATING
C1666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n2 GND 0.03fF $ **FLOATING
C1667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n3 GND 0.07fF $ **FLOATING
C1668 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n4 GND 0.02fF $ **FLOATING
C1669 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n5 GND 0.04fF $ **FLOATING
C1670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n6 GND 0.02fF $ **FLOATING
C1671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n7 GND 0.05fF $ **FLOATING
C1672 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n8 GND 0.02fF $ **FLOATING
C1673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n9 GND 0.03fF $ **FLOATING
C1674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n10 GND 0.05fF $ **FLOATING
C1675 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n11 GND 0.02fF $ **FLOATING
C1676 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n12 GND 0.05fF $ **FLOATING
C1677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n13 GND 0.02fF $ **FLOATING
C1678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n14 GND 0.05fF $ **FLOATING
C1679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n15 GND 0.02fF $ **FLOATING
C1680 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t220 GND 0.02fF
C1681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t24 GND 0.01fF
C1682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n16 GND 0.10fF $ **FLOATING
C1683 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n17 GND 0.02fF $ **FLOATING
C1684 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n18 GND 0.05fF $ **FLOATING
C1685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n19 GND 0.04fF $ **FLOATING
C1686 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n20 GND 0.10fF $ **FLOATING
C1687 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n21 GND 0.21fF $ **FLOATING
C1688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n22 GND 0.02fF $ **FLOATING
C1689 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n23 GND 0.05fF $ **FLOATING
C1690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n24 GND 0.06fF $ **FLOATING
C1691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n25 GND 0.02fF $ **FLOATING
C1692 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n26 GND 0.04fF $ **FLOATING
C1693 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n27 GND 0.06fF $ **FLOATING
C1694 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t221 GND 0.02fF
C1695 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n28 GND 0.06fF $ **FLOATING
C1696 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n29 GND 0.05fF $ **FLOATING
C1697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t83 GND 0.01fF
C1698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n30 GND 0.03fF $ **FLOATING
C1699 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n31 GND 0.05fF $ **FLOATING
C1700 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n32 GND 0.02fF $ **FLOATING
C1701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n33 GND 0.04fF $ **FLOATING
C1702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n34 GND 0.06fF $ **FLOATING
C1703 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n35 GND 0.02fF $ **FLOATING
C1704 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n36 GND 0.04fF $ **FLOATING
C1705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n37 GND 0.06fF $ **FLOATING
C1706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t191 GND 0.01fF
C1707 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t222 GND 0.02fF
C1708 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n38 GND 0.04fF $ **FLOATING
C1709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n39 GND 0.04fF $ **FLOATING
C1710 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n40 GND 0.02fF $ **FLOATING
C1711 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n41 GND 0.03fF $ **FLOATING
C1712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n42 GND 0.06fF $ **FLOATING
C1713 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n43 GND 0.02fF $ **FLOATING
C1714 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n44 GND 0.05fF $ **FLOATING
C1715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n45 GND 0.06fF $ **FLOATING
C1716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n46 GND 0.02fF $ **FLOATING
C1717 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n47 GND 0.05fF $ **FLOATING
C1718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n48 GND 0.06fF $ **FLOATING
C1719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n49 GND 0.02fF $ **FLOATING
C1720 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n50 GND 0.05fF $ **FLOATING
C1721 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n51 GND 0.06fF $ **FLOATING
C1722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t209 GND 0.04fF
C1723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n52 GND 0.09fF $ **FLOATING
C1724 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n53 GND 0.02fF $ **FLOATING
C1725 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n54 GND 0.03fF $ **FLOATING
C1726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n55 GND 0.06fF $ **FLOATING
C1727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n56 GND 0.02fF $ **FLOATING
C1728 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n57 GND 0.04fF $ **FLOATING
C1729 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n58 GND 0.06fF $ **FLOATING
C1730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t176 GND 0.01fF
C1731 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t208 GND 0.01fF
C1732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n59 GND 0.04fF $ **FLOATING
C1733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n60 GND 0.05fF $ **FLOATING
C1734 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n61 GND 0.02fF $ **FLOATING
C1735 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n62 GND 0.04fF $ **FLOATING
C1736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n63 GND 0.06fF $ **FLOATING
C1737 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n64 GND 0.02fF $ **FLOATING
C1738 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n65 GND 0.04fF $ **FLOATING
C1739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n66 GND 0.06fF $ **FLOATING
C1740 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n67 GND 0.02fF $ **FLOATING
C1741 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n68 GND 0.05fF $ **FLOATING
C1742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n69 GND 0.06fF $ **FLOATING
C1743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n70 GND 0.02fF $ **FLOATING
C1744 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n71 GND 0.05fF $ **FLOATING
C1745 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n72 GND 0.06fF $ **FLOATING
C1746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n73 GND 0.02fF $ **FLOATING
C1747 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n74 GND 0.05fF $ **FLOATING
C1748 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n75 GND 0.06fF $ **FLOATING
C1749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t25 GND 0.02fF
C1750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n76 GND 0.07fF $ **FLOATING
C1751 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n77 GND 0.02fF $ **FLOATING
C1752 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n78 GND 0.03fF $ **FLOATING
C1753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n79 GND 0.06fF $ **FLOATING
C1754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n80 GND 0.02fF $ **FLOATING
C1755 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n81 GND 0.04fF $ **FLOATING
C1756 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n82 GND 0.06fF $ **FLOATING
C1757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n83 GND 0.02fF $ **FLOATING
C1758 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n84 GND 0.05fF $ **FLOATING
C1759 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n85 GND 0.06fF $ **FLOATING
C1760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t1 GND 0.01fF
C1761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t238 GND 0.01fF
C1762 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n86 GND 0.04fF $ **FLOATING
C1763 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n87 GND 0.05fF $ **FLOATING
C1764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n88 GND 0.02fF $ **FLOATING
C1765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n89 GND 0.03fF $ **FLOATING
C1766 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n90 GND 0.06fF $ **FLOATING
C1767 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n91 GND 0.02fF $ **FLOATING
C1768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n92 GND 0.05fF $ **FLOATING
C1769 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n93 GND 0.06fF $ **FLOATING
C1770 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n94 GND 0.02fF $ **FLOATING
C1771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n95 GND 0.05fF $ **FLOATING
C1772 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n96 GND 0.06fF $ **FLOATING
C1773 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t153 GND 0.02fF
C1774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t129 GND 0.01fF
C1775 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n97 GND 0.10fF $ **FLOATING
C1776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n98 GND 0.04fF $ **FLOATING
C1777 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n99 GND 0.02fF $ **FLOATING
C1778 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n100 GND 0.03fF $ **FLOATING
C1779 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n101 GND 0.06fF $ **FLOATING
C1780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n102 GND 0.02fF $ **FLOATING
C1781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n103 GND 0.05fF $ **FLOATING
C1782 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n104 GND 0.06fF $ **FLOATING
C1783 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n105 GND 0.02fF $ **FLOATING
C1784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n106 GND 0.05fF $ **FLOATING
C1785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n107 GND 0.06fF $ **FLOATING
C1786 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n108 GND 0.02fF $ **FLOATING
C1787 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n109 GND 0.04fF $ **FLOATING
C1788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n110 GND 0.06fF $ **FLOATING
C1789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t154 GND 0.02fF
C1790 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n111 GND 0.06fF $ **FLOATING
C1791 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n112 GND 0.05fF $ **FLOATING
C1792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t108 GND 0.01fF
C1793 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n113 GND 0.03fF $ **FLOATING
C1794 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n114 GND 0.05fF $ **FLOATING
C1795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n115 GND 0.02fF $ **FLOATING
C1796 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n116 GND 0.04fF $ **FLOATING
C1797 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n117 GND 0.06fF $ **FLOATING
C1798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n118 GND 0.02fF $ **FLOATING
C1799 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n119 GND 0.04fF $ **FLOATING
C1800 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n120 GND 0.06fF $ **FLOATING
C1801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t164 GND 0.01fF
C1802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t152 GND 0.02fF
C1803 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n121 GND 0.04fF $ **FLOATING
C1804 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n122 GND 0.04fF $ **FLOATING
C1805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n123 GND 0.02fF $ **FLOATING
C1806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n124 GND 0.03fF $ **FLOATING
C1807 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n125 GND 0.06fF $ **FLOATING
C1808 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n126 GND 0.02fF $ **FLOATING
C1809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n127 GND 0.05fF $ **FLOATING
C1810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n128 GND 0.06fF $ **FLOATING
C1811 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n129 GND 0.02fF $ **FLOATING
C1812 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n130 GND 0.05fF $ **FLOATING
C1813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n131 GND 0.06fF $ **FLOATING
C1814 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n132 GND 0.02fF $ **FLOATING
C1815 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n133 GND 0.05fF $ **FLOATING
C1816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n134 GND 0.06fF $ **FLOATING
C1817 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t56 GND 0.04fF
C1818 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n135 GND 0.09fF $ **FLOATING
C1819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n136 GND 0.02fF $ **FLOATING
C1820 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n137 GND 0.03fF $ **FLOATING
C1821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n138 GND 0.06fF $ **FLOATING
C1822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n139 GND 0.02fF $ **FLOATING
C1823 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n140 GND 0.04fF $ **FLOATING
C1824 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n141 GND 0.06fF $ **FLOATING
C1825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t180 GND 0.01fF
C1826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t2 GND 0.01fF
C1827 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n142 GND 0.04fF $ **FLOATING
C1828 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n143 GND 0.05fF $ **FLOATING
C1829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n144 GND 0.02fF $ **FLOATING
C1830 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n145 GND 0.04fF $ **FLOATING
C1831 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n146 GND 0.06fF $ **FLOATING
C1832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n147 GND 0.02fF $ **FLOATING
C1833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n148 GND 0.04fF $ **FLOATING
C1834 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n149 GND 0.06fF $ **FLOATING
C1835 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n150 GND 0.02fF $ **FLOATING
C1836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n151 GND 0.05fF $ **FLOATING
C1837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n152 GND 0.06fF $ **FLOATING
C1838 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n153 GND 0.02fF $ **FLOATING
C1839 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n154 GND 0.05fF $ **FLOATING
C1840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n155 GND 0.06fF $ **FLOATING
C1841 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n156 GND 0.02fF $ **FLOATING
C1842 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n157 GND 0.05fF $ **FLOATING
C1843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n158 GND 0.06fF $ **FLOATING
C1844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t237 GND 0.02fF
C1845 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n159 GND 0.07fF $ **FLOATING
C1846 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n160 GND 0.02fF $ **FLOATING
C1847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n161 GND 0.03fF $ **FLOATING
C1848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n162 GND 0.06fF $ **FLOATING
C1849 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n163 GND 0.02fF $ **FLOATING
C1850 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n164 GND 0.04fF $ **FLOATING
C1851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n165 GND 0.06fF $ **FLOATING
C1852 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n166 GND 0.02fF $ **FLOATING
C1853 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n167 GND 0.05fF $ **FLOATING
C1854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n168 GND 0.06fF $ **FLOATING
C1855 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t8 GND 0.01fF
C1856 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t55 GND 0.01fF
C1857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n169 GND 0.04fF $ **FLOATING
C1858 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n170 GND 0.05fF $ **FLOATING
C1859 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n171 GND 0.02fF $ **FLOATING
C1860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n172 GND 0.03fF $ **FLOATING
C1861 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n173 GND 0.06fF $ **FLOATING
C1862 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n174 GND 0.02fF $ **FLOATING
C1863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n175 GND 0.05fF $ **FLOATING
C1864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n176 GND 0.06fF $ **FLOATING
C1865 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n177 GND 0.02fF $ **FLOATING
C1866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n178 GND 0.05fF $ **FLOATING
C1867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n179 GND 0.06fF $ **FLOATING
C1868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t229 GND 0.02fF
C1869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t15 GND 0.01fF
C1870 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n180 GND 0.10fF $ **FLOATING
C1871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n181 GND 0.04fF $ **FLOATING
C1872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n182 GND 0.02fF $ **FLOATING
C1873 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n183 GND 0.03fF $ **FLOATING
C1874 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n184 GND 0.06fF $ **FLOATING
C1875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n185 GND 0.02fF $ **FLOATING
C1876 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n186 GND 0.05fF $ **FLOATING
C1877 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n187 GND 0.06fF $ **FLOATING
C1878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n188 GND 0.02fF $ **FLOATING
C1879 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n189 GND 0.05fF $ **FLOATING
C1880 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n190 GND 0.06fF $ **FLOATING
C1881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n191 GND 0.02fF $ **FLOATING
C1882 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n192 GND 0.04fF $ **FLOATING
C1883 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n193 GND 0.06fF $ **FLOATING
C1884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t230 GND 0.02fF
C1885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n194 GND 0.06fF $ **FLOATING
C1886 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n195 GND 0.05fF $ **FLOATING
C1887 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t43 GND 0.01fF
C1888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n196 GND 0.03fF $ **FLOATING
C1889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n197 GND 0.05fF $ **FLOATING
C1890 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n198 GND 0.02fF $ **FLOATING
C1891 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n199 GND 0.04fF $ **FLOATING
C1892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n200 GND 0.06fF $ **FLOATING
C1893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n201 GND 0.02fF $ **FLOATING
C1894 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n202 GND 0.04fF $ **FLOATING
C1895 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n203 GND 0.06fF $ **FLOATING
C1896 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t160 GND 0.01fF
C1897 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t228 GND 0.02fF
C1898 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n204 GND 0.04fF $ **FLOATING
C1899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n205 GND 0.04fF $ **FLOATING
C1900 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n206 GND 0.02fF $ **FLOATING
C1901 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n207 GND 0.03fF $ **FLOATING
C1902 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n208 GND 0.06fF $ **FLOATING
C1903 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n209 GND 0.02fF $ **FLOATING
C1904 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n210 GND 0.05fF $ **FLOATING
C1905 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n211 GND 0.06fF $ **FLOATING
C1906 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n212 GND 0.02fF $ **FLOATING
C1907 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n213 GND 0.05fF $ **FLOATING
C1908 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n214 GND 0.06fF $ **FLOATING
C1909 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n215 GND 0.02fF $ **FLOATING
C1910 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n216 GND 0.05fF $ **FLOATING
C1911 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n217 GND 0.06fF $ **FLOATING
C1912 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t219 GND 0.04fF
C1913 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n218 GND 0.09fF $ **FLOATING
C1914 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n219 GND 0.02fF $ **FLOATING
C1915 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n220 GND 0.03fF $ **FLOATING
C1916 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n221 GND 0.06fF $ **FLOATING
C1917 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n222 GND 0.02fF $ **FLOATING
C1918 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n223 GND 0.04fF $ **FLOATING
C1919 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n224 GND 0.06fF $ **FLOATING
C1920 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t188 GND 0.01fF
C1921 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t110 GND 0.01fF
C1922 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n225 GND 0.04fF $ **FLOATING
C1923 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n226 GND 0.05fF $ **FLOATING
C1924 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n227 GND 0.02fF $ **FLOATING
C1925 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n228 GND 0.04fF $ **FLOATING
C1926 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n229 GND 0.06fF $ **FLOATING
C1927 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n230 GND 0.02fF $ **FLOATING
C1928 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n231 GND 0.04fF $ **FLOATING
C1929 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n232 GND 0.06fF $ **FLOATING
C1930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n233 GND 0.02fF $ **FLOATING
C1931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n234 GND 0.05fF $ **FLOATING
C1932 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n235 GND 0.06fF $ **FLOATING
C1933 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n236 GND 0.02fF $ **FLOATING
C1934 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n237 GND 0.05fF $ **FLOATING
C1935 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n238 GND 0.06fF $ **FLOATING
C1936 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n239 GND 0.02fF $ **FLOATING
C1937 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n240 GND 0.05fF $ **FLOATING
C1938 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n241 GND 0.06fF $ **FLOATING
C1939 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t54 GND 0.02fF
C1940 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n242 GND 0.07fF $ **FLOATING
C1941 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n243 GND 0.02fF $ **FLOATING
C1942 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n244 GND 0.03fF $ **FLOATING
C1943 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n245 GND 0.06fF $ **FLOATING
C1944 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n246 GND 0.02fF $ **FLOATING
C1945 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n247 GND 0.04fF $ **FLOATING
C1946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n248 GND 0.06fF $ **FLOATING
C1947 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n249 GND 0.02fF $ **FLOATING
C1948 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n250 GND 0.05fF $ **FLOATING
C1949 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n251 GND 0.06fF $ **FLOATING
C1950 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t94 GND 0.01fF
C1951 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t50 GND 0.01fF
C1952 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n252 GND 0.04fF $ **FLOATING
C1953 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n253 GND 0.05fF $ **FLOATING
C1954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n254 GND 0.02fF $ **FLOATING
C1955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n255 GND 0.03fF $ **FLOATING
C1956 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n256 GND 0.06fF $ **FLOATING
C1957 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n257 GND 0.02fF $ **FLOATING
C1958 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n258 GND 0.05fF $ **FLOATING
C1959 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n259 GND 0.06fF $ **FLOATING
C1960 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n260 GND 0.02fF $ **FLOATING
C1961 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n261 GND 0.05fF $ **FLOATING
C1962 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n262 GND 0.06fF $ **FLOATING
C1963 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t65 GND 0.02fF
C1964 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t71 GND 0.01fF
C1965 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n263 GND 0.10fF $ **FLOATING
C1966 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n264 GND 0.04fF $ **FLOATING
C1967 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n265 GND 0.02fF $ **FLOATING
C1968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n266 GND 0.03fF $ **FLOATING
C1969 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n267 GND 0.06fF $ **FLOATING
C1970 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n268 GND 0.02fF $ **FLOATING
C1971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n269 GND 0.05fF $ **FLOATING
C1972 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n270 GND 0.06fF $ **FLOATING
C1973 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n271 GND 0.02fF $ **FLOATING
C1974 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n272 GND 0.05fF $ **FLOATING
C1975 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n273 GND 0.06fF $ **FLOATING
C1976 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n274 GND 0.02fF $ **FLOATING
C1977 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n275 GND 0.04fF $ **FLOATING
C1978 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n276 GND 0.06fF $ **FLOATING
C1979 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t66 GND 0.02fF
C1980 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n277 GND 0.06fF $ **FLOATING
C1981 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n278 GND 0.05fF $ **FLOATING
C1982 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t150 GND 0.01fF
C1983 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n279 GND 0.03fF $ **FLOATING
C1984 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n280 GND 0.05fF $ **FLOATING
C1985 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n281 GND 0.02fF $ **FLOATING
C1986 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n282 GND 0.04fF $ **FLOATING
C1987 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n283 GND 0.06fF $ **FLOATING
C1988 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n284 GND 0.02fF $ **FLOATING
C1989 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n285 GND 0.04fF $ **FLOATING
C1990 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n286 GND 0.06fF $ **FLOATING
C1991 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t173 GND 0.01fF
C1992 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t64 GND 0.02fF
C1993 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n287 GND 0.04fF $ **FLOATING
C1994 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n288 GND 0.04fF $ **FLOATING
C1995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n289 GND 0.02fF $ **FLOATING
C1996 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n290 GND 0.03fF $ **FLOATING
C1997 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n291 GND 0.06fF $ **FLOATING
C1998 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n292 GND 0.02fF $ **FLOATING
C1999 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n293 GND 0.05fF $ **FLOATING
C2000 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n294 GND 0.06fF $ **FLOATING
C2001 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n295 GND 0.02fF $ **FLOATING
C2002 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n296 GND 0.05fF $ **FLOATING
C2003 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n297 GND 0.06fF $ **FLOATING
C2004 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n298 GND 0.02fF $ **FLOATING
C2005 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n299 GND 0.05fF $ **FLOATING
C2006 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n300 GND 0.06fF $ **FLOATING
C2007 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t111 GND 0.04fF
C2008 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n301 GND 0.09fF $ **FLOATING
C2009 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n302 GND 0.02fF $ **FLOATING
C2010 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n303 GND 0.03fF $ **FLOATING
C2011 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n304 GND 0.06fF $ **FLOATING
C2012 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n305 GND 0.02fF $ **FLOATING
C2013 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n306 GND 0.04fF $ **FLOATING
C2014 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n307 GND 0.06fF $ **FLOATING
C2015 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t185 GND 0.01fF
C2016 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t82 GND 0.01fF
C2017 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n308 GND 0.04fF $ **FLOATING
C2018 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n309 GND 0.05fF $ **FLOATING
C2019 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n310 GND 0.02fF $ **FLOATING
C2020 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n311 GND 0.04fF $ **FLOATING
C2021 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n312 GND 0.06fF $ **FLOATING
C2022 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n313 GND 0.02fF $ **FLOATING
C2023 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n314 GND 0.04fF $ **FLOATING
C2024 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n315 GND 0.06fF $ **FLOATING
C2025 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n316 GND 0.02fF $ **FLOATING
C2026 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n317 GND 0.05fF $ **FLOATING
C2027 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n318 GND 0.06fF $ **FLOATING
C2028 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n319 GND 0.02fF $ **FLOATING
C2029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n320 GND 0.05fF $ **FLOATING
C2030 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n321 GND 0.06fF $ **FLOATING
C2031 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n322 GND 0.02fF $ **FLOATING
C2032 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n323 GND 0.05fF $ **FLOATING
C2033 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n324 GND 0.06fF $ **FLOATING
C2034 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t49 GND 0.02fF
C2035 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n325 GND 0.07fF $ **FLOATING
C2036 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n326 GND 0.02fF $ **FLOATING
C2037 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n327 GND 0.03fF $ **FLOATING
C2038 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n328 GND 0.06fF $ **FLOATING
C2039 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n329 GND 0.02fF $ **FLOATING
C2040 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n330 GND 0.04fF $ **FLOATING
C2041 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n331 GND 0.06fF $ **FLOATING
C2042 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n332 GND 0.02fF $ **FLOATING
C2043 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n333 GND 0.05fF $ **FLOATING
C2044 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n334 GND 0.06fF $ **FLOATING
C2045 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t89 GND 0.01fF
C2046 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t91 GND 0.01fF
C2047 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n335 GND 0.04fF $ **FLOATING
C2048 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n336 GND 0.05fF $ **FLOATING
C2049 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n337 GND 0.02fF $ **FLOATING
C2050 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n338 GND 0.03fF $ **FLOATING
C2051 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n339 GND 0.06fF $ **FLOATING
C2052 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n340 GND 0.02fF $ **FLOATING
C2053 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n341 GND 0.05fF $ **FLOATING
C2054 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n342 GND 0.06fF $ **FLOATING
C2055 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n343 GND 0.02fF $ **FLOATING
C2056 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n344 GND 0.05fF $ **FLOATING
C2057 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n345 GND 0.06fF $ **FLOATING
C2058 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t200 GND 0.02fF
C2059 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t113 GND 0.01fF
C2060 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n346 GND 0.10fF $ **FLOATING
C2061 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n347 GND 0.04fF $ **FLOATING
C2062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n348 GND 0.02fF $ **FLOATING
C2063 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n349 GND 0.03fF $ **FLOATING
C2064 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n350 GND 0.06fF $ **FLOATING
C2065 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n351 GND 0.02fF $ **FLOATING
C2066 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n352 GND 0.05fF $ **FLOATING
C2067 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n353 GND 0.06fF $ **FLOATING
C2068 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n354 GND 0.02fF $ **FLOATING
C2069 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n355 GND 0.05fF $ **FLOATING
C2070 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n356 GND 0.06fF $ **FLOATING
C2071 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n357 GND 0.02fF $ **FLOATING
C2072 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n358 GND 0.04fF $ **FLOATING
C2073 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n359 GND 0.06fF $ **FLOATING
C2074 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t198 GND 0.02fF
C2075 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n360 GND 0.06fF $ **FLOATING
C2076 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n361 GND 0.05fF $ **FLOATING
C2077 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t112 GND 0.01fF
C2078 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n362 GND 0.03fF $ **FLOATING
C2079 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n363 GND 0.05fF $ **FLOATING
C2080 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n364 GND 0.02fF $ **FLOATING
C2081 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n365 GND 0.04fF $ **FLOATING
C2082 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n366 GND 0.06fF $ **FLOATING
C2083 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n367 GND 0.02fF $ **FLOATING
C2084 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n368 GND 0.04fF $ **FLOATING
C2085 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n369 GND 0.06fF $ **FLOATING
C2086 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t175 GND 0.01fF
C2087 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t199 GND 0.02fF
C2088 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n370 GND 0.04fF $ **FLOATING
C2089 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n371 GND 0.04fF $ **FLOATING
C2090 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n372 GND 0.02fF $ **FLOATING
C2091 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n373 GND 0.03fF $ **FLOATING
C2092 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n374 GND 0.06fF $ **FLOATING
C2093 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n375 GND 0.02fF $ **FLOATING
C2094 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n376 GND 0.05fF $ **FLOATING
C2095 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n377 GND 0.06fF $ **FLOATING
C2096 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n378 GND 0.02fF $ **FLOATING
C2097 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n379 GND 0.05fF $ **FLOATING
C2098 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n380 GND 0.06fF $ **FLOATING
C2099 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n381 GND 0.02fF $ **FLOATING
C2100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n382 GND 0.05fF $ **FLOATING
C2101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n383 GND 0.06fF $ **FLOATING
C2102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t16 GND 0.04fF
C2103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n384 GND 0.09fF $ **FLOATING
C2104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n385 GND 0.02fF $ **FLOATING
C2105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n386 GND 0.03fF $ **FLOATING
C2106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n387 GND 0.06fF $ **FLOATING
C2107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n388 GND 0.02fF $ **FLOATING
C2108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n389 GND 0.04fF $ **FLOATING
C2109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n390 GND 0.06fF $ **FLOATING
C2110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t193 GND 0.01fF
C2111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t72 GND 0.01fF
C2112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n391 GND 0.04fF $ **FLOATING
C2113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n392 GND 0.05fF $ **FLOATING
C2114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n393 GND 0.02fF $ **FLOATING
C2115 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n394 GND 0.04fF $ **FLOATING
C2116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n395 GND 0.06fF $ **FLOATING
C2117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n396 GND 0.02fF $ **FLOATING
C2118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n397 GND 0.04fF $ **FLOATING
C2119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n398 GND 0.06fF $ **FLOATING
C2120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n399 GND 0.02fF $ **FLOATING
C2121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n400 GND 0.05fF $ **FLOATING
C2122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n401 GND 0.06fF $ **FLOATING
C2123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n402 GND 0.02fF $ **FLOATING
C2124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n403 GND 0.05fF $ **FLOATING
C2125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n404 GND 0.06fF $ **FLOATING
C2126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n405 GND 0.02fF $ **FLOATING
C2127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n406 GND 0.05fF $ **FLOATING
C2128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n407 GND 0.06fF $ **FLOATING
C2129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t92 GND 0.02fF
C2130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n408 GND 0.07fF $ **FLOATING
C2131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n409 GND 0.02fF $ **FLOATING
C2132 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n410 GND 0.03fF $ **FLOATING
C2133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n411 GND 0.06fF $ **FLOATING
C2134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n412 GND 0.02fF $ **FLOATING
C2135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n413 GND 0.04fF $ **FLOATING
C2136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n414 GND 0.06fF $ **FLOATING
C2137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n415 GND 0.02fF $ **FLOATING
C2138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n416 GND 0.05fF $ **FLOATING
C2139 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n417 GND 0.06fF $ **FLOATING
C2140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t48 GND 0.01fF
C2141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t75 GND 0.01fF
C2142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n418 GND 0.04fF $ **FLOATING
C2143 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n419 GND 0.05fF $ **FLOATING
C2144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n420 GND 0.02fF $ **FLOATING
C2145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n421 GND 0.03fF $ **FLOATING
C2146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n422 GND 0.06fF $ **FLOATING
C2147 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n423 GND 0.02fF $ **FLOATING
C2148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n424 GND 0.05fF $ **FLOATING
C2149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n425 GND 0.06fF $ **FLOATING
C2150 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n426 GND 0.02fF $ **FLOATING
C2151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n427 GND 0.05fF $ **FLOATING
C2152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n428 GND 0.06fF $ **FLOATING
C2153 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t11 GND 0.02fF
C2154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t57 GND 0.01fF
C2155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n429 GND 0.10fF $ **FLOATING
C2156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n430 GND 0.04fF $ **FLOATING
C2157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n431 GND 0.02fF $ **FLOATING
C2158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n432 GND 0.03fF $ **FLOATING
C2159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n433 GND 0.06fF $ **FLOATING
C2160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n434 GND 0.02fF $ **FLOATING
C2161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n435 GND 0.05fF $ **FLOATING
C2162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n436 GND 0.06fF $ **FLOATING
C2163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n437 GND 0.02fF $ **FLOATING
C2164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n438 GND 0.05fF $ **FLOATING
C2165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n439 GND 0.06fF $ **FLOATING
C2166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n440 GND 0.02fF $ **FLOATING
C2167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n441 GND 0.04fF $ **FLOATING
C2168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n442 GND 0.06fF $ **FLOATING
C2169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t12 GND 0.02fF
C2170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n443 GND 0.06fF $ **FLOATING
C2171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n444 GND 0.05fF $ **FLOATING
C2172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t99 GND 0.01fF
C2173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n445 GND 0.03fF $ **FLOATING
C2174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n446 GND 0.05fF $ **FLOATING
C2175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n447 GND 0.02fF $ **FLOATING
C2176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n448 GND 0.04fF $ **FLOATING
C2177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n449 GND 0.06fF $ **FLOATING
C2178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n450 GND 0.02fF $ **FLOATING
C2179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n451 GND 0.04fF $ **FLOATING
C2180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n452 GND 0.06fF $ **FLOATING
C2181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t174 GND 0.01fF
C2182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t10 GND 0.02fF
C2183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n453 GND 0.04fF $ **FLOATING
C2184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n454 GND 0.04fF $ **FLOATING
C2185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n455 GND 0.02fF $ **FLOATING
C2186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n456 GND 0.03fF $ **FLOATING
C2187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n457 GND 0.06fF $ **FLOATING
C2188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n458 GND 0.02fF $ **FLOATING
C2189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n459 GND 0.05fF $ **FLOATING
C2190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n460 GND 0.06fF $ **FLOATING
C2191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n461 GND 0.02fF $ **FLOATING
C2192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n462 GND 0.05fF $ **FLOATING
C2193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n463 GND 0.06fF $ **FLOATING
C2194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n464 GND 0.02fF $ **FLOATING
C2195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n465 GND 0.05fF $ **FLOATING
C2196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n466 GND 0.06fF $ **FLOATING
C2197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t223 GND 0.04fF
C2198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n467 GND 0.09fF $ **FLOATING
C2199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n468 GND 0.02fF $ **FLOATING
C2200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n469 GND 0.03fF $ **FLOATING
C2201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n470 GND 0.06fF $ **FLOATING
C2202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n471 GND 0.02fF $ **FLOATING
C2203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n472 GND 0.04fF $ **FLOATING
C2204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n473 GND 0.06fF $ **FLOATING
C2205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t195 GND 0.01fF
C2206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t216 GND 0.01fF
C2207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n474 GND 0.04fF $ **FLOATING
C2208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n475 GND 0.05fF $ **FLOATING
C2209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n476 GND 0.02fF $ **FLOATING
C2210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n477 GND 0.04fF $ **FLOATING
C2211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n478 GND 0.06fF $ **FLOATING
C2212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n479 GND 0.02fF $ **FLOATING
C2213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n480 GND 0.04fF $ **FLOATING
C2214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n481 GND 0.06fF $ **FLOATING
C2215 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n482 GND 0.02fF $ **FLOATING
C2216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n483 GND 0.05fF $ **FLOATING
C2217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n484 GND 0.06fF $ **FLOATING
C2218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n485 GND 0.02fF $ **FLOATING
C2219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n486 GND 0.05fF $ **FLOATING
C2220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n487 GND 0.06fF $ **FLOATING
C2221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n488 GND 0.02fF $ **FLOATING
C2222 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n489 GND 0.05fF $ **FLOATING
C2223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n490 GND 0.06fF $ **FLOATING
C2224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t76 GND 0.02fF
C2225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n491 GND 0.07fF $ **FLOATING
C2226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n492 GND 0.02fF $ **FLOATING
C2227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n493 GND 0.03fF $ **FLOATING
C2228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n494 GND 0.06fF $ **FLOATING
C2229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n495 GND 0.02fF $ **FLOATING
C2230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n496 GND 0.04fF $ **FLOATING
C2231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n497 GND 0.06fF $ **FLOATING
C2232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n498 GND 0.02fF $ **FLOATING
C2233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n499 GND 0.05fF $ **FLOATING
C2234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n500 GND 0.06fF $ **FLOATING
C2235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t232 GND 0.01fF
C2236 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t101 GND 0.01fF
C2237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n501 GND 0.04fF $ **FLOATING
C2238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n502 GND 0.05fF $ **FLOATING
C2239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n503 GND 0.02fF $ **FLOATING
C2240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n504 GND 0.03fF $ **FLOATING
C2241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n505 GND 0.06fF $ **FLOATING
C2242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n506 GND 0.02fF $ **FLOATING
C2243 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n507 GND 0.05fF $ **FLOATING
C2244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n508 GND 0.06fF $ **FLOATING
C2245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n509 GND 0.02fF $ **FLOATING
C2246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n510 GND 0.05fF $ **FLOATING
C2247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n511 GND 0.06fF $ **FLOATING
C2248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t67 GND 0.02fF
C2249 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t155 GND 0.01fF
C2250 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n512 GND 0.10fF $ **FLOATING
C2251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n513 GND 0.04fF $ **FLOATING
C2252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n514 GND 0.02fF $ **FLOATING
C2253 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n515 GND 0.03fF $ **FLOATING
C2254 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n516 GND 0.06fF $ **FLOATING
C2255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n517 GND 0.02fF $ **FLOATING
C2256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n518 GND 0.05fF $ **FLOATING
C2257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n519 GND 0.06fF $ **FLOATING
C2258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n520 GND 0.02fF $ **FLOATING
C2259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n521 GND 0.05fF $ **FLOATING
C2260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n522 GND 0.06fF $ **FLOATING
C2261 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n523 GND 0.02fF $ **FLOATING
C2262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n524 GND 0.04fF $ **FLOATING
C2263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n525 GND 0.06fF $ **FLOATING
C2264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t68 GND 0.02fF
C2265 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n526 GND 0.06fF $ **FLOATING
C2266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n527 GND 0.05fF $ **FLOATING
C2267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t7 GND 0.01fF
C2268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n528 GND 0.03fF $ **FLOATING
C2269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n529 GND 0.05fF $ **FLOATING
C2270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n530 GND 0.02fF $ **FLOATING
C2271 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n531 GND 0.04fF $ **FLOATING
C2272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n532 GND 0.06fF $ **FLOATING
C2273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n533 GND 0.02fF $ **FLOATING
C2274 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n534 GND 0.04fF $ **FLOATING
C2275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n535 GND 0.06fF $ **FLOATING
C2276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t179 GND 0.01fF
C2277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t69 GND 0.02fF
C2278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n536 GND 0.04fF $ **FLOATING
C2279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n537 GND 0.04fF $ **FLOATING
C2280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n538 GND 0.02fF $ **FLOATING
C2281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n539 GND 0.03fF $ **FLOATING
C2282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n540 GND 0.06fF $ **FLOATING
C2283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n541 GND 0.02fF $ **FLOATING
C2284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n542 GND 0.05fF $ **FLOATING
C2285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n543 GND 0.06fF $ **FLOATING
C2286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n544 GND 0.02fF $ **FLOATING
C2287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n545 GND 0.05fF $ **FLOATING
C2288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n546 GND 0.06fF $ **FLOATING
C2289 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n547 GND 0.02fF $ **FLOATING
C2290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n548 GND 0.05fF $ **FLOATING
C2291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n549 GND 0.06fF $ **FLOATING
C2292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t42 GND 0.04fF
C2293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n550 GND 0.09fF $ **FLOATING
C2294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n551 GND 0.02fF $ **FLOATING
C2295 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n552 GND 0.03fF $ **FLOATING
C2296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n553 GND 0.06fF $ **FLOATING
C2297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n554 GND 0.02fF $ **FLOATING
C2298 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n555 GND 0.04fF $ **FLOATING
C2299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n556 GND 0.06fF $ **FLOATING
C2300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t168 GND 0.01fF
C2301 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t204 GND 0.01fF
C2302 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n557 GND 0.04fF $ **FLOATING
C2303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n558 GND 0.05fF $ **FLOATING
C2304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n559 GND 0.02fF $ **FLOATING
C2305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n560 GND 0.04fF $ **FLOATING
C2306 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n561 GND 0.06fF $ **FLOATING
C2307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n562 GND 0.02fF $ **FLOATING
C2308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n563 GND 0.04fF $ **FLOATING
C2309 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n564 GND 0.06fF $ **FLOATING
C2310 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n565 GND 0.02fF $ **FLOATING
C2311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n566 GND 0.05fF $ **FLOATING
C2312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n567 GND 0.06fF $ **FLOATING
C2313 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n568 GND 0.02fF $ **FLOATING
C2314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n569 GND 0.05fF $ **FLOATING
C2315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n570 GND 0.06fF $ **FLOATING
C2316 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n571 GND 0.02fF $ **FLOATING
C2317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n572 GND 0.05fF $ **FLOATING
C2318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n573 GND 0.06fF $ **FLOATING
C2319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t100 GND 0.02fF
C2320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n574 GND 0.07fF $ **FLOATING
C2321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n575 GND 0.02fF $ **FLOATING
C2322 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n576 GND 0.03fF $ **FLOATING
C2323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n577 GND 0.06fF $ **FLOATING
C2324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n578 GND 0.02fF $ **FLOATING
C2325 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n579 GND 0.04fF $ **FLOATING
C2326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n580 GND 0.06fF $ **FLOATING
C2327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n581 GND 0.02fF $ **FLOATING
C2328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n582 GND 0.05fF $ **FLOATING
C2329 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n583 GND 0.06fF $ **FLOATING
C2330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t136 GND 0.01fF
C2331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t51 GND 0.01fF
C2332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n584 GND 0.04fF $ **FLOATING
C2333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n585 GND 0.05fF $ **FLOATING
C2334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n586 GND 0.02fF $ **FLOATING
C2335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n587 GND 0.03fF $ **FLOATING
C2336 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n588 GND 0.06fF $ **FLOATING
C2337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n589 GND 0.02fF $ **FLOATING
C2338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n590 GND 0.05fF $ **FLOATING
C2339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n591 GND 0.06fF $ **FLOATING
C2340 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n592 GND 0.02fF $ **FLOATING
C2341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n593 GND 0.05fF $ **FLOATING
C2342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n594 GND 0.06fF $ **FLOATING
C2343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t26 GND 0.02fF
C2344 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t218 GND 0.01fF
C2345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n595 GND 0.10fF $ **FLOATING
C2346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n596 GND 0.04fF $ **FLOATING
C2347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n597 GND 0.02fF $ **FLOATING
C2348 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n598 GND 0.03fF $ **FLOATING
C2349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n599 GND 0.06fF $ **FLOATING
C2350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n600 GND 0.02fF $ **FLOATING
C2351 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n601 GND 0.05fF $ **FLOATING
C2352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n602 GND 0.06fF $ **FLOATING
C2353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n603 GND 0.02fF $ **FLOATING
C2354 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n604 GND 0.05fF $ **FLOATING
C2355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n605 GND 0.06fF $ **FLOATING
C2356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n606 GND 0.02fF $ **FLOATING
C2357 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n607 GND 0.04fF $ **FLOATING
C2358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n608 GND 0.06fF $ **FLOATING
C2359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t27 GND 0.02fF
C2360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n609 GND 0.06fF $ **FLOATING
C2361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n610 GND 0.05fF $ **FLOATING
C2362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t98 GND 0.01fF
C2363 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n611 GND 0.03fF $ **FLOATING
C2364 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n612 GND 0.05fF $ **FLOATING
C2365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n613 GND 0.02fF $ **FLOATING
C2366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n614 GND 0.04fF $ **FLOATING
C2367 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n615 GND 0.06fF $ **FLOATING
C2368 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n616 GND 0.02fF $ **FLOATING
C2369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n617 GND 0.04fF $ **FLOATING
C2370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n618 GND 0.06fF $ **FLOATING
C2371 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t178 GND 0.01fF
C2372 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t28 GND 0.02fF
C2373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n619 GND 0.04fF $ **FLOATING
C2374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n620 GND 0.04fF $ **FLOATING
C2375 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n621 GND 0.02fF $ **FLOATING
C2376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n622 GND 0.03fF $ **FLOATING
C2377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n623 GND 0.06fF $ **FLOATING
C2378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n624 GND 0.02fF $ **FLOATING
C2379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n625 GND 0.05fF $ **FLOATING
C2380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n626 GND 0.06fF $ **FLOATING
C2381 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n627 GND 0.02fF $ **FLOATING
C2382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n628 GND 0.05fF $ **FLOATING
C2383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n629 GND 0.06fF $ **FLOATING
C2384 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n630 GND 0.02fF $ **FLOATING
C2385 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n631 GND 0.05fF $ **FLOATING
C2386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n632 GND 0.06fF $ **FLOATING
C2387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t105 GND 0.04fF
C2388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n633 GND 0.09fF $ **FLOATING
C2389 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n634 GND 0.02fF $ **FLOATING
C2390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n635 GND 0.03fF $ **FLOATING
C2391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n636 GND 0.06fF $ **FLOATING
C2392 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n637 GND 0.02fF $ **FLOATING
C2393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n638 GND 0.04fF $ **FLOATING
C2394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n639 GND 0.06fF $ **FLOATING
C2395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t171 GND 0.01fF
C2396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t70 GND 0.01fF
C2397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n640 GND 0.04fF $ **FLOATING
C2398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n641 GND 0.05fF $ **FLOATING
C2399 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n642 GND 0.02fF $ **FLOATING
C2400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n643 GND 0.04fF $ **FLOATING
C2401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n644 GND 0.06fF $ **FLOATING
C2402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n645 GND 0.02fF $ **FLOATING
C2403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n646 GND 0.04fF $ **FLOATING
C2404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n647 GND 0.06fF $ **FLOATING
C2405 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n648 GND 0.02fF $ **FLOATING
C2406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n649 GND 0.05fF $ **FLOATING
C2407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n650 GND 0.06fF $ **FLOATING
C2408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n651 GND 0.02fF $ **FLOATING
C2409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n652 GND 0.05fF $ **FLOATING
C2410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n653 GND 0.06fF $ **FLOATING
C2411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n654 GND 0.02fF $ **FLOATING
C2412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n655 GND 0.05fF $ **FLOATING
C2413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n656 GND 0.06fF $ **FLOATING
C2414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t52 GND 0.02fF
C2415 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n657 GND 0.07fF $ **FLOATING
C2416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n658 GND 0.02fF $ **FLOATING
C2417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n659 GND 0.03fF $ **FLOATING
C2418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n660 GND 0.06fF $ **FLOATING
C2419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n661 GND 0.02fF $ **FLOATING
C2420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n662 GND 0.04fF $ **FLOATING
C2421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n663 GND 0.06fF $ **FLOATING
C2422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n664 GND 0.02fF $ **FLOATING
C2423 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n665 GND 0.05fF $ **FLOATING
C2424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n666 GND 0.06fF $ **FLOATING
C2425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t97 GND 0.01fF
C2426 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t106 GND 0.01fF
C2427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n667 GND 0.04fF $ **FLOATING
C2428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n668 GND 0.05fF $ **FLOATING
C2429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n669 GND 0.02fF $ **FLOATING
C2430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n670 GND 0.03fF $ **FLOATING
C2431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n671 GND 0.06fF $ **FLOATING
C2432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n672 GND 0.02fF $ **FLOATING
C2433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n673 GND 0.05fF $ **FLOATING
C2434 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n674 GND 0.06fF $ **FLOATING
C2435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n675 GND 0.02fF $ **FLOATING
C2436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n676 GND 0.05fF $ **FLOATING
C2437 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n677 GND 0.06fF $ **FLOATING
C2438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t80 GND 0.02fF
C2439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t206 GND 0.01fF
C2440 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n678 GND 0.10fF $ **FLOATING
C2441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n679 GND 0.04fF $ **FLOATING
C2442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n680 GND 0.02fF $ **FLOATING
C2443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n681 GND 0.03fF $ **FLOATING
C2444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n682 GND 0.06fF $ **FLOATING
C2445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n683 GND 0.02fF $ **FLOATING
C2446 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n684 GND 0.05fF $ **FLOATING
C2447 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n685 GND 0.06fF $ **FLOATING
C2448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n686 GND 0.02fF $ **FLOATING
C2449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n687 GND 0.05fF $ **FLOATING
C2450 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n688 GND 0.06fF $ **FLOATING
C2451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n689 GND 0.02fF $ **FLOATING
C2452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n690 GND 0.04fF $ **FLOATING
C2453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n691 GND 0.06fF $ **FLOATING
C2454 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t79 GND 0.02fF
C2455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n692 GND 0.06fF $ **FLOATING
C2456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n693 GND 0.05fF $ **FLOATING
C2457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t224 GND 0.01fF
C2458 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n694 GND 0.03fF $ **FLOATING
C2459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n695 GND 0.05fF $ **FLOATING
C2460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n696 GND 0.02fF $ **FLOATING
C2461 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n697 GND 0.04fF $ **FLOATING
C2462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n698 GND 0.06fF $ **FLOATING
C2463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n699 GND 0.02fF $ **FLOATING
C2464 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n700 GND 0.04fF $ **FLOATING
C2465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n701 GND 0.06fF $ **FLOATING
C2466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t177 GND 0.01fF
C2467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t81 GND 0.02fF
C2468 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n702 GND 0.04fF $ **FLOATING
C2469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n703 GND 0.04fF $ **FLOATING
C2470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n704 GND 0.02fF $ **FLOATING
C2471 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n705 GND 0.03fF $ **FLOATING
C2472 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n706 GND 0.06fF $ **FLOATING
C2473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n707 GND 0.02fF $ **FLOATING
C2474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n708 GND 0.05fF $ **FLOATING
C2475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n709 GND 0.06fF $ **FLOATING
C2476 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n710 GND 0.02fF $ **FLOATING
C2477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n711 GND 0.05fF $ **FLOATING
C2478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n712 GND 0.06fF $ **FLOATING
C2479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n713 GND 0.02fF $ **FLOATING
C2480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n714 GND 0.05fF $ **FLOATING
C2481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n715 GND 0.06fF $ **FLOATING
C2482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t87 GND 0.04fF
C2483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n716 GND 0.09fF $ **FLOATING
C2484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n717 GND 0.02fF $ **FLOATING
C2485 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n718 GND 0.03fF $ **FLOATING
C2486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n719 GND 0.06fF $ **FLOATING
C2487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n720 GND 0.02fF $ **FLOATING
C2488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n721 GND 0.04fF $ **FLOATING
C2489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n722 GND 0.06fF $ **FLOATING
C2490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t170 GND 0.01fF
C2491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t127 GND 0.01fF
C2492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n723 GND 0.04fF $ **FLOATING
C2493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n724 GND 0.05fF $ **FLOATING
C2494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n725 GND 0.02fF $ **FLOATING
C2495 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n726 GND 0.04fF $ **FLOATING
C2496 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n727 GND 0.06fF $ **FLOATING
C2497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n728 GND 0.02fF $ **FLOATING
C2498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n729 GND 0.04fF $ **FLOATING
C2499 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n730 GND 0.06fF $ **FLOATING
C2500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n731 GND 0.02fF $ **FLOATING
C2501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n732 GND 0.05fF $ **FLOATING
C2502 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n733 GND 0.06fF $ **FLOATING
C2503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n734 GND 0.02fF $ **FLOATING
C2504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n735 GND 0.05fF $ **FLOATING
C2505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n736 GND 0.06fF $ **FLOATING
C2506 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n737 GND 0.02fF $ **FLOATING
C2507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n738 GND 0.05fF $ **FLOATING
C2508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n739 GND 0.06fF $ **FLOATING
C2509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t107 GND 0.02fF
C2510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n740 GND 0.07fF $ **FLOATING
C2511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n741 GND 0.02fF $ **FLOATING
C2512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n742 GND 0.03fF $ **FLOATING
C2513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n743 GND 0.06fF $ **FLOATING
C2514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n744 GND 0.02fF $ **FLOATING
C2515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n745 GND 0.04fF $ **FLOATING
C2516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n746 GND 0.06fF $ **FLOATING
C2517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n747 GND 0.02fF $ **FLOATING
C2518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n748 GND 0.05fF $ **FLOATING
C2519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n749 GND 0.06fF $ **FLOATING
C2520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t145 GND 0.01fF
C2521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t36 GND 0.01fF
C2522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n750 GND 0.04fF $ **FLOATING
C2523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n751 GND 0.05fF $ **FLOATING
C2524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n752 GND 0.02fF $ **FLOATING
C2525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n753 GND 0.03fF $ **FLOATING
C2526 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n754 GND 0.06fF $ **FLOATING
C2527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n755 GND 0.02fF $ **FLOATING
C2528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n756 GND 0.05fF $ **FLOATING
C2529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n757 GND 0.06fF $ **FLOATING
C2530 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n758 GND 0.02fF $ **FLOATING
C2531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n759 GND 0.05fF $ **FLOATING
C2532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n760 GND 0.06fF $ **FLOATING
C2533 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t143 GND 0.02fF
C2534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t120 GND 0.01fF
C2535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n761 GND 0.10fF $ **FLOATING
C2536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n762 GND 0.04fF $ **FLOATING
C2537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n763 GND 0.02fF $ **FLOATING
C2538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n764 GND 0.03fF $ **FLOATING
C2539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n765 GND 0.06fF $ **FLOATING
C2540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n766 GND 0.02fF $ **FLOATING
C2541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n767 GND 0.05fF $ **FLOATING
C2542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n768 GND 0.06fF $ **FLOATING
C2543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n769 GND 0.02fF $ **FLOATING
C2544 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n770 GND 0.05fF $ **FLOATING
C2545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n771 GND 0.06fF $ **FLOATING
C2546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n772 GND 0.02fF $ **FLOATING
C2547 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n773 GND 0.04fF $ **FLOATING
C2548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n774 GND 0.06fF $ **FLOATING
C2549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t142 GND 0.02fF
C2550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n775 GND 0.06fF $ **FLOATING
C2551 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n776 GND 0.05fF $ **FLOATING
C2552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t93 GND 0.01fF
C2553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n777 GND 0.03fF $ **FLOATING
C2554 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n778 GND 0.05fF $ **FLOATING
C2555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n779 GND 0.02fF $ **FLOATING
C2556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n780 GND 0.04fF $ **FLOATING
C2557 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n781 GND 0.06fF $ **FLOATING
C2558 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n782 GND 0.02fF $ **FLOATING
C2559 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n783 GND 0.04fF $ **FLOATING
C2560 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n784 GND 0.06fF $ **FLOATING
C2561 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t192 GND 0.01fF
C2562 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t141 GND 0.02fF
C2563 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n785 GND 0.04fF $ **FLOATING
C2564 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n786 GND 0.04fF $ **FLOATING
C2565 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n787 GND 0.02fF $ **FLOATING
C2566 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n788 GND 0.03fF $ **FLOATING
C2567 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n789 GND 0.06fF $ **FLOATING
C2568 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n790 GND 0.02fF $ **FLOATING
C2569 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n791 GND 0.05fF $ **FLOATING
C2570 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n792 GND 0.06fF $ **FLOATING
C2571 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n793 GND 0.02fF $ **FLOATING
C2572 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n794 GND 0.05fF $ **FLOATING
C2573 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n795 GND 0.06fF $ **FLOATING
C2574 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n796 GND 0.02fF $ **FLOATING
C2575 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n797 GND 0.05fF $ **FLOATING
C2576 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n798 GND 0.06fF $ **FLOATING
C2577 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t212 GND 0.04fF
C2578 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n799 GND 0.09fF $ **FLOATING
C2579 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n800 GND 0.02fF $ **FLOATING
C2580 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n801 GND 0.03fF $ **FLOATING
C2581 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n802 GND 0.06fF $ **FLOATING
C2582 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n803 GND 0.02fF $ **FLOATING
C2583 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n804 GND 0.04fF $ **FLOATING
C2584 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n805 GND 0.06fF $ **FLOATING
C2585 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t169 GND 0.01fF
C2586 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t74 GND 0.01fF
C2587 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n806 GND 0.04fF $ **FLOATING
C2588 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n807 GND 0.05fF $ **FLOATING
C2589 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n808 GND 0.02fF $ **FLOATING
C2590 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n809 GND 0.04fF $ **FLOATING
C2591 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n810 GND 0.06fF $ **FLOATING
C2592 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n811 GND 0.02fF $ **FLOATING
C2593 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n812 GND 0.04fF $ **FLOATING
C2594 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n813 GND 0.06fF $ **FLOATING
C2595 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n814 GND 0.02fF $ **FLOATING
C2596 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n815 GND 0.05fF $ **FLOATING
C2597 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n816 GND 0.06fF $ **FLOATING
C2598 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n817 GND 0.02fF $ **FLOATING
C2599 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n818 GND 0.05fF $ **FLOATING
C2600 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n819 GND 0.06fF $ **FLOATING
C2601 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n820 GND 0.02fF $ **FLOATING
C2602 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n821 GND 0.05fF $ **FLOATING
C2603 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n822 GND 0.06fF $ **FLOATING
C2604 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t35 GND 0.02fF
C2605 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n823 GND 0.07fF $ **FLOATING
C2606 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n824 GND 0.02fF $ **FLOATING
C2607 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n825 GND 0.03fF $ **FLOATING
C2608 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n826 GND 0.06fF $ **FLOATING
C2609 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n827 GND 0.02fF $ **FLOATING
C2610 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n828 GND 0.04fF $ **FLOATING
C2611 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n829 GND 0.06fF $ **FLOATING
C2612 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n830 GND 0.02fF $ **FLOATING
C2613 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n831 GND 0.05fF $ **FLOATING
C2614 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n832 GND 0.06fF $ **FLOATING
C2615 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t73 GND 0.01fF
C2616 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t18 GND 0.01fF
C2617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n833 GND 0.04fF $ **FLOATING
C2618 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n834 GND 0.05fF $ **FLOATING
C2619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n835 GND 0.02fF $ **FLOATING
C2620 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n836 GND 0.03fF $ **FLOATING
C2621 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n837 GND 0.06fF $ **FLOATING
C2622 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n838 GND 0.02fF $ **FLOATING
C2623 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n839 GND 0.05fF $ **FLOATING
C2624 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n840 GND 0.06fF $ **FLOATING
C2625 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n841 GND 0.02fF $ **FLOATING
C2626 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n842 GND 0.05fF $ **FLOATING
C2627 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n843 GND 0.06fF $ **FLOATING
C2628 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t102 GND 0.02fF
C2629 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t17 GND 0.01fF
C2630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n844 GND 0.10fF $ **FLOATING
C2631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n845 GND 0.04fF $ **FLOATING
C2632 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n846 GND 0.02fF $ **FLOATING
C2633 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n847 GND 0.03fF $ **FLOATING
C2634 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n848 GND 0.06fF $ **FLOATING
C2635 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n849 GND 0.02fF $ **FLOATING
C2636 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n850 GND 0.05fF $ **FLOATING
C2637 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n851 GND 0.06fF $ **FLOATING
C2638 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n852 GND 0.02fF $ **FLOATING
C2639 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n853 GND 0.05fF $ **FLOATING
C2640 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n854 GND 0.06fF $ **FLOATING
C2641 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n855 GND 0.02fF $ **FLOATING
C2642 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n856 GND 0.04fF $ **FLOATING
C2643 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n857 GND 0.06fF $ **FLOATING
C2644 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t103 GND 0.02fF
C2645 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n858 GND 0.06fF $ **FLOATING
C2646 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n859 GND 0.05fF $ **FLOATING
C2647 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t151 GND 0.01fF
C2648 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n860 GND 0.03fF $ **FLOATING
C2649 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n861 GND 0.05fF $ **FLOATING
C2650 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n862 GND 0.02fF $ **FLOATING
C2651 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n863 GND 0.04fF $ **FLOATING
C2652 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n864 GND 0.06fF $ **FLOATING
C2653 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n865 GND 0.02fF $ **FLOATING
C2654 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n866 GND 0.04fF $ **FLOATING
C2655 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n867 GND 0.06fF $ **FLOATING
C2656 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t190 GND 0.01fF
C2657 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t104 GND 0.02fF
C2658 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n868 GND 0.04fF $ **FLOATING
C2659 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n869 GND 0.04fF $ **FLOATING
C2660 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n870 GND 0.02fF $ **FLOATING
C2661 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n871 GND 0.03fF $ **FLOATING
C2662 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n872 GND 0.06fF $ **FLOATING
C2663 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n873 GND 0.02fF $ **FLOATING
C2664 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n874 GND 0.05fF $ **FLOATING
C2665 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n875 GND 0.06fF $ **FLOATING
C2666 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n876 GND 0.02fF $ **FLOATING
C2667 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n877 GND 0.05fF $ **FLOATING
C2668 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n878 GND 0.06fF $ **FLOATING
C2669 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n879 GND 0.02fF $ **FLOATING
C2670 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n880 GND 0.05fF $ **FLOATING
C2671 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n881 GND 0.06fF $ **FLOATING
C2672 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t6 GND 0.04fF
C2673 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n882 GND 0.09fF $ **FLOATING
C2674 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n883 GND 0.02fF $ **FLOATING
C2675 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n884 GND 0.03fF $ **FLOATING
C2676 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n885 GND 0.06fF $ **FLOATING
C2677 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n886 GND 0.02fF $ **FLOATING
C2678 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n887 GND 0.04fF $ **FLOATING
C2679 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n888 GND 0.06fF $ **FLOATING
C2680 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t172 GND 0.01fF
C2681 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t196 GND 0.01fF
C2682 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n889 GND 0.04fF $ **FLOATING
C2683 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n890 GND 0.05fF $ **FLOATING
C2684 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n891 GND 0.02fF $ **FLOATING
C2685 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n892 GND 0.04fF $ **FLOATING
C2686 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n893 GND 0.06fF $ **FLOATING
C2687 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n894 GND 0.02fF $ **FLOATING
C2688 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n895 GND 0.04fF $ **FLOATING
C2689 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n896 GND 0.06fF $ **FLOATING
C2690 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n897 GND 0.02fF $ **FLOATING
C2691 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n898 GND 0.05fF $ **FLOATING
C2692 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n899 GND 0.06fF $ **FLOATING
C2693 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n900 GND 0.02fF $ **FLOATING
C2694 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n901 GND 0.05fF $ **FLOATING
C2695 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n902 GND 0.06fF $ **FLOATING
C2696 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n903 GND 0.02fF $ **FLOATING
C2697 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n904 GND 0.05fF $ **FLOATING
C2698 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n905 GND 0.06fF $ **FLOATING
C2699 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t19 GND 0.02fF
C2700 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n906 GND 0.07fF $ **FLOATING
C2701 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n907 GND 0.02fF $ **FLOATING
C2702 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n908 GND 0.03fF $ **FLOATING
C2703 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n909 GND 0.06fF $ **FLOATING
C2704 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n910 GND 0.02fF $ **FLOATING
C2705 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n911 GND 0.04fF $ **FLOATING
C2706 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n912 GND 0.06fF $ **FLOATING
C2707 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n913 GND 0.02fF $ **FLOATING
C2708 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n914 GND 0.05fF $ **FLOATING
C2709 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n915 GND 0.06fF $ **FLOATING
C2710 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t231 GND 0.01fF
C2711 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t38 GND 0.01fF
C2712 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n916 GND 0.04fF $ **FLOATING
C2713 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n917 GND 0.05fF $ **FLOATING
C2714 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n918 GND 0.02fF $ **FLOATING
C2715 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n919 GND 0.03fF $ **FLOATING
C2716 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n920 GND 0.06fF $ **FLOATING
C2717 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n921 GND 0.02fF $ **FLOATING
C2718 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n922 GND 0.05fF $ **FLOATING
C2719 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n923 GND 0.06fF $ **FLOATING
C2720 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n924 GND 0.02fF $ **FLOATING
C2721 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n925 GND 0.05fF $ **FLOATING
C2722 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n926 GND 0.06fF $ **FLOATING
C2723 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t122 GND 0.02fF
C2724 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t124 GND 0.01fF
C2725 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n927 GND 0.10fF $ **FLOATING
C2726 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n928 GND 0.04fF $ **FLOATING
C2727 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n929 GND 0.02fF $ **FLOATING
C2728 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n930 GND 0.03fF $ **FLOATING
C2729 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n931 GND 0.06fF $ **FLOATING
C2730 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n932 GND 0.02fF $ **FLOATING
C2731 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n933 GND 0.05fF $ **FLOATING
C2732 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n934 GND 0.06fF $ **FLOATING
C2733 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n935 GND 0.02fF $ **FLOATING
C2734 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n936 GND 0.05fF $ **FLOATING
C2735 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n937 GND 0.06fF $ **FLOATING
C2736 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n938 GND 0.02fF $ **FLOATING
C2737 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n939 GND 0.04fF $ **FLOATING
C2738 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n940 GND 0.06fF $ **FLOATING
C2739 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t123 GND 0.02fF
C2740 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n941 GND 0.06fF $ **FLOATING
C2741 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n942 GND 0.05fF $ **FLOATING
C2742 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t109 GND 0.01fF
C2743 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n943 GND 0.03fF $ **FLOATING
C2744 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n944 GND 0.05fF $ **FLOATING
C2745 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n945 GND 0.02fF $ **FLOATING
C2746 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n946 GND 0.04fF $ **FLOATING
C2747 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n947 GND 0.06fF $ **FLOATING
C2748 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n948 GND 0.02fF $ **FLOATING
C2749 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n949 GND 0.04fF $ **FLOATING
C2750 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n950 GND 0.06fF $ **FLOATING
C2751 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t163 GND 0.01fF
C2752 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t121 GND 0.02fF
C2753 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n951 GND 0.04fF $ **FLOATING
C2754 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n952 GND 0.04fF $ **FLOATING
C2755 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n953 GND 0.02fF $ **FLOATING
C2756 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n954 GND 0.03fF $ **FLOATING
C2757 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n955 GND 0.06fF $ **FLOATING
C2758 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n956 GND 0.02fF $ **FLOATING
C2759 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n957 GND 0.05fF $ **FLOATING
C2760 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n958 GND 0.06fF $ **FLOATING
C2761 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n959 GND 0.02fF $ **FLOATING
C2762 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n960 GND 0.05fF $ **FLOATING
C2763 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n961 GND 0.06fF $ **FLOATING
C2764 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n962 GND 0.02fF $ **FLOATING
C2765 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n963 GND 0.05fF $ **FLOATING
C2766 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n964 GND 0.06fF $ **FLOATING
C2767 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t197 GND 0.04fF
C2768 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n965 GND 0.09fF $ **FLOATING
C2769 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n966 GND 0.02fF $ **FLOATING
C2770 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n967 GND 0.03fF $ **FLOATING
C2771 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n968 GND 0.06fF $ **FLOATING
C2772 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n969 GND 0.02fF $ **FLOATING
C2773 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n970 GND 0.04fF $ **FLOATING
C2774 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n971 GND 0.06fF $ **FLOATING
C2775 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t181 GND 0.01fF
C2776 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t53 GND 0.01fF
C2777 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n972 GND 0.04fF $ **FLOATING
C2778 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n973 GND 0.05fF $ **FLOATING
C2779 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n974 GND 0.02fF $ **FLOATING
C2780 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n975 GND 0.04fF $ **FLOATING
C2781 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n976 GND 0.06fF $ **FLOATING
C2782 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n977 GND 0.02fF $ **FLOATING
C2783 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n978 GND 0.04fF $ **FLOATING
C2784 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n979 GND 0.06fF $ **FLOATING
C2785 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n980 GND 0.02fF $ **FLOATING
C2786 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n981 GND 0.05fF $ **FLOATING
C2787 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n982 GND 0.06fF $ **FLOATING
C2788 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n983 GND 0.02fF $ **FLOATING
C2789 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n984 GND 0.05fF $ **FLOATING
C2790 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n985 GND 0.06fF $ **FLOATING
C2791 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n986 GND 0.02fF $ **FLOATING
C2792 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n987 GND 0.05fF $ **FLOATING
C2793 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n988 GND 0.06fF $ **FLOATING
C2794 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t37 GND 0.02fF
C2795 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n989 GND 0.07fF $ **FLOATING
C2796 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n990 GND 0.02fF $ **FLOATING
C2797 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n991 GND 0.03fF $ **FLOATING
C2798 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n992 GND 0.06fF $ **FLOATING
C2799 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n993 GND 0.02fF $ **FLOATING
C2800 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n994 GND 0.04fF $ **FLOATING
C2801 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n995 GND 0.06fF $ **FLOATING
C2802 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n996 GND 0.02fF $ **FLOATING
C2803 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n997 GND 0.05fF $ **FLOATING
C2804 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n998 GND 0.06fF $ **FLOATING
C2805 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t135 GND 0.01fF
C2806 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t134 GND 0.01fF
C2807 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n999 GND 0.04fF $ **FLOATING
C2808 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1000 GND 0.05fF $ **FLOATING
C2809 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1001 GND 0.02fF $ **FLOATING
C2810 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1002 GND 0.03fF $ **FLOATING
C2811 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1003 GND 0.06fF $ **FLOATING
C2812 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1004 GND 0.02fF $ **FLOATING
C2813 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1005 GND 0.05fF $ **FLOATING
C2814 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1006 GND 0.06fF $ **FLOATING
C2815 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1007 GND 0.02fF $ **FLOATING
C2816 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1008 GND 0.05fF $ **FLOATING
C2817 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1009 GND 0.06fF $ **FLOATING
C2818 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t139 GND 0.02fF
C2819 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t40 GND 0.01fF
C2820 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1010 GND 0.10fF $ **FLOATING
C2821 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1011 GND 0.04fF $ **FLOATING
C2822 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1012 GND 0.02fF $ **FLOATING
C2823 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1013 GND 0.03fF $ **FLOATING
C2824 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1014 GND 0.06fF $ **FLOATING
C2825 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1015 GND 0.02fF $ **FLOATING
C2826 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1016 GND 0.05fF $ **FLOATING
C2827 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1017 GND 0.06fF $ **FLOATING
C2828 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1018 GND 0.02fF $ **FLOATING
C2829 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1019 GND 0.05fF $ **FLOATING
C2830 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1020 GND 0.06fF $ **FLOATING
C2831 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1021 GND 0.02fF $ **FLOATING
C2832 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1022 GND 0.04fF $ **FLOATING
C2833 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1023 GND 0.06fF $ **FLOATING
C2834 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t140 GND 0.02fF
C2835 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1024 GND 0.06fF $ **FLOATING
C2836 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1025 GND 0.05fF $ **FLOATING
C2837 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t20 GND 0.01fF
C2838 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1026 GND 0.03fF $ **FLOATING
C2839 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1027 GND 0.05fF $ **FLOATING
C2840 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1028 GND 0.02fF $ **FLOATING
C2841 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1029 GND 0.04fF $ **FLOATING
C2842 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1030 GND 0.06fF $ **FLOATING
C2843 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1031 GND 0.02fF $ **FLOATING
C2844 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1032 GND 0.04fF $ **FLOATING
C2845 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1033 GND 0.06fF $ **FLOATING
C2846 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t161 GND 0.01fF
C2847 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t138 GND 0.02fF
C2848 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1034 GND 0.04fF $ **FLOATING
C2849 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1035 GND 0.04fF $ **FLOATING
C2850 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1036 GND 0.02fF $ **FLOATING
C2851 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1037 GND 0.03fF $ **FLOATING
C2852 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1038 GND 0.06fF $ **FLOATING
C2853 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1039 GND 0.02fF $ **FLOATING
C2854 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1040 GND 0.05fF $ **FLOATING
C2855 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1041 GND 0.06fF $ **FLOATING
C2856 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1042 GND 0.02fF $ **FLOATING
C2857 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1043 GND 0.05fF $ **FLOATING
C2858 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1044 GND 0.06fF $ **FLOATING
C2859 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1045 GND 0.02fF $ **FLOATING
C2860 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1046 GND 0.05fF $ **FLOATING
C2861 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1047 GND 0.06fF $ **FLOATING
C2862 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t0 GND 0.04fF
C2863 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1048 GND 0.09fF $ **FLOATING
C2864 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1049 GND 0.02fF $ **FLOATING
C2865 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1050 GND 0.03fF $ **FLOATING
C2866 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1051 GND 0.06fF $ **FLOATING
C2867 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1052 GND 0.02fF $ **FLOATING
C2868 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1053 GND 0.04fF $ **FLOATING
C2869 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1054 GND 0.06fF $ **FLOATING
C2870 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t189 GND 0.01fF
C2871 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t29 GND 0.01fF
C2872 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1055 GND 0.04fF $ **FLOATING
C2873 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1056 GND 0.05fF $ **FLOATING
C2874 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1057 GND 0.02fF $ **FLOATING
C2875 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1058 GND 0.04fF $ **FLOATING
C2876 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1059 GND 0.06fF $ **FLOATING
C2877 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1060 GND 0.02fF $ **FLOATING
C2878 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1061 GND 0.04fF $ **FLOATING
C2879 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1062 GND 0.06fF $ **FLOATING
C2880 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1063 GND 0.02fF $ **FLOATING
C2881 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1064 GND 0.05fF $ **FLOATING
C2882 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1065 GND 0.06fF $ **FLOATING
C2883 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1066 GND 0.02fF $ **FLOATING
C2884 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1067 GND 0.05fF $ **FLOATING
C2885 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1068 GND 0.06fF $ **FLOATING
C2886 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1069 GND 0.02fF $ **FLOATING
C2887 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1070 GND 0.05fF $ **FLOATING
C2888 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1071 GND 0.06fF $ **FLOATING
C2889 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t133 GND 0.02fF
C2890 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1072 GND 0.07fF $ **FLOATING
C2891 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1073 GND 0.02fF $ **FLOATING
C2892 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1074 GND 0.03fF $ **FLOATING
C2893 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1075 GND 0.06fF $ **FLOATING
C2894 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1076 GND 0.02fF $ **FLOATING
C2895 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1077 GND 0.04fF $ **FLOATING
C2896 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1078 GND 0.06fF $ **FLOATING
C2897 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1079 GND 0.02fF $ **FLOATING
C2898 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1080 GND 0.05fF $ **FLOATING
C2899 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1081 GND 0.06fF $ **FLOATING
C2900 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t144 GND 0.01fF
C2901 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t214 GND 0.01fF
C2902 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1082 GND 0.04fF $ **FLOATING
C2903 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1083 GND 0.05fF $ **FLOATING
C2904 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1084 GND 0.02fF $ **FLOATING
C2905 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1085 GND 0.03fF $ **FLOATING
C2906 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1086 GND 0.06fF $ **FLOATING
C2907 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1087 GND 0.02fF $ **FLOATING
C2908 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1088 GND 0.05fF $ **FLOATING
C2909 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1089 GND 0.06fF $ **FLOATING
C2910 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1090 GND 0.02fF $ **FLOATING
C2911 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1091 GND 0.05fF $ **FLOATING
C2912 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1092 GND 0.06fF $ **FLOATING
C2913 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t62 GND 0.02fF
C2914 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t88 GND 0.01fF
C2915 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1093 GND 0.10fF $ **FLOATING
C2916 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1094 GND 0.04fF $ **FLOATING
C2917 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1095 GND 0.02fF $ **FLOATING
C2918 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1096 GND 0.03fF $ **FLOATING
C2919 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1097 GND 0.06fF $ **FLOATING
C2920 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1098 GND 0.02fF $ **FLOATING
C2921 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1099 GND 0.05fF $ **FLOATING
C2922 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1100 GND 0.06fF $ **FLOATING
C2923 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1101 GND 0.02fF $ **FLOATING
C2924 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1102 GND 0.05fF $ **FLOATING
C2925 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1103 GND 0.06fF $ **FLOATING
C2926 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1104 GND 0.02fF $ **FLOATING
C2927 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1105 GND 0.04fF $ **FLOATING
C2928 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1106 GND 0.06fF $ **FLOATING
C2929 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t63 GND 0.02fF
C2930 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1107 GND 0.06fF $ **FLOATING
C2931 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1108 GND 0.05fF $ **FLOATING
C2932 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t90 GND 0.01fF
C2933 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1109 GND 0.03fF $ **FLOATING
C2934 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1110 GND 0.05fF $ **FLOATING
C2935 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1111 GND 0.02fF $ **FLOATING
C2936 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1112 GND 0.04fF $ **FLOATING
C2937 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1113 GND 0.06fF $ **FLOATING
C2938 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1114 GND 0.02fF $ **FLOATING
C2939 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1115 GND 0.04fF $ **FLOATING
C2940 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1116 GND 0.06fF $ **FLOATING
C2941 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t157 GND 0.01fF
C2942 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t61 GND 0.02fF
C2943 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1117 GND 0.04fF $ **FLOATING
C2944 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1118 GND 0.04fF $ **FLOATING
C2945 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1119 GND 0.02fF $ **FLOATING
C2946 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1120 GND 0.03fF $ **FLOATING
C2947 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1121 GND 0.06fF $ **FLOATING
C2948 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1122 GND 0.02fF $ **FLOATING
C2949 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1123 GND 0.05fF $ **FLOATING
C2950 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1124 GND 0.06fF $ **FLOATING
C2951 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1125 GND 0.02fF $ **FLOATING
C2952 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1126 GND 0.05fF $ **FLOATING
C2953 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1127 GND 0.06fF $ **FLOATING
C2954 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1128 GND 0.02fF $ **FLOATING
C2955 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1129 GND 0.05fF $ **FLOATING
C2956 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1130 GND 0.06fF $ **FLOATING
C2957 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t39 GND 0.04fF
C2958 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1131 GND 0.09fF $ **FLOATING
C2959 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1132 GND 0.02fF $ **FLOATING
C2960 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1133 GND 0.03fF $ **FLOATING
C2961 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1134 GND 0.06fF $ **FLOATING
C2962 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1135 GND 0.02fF $ **FLOATING
C2963 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1136 GND 0.04fF $ **FLOATING
C2964 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1137 GND 0.06fF $ **FLOATING
C2965 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t186 GND 0.01fF
C2966 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t96 GND 0.01fF
C2967 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1138 GND 0.04fF $ **FLOATING
C2968 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1139 GND 0.05fF $ **FLOATING
C2969 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1140 GND 0.02fF $ **FLOATING
C2970 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1141 GND 0.04fF $ **FLOATING
C2971 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1142 GND 0.06fF $ **FLOATING
C2972 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1143 GND 0.02fF $ **FLOATING
C2973 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1144 GND 0.04fF $ **FLOATING
C2974 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1145 GND 0.06fF $ **FLOATING
C2975 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1146 GND 0.02fF $ **FLOATING
C2976 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1147 GND 0.05fF $ **FLOATING
C2977 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1148 GND 0.06fF $ **FLOATING
C2978 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1149 GND 0.02fF $ **FLOATING
C2979 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1150 GND 0.05fF $ **FLOATING
C2980 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1151 GND 0.06fF $ **FLOATING
C2981 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1152 GND 0.02fF $ **FLOATING
C2982 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1153 GND 0.05fF $ **FLOATING
C2983 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1154 GND 0.06fF $ **FLOATING
C2984 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t213 GND 0.02fF
C2985 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1155 GND 0.07fF $ **FLOATING
C2986 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1156 GND 0.02fF $ **FLOATING
C2987 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1157 GND 0.03fF $ **FLOATING
C2988 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1158 GND 0.06fF $ **FLOATING
C2989 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1159 GND 0.02fF $ **FLOATING
C2990 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1160 GND 0.04fF $ **FLOATING
C2991 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1161 GND 0.06fF $ **FLOATING
C2992 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1162 GND 0.02fF $ **FLOATING
C2993 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1163 GND 0.05fF $ **FLOATING
C2994 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1164 GND 0.06fF $ **FLOATING
C2995 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t239 GND 0.01fF
C2996 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t147 GND 0.01fF
C2997 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1165 GND 0.04fF $ **FLOATING
C2998 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1166 GND 0.05fF $ **FLOATING
C2999 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1167 GND 0.02fF $ **FLOATING
C3000 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1168 GND 0.03fF $ **FLOATING
C3001 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1169 GND 0.06fF $ **FLOATING
C3002 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1170 GND 0.02fF $ **FLOATING
C3003 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1171 GND 0.05fF $ **FLOATING
C3004 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1172 GND 0.06fF $ **FLOATING
C3005 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1173 GND 0.02fF $ **FLOATING
C3006 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1174 GND 0.05fF $ **FLOATING
C3007 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1175 GND 0.06fF $ **FLOATING
C3008 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t116 GND 0.02fF
C3009 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t207 GND 0.01fF
C3010 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1176 GND 0.10fF $ **FLOATING
C3011 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1177 GND 0.04fF $ **FLOATING
C3012 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1178 GND 0.02fF $ **FLOATING
C3013 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1179 GND 0.03fF $ **FLOATING
C3014 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1180 GND 0.06fF $ **FLOATING
C3015 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1181 GND 0.02fF $ **FLOATING
C3016 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1182 GND 0.05fF $ **FLOATING
C3017 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1183 GND 0.06fF $ **FLOATING
C3018 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1184 GND 0.02fF $ **FLOATING
C3019 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1185 GND 0.05fF $ **FLOATING
C3020 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1186 GND 0.06fF $ **FLOATING
C3021 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1187 GND 0.02fF $ **FLOATING
C3022 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1188 GND 0.04fF $ **FLOATING
C3023 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1189 GND 0.06fF $ **FLOATING
C3024 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t114 GND 0.02fF
C3025 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1190 GND 0.06fF $ **FLOATING
C3026 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1191 GND 0.05fF $ **FLOATING
C3027 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t23 GND 0.01fF
C3028 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1192 GND 0.03fF $ **FLOATING
C3029 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1193 GND 0.05fF $ **FLOATING
C3030 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1194 GND 0.02fF $ **FLOATING
C3031 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1195 GND 0.04fF $ **FLOATING
C3032 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1196 GND 0.06fF $ **FLOATING
C3033 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1197 GND 0.02fF $ **FLOATING
C3034 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1198 GND 0.04fF $ **FLOATING
C3035 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1199 GND 0.06fF $ **FLOATING
C3036 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t165 GND 0.01fF
C3037 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t115 GND 0.02fF
C3038 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1200 GND 0.04fF $ **FLOATING
C3039 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1201 GND 0.04fF $ **FLOATING
C3040 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1202 GND 0.02fF $ **FLOATING
C3041 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1203 GND 0.03fF $ **FLOATING
C3042 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1204 GND 0.06fF $ **FLOATING
C3043 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1205 GND 0.02fF $ **FLOATING
C3044 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1206 GND 0.05fF $ **FLOATING
C3045 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1207 GND 0.06fF $ **FLOATING
C3046 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1208 GND 0.02fF $ **FLOATING
C3047 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1209 GND 0.05fF $ **FLOATING
C3048 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1210 GND 0.06fF $ **FLOATING
C3049 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1211 GND 0.02fF $ **FLOATING
C3050 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1212 GND 0.05fF $ **FLOATING
C3051 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1213 GND 0.06fF $ **FLOATING
C3052 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t126 GND 0.04fF
C3053 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1214 GND 0.09fF $ **FLOATING
C3054 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1215 GND 0.02fF $ **FLOATING
C3055 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1216 GND 0.03fF $ **FLOATING
C3056 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1217 GND 0.06fF $ **FLOATING
C3057 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1218 GND 0.02fF $ **FLOATING
C3058 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1219 GND 0.04fF $ **FLOATING
C3059 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1220 GND 0.06fF $ **FLOATING
C3060 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t183 GND 0.01fF
C3061 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t30 GND 0.01fF
C3062 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1221 GND 0.04fF $ **FLOATING
C3063 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1222 GND 0.05fF $ **FLOATING
C3064 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1223 GND 0.02fF $ **FLOATING
C3065 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1224 GND 0.04fF $ **FLOATING
C3066 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1225 GND 0.06fF $ **FLOATING
C3067 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1226 GND 0.02fF $ **FLOATING
C3068 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1227 GND 0.04fF $ **FLOATING
C3069 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1228 GND 0.06fF $ **FLOATING
C3070 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1229 GND 0.02fF $ **FLOATING
C3071 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1230 GND 0.05fF $ **FLOATING
C3072 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1231 GND 0.06fF $ **FLOATING
C3073 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1232 GND 0.02fF $ **FLOATING
C3074 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1233 GND 0.05fF $ **FLOATING
C3075 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1234 GND 0.06fF $ **FLOATING
C3076 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1235 GND 0.02fF $ **FLOATING
C3077 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1236 GND 0.05fF $ **FLOATING
C3078 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1237 GND 0.06fF $ **FLOATING
C3079 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t146 GND 0.02fF
C3080 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1238 GND 0.07fF $ **FLOATING
C3081 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1239 GND 0.02fF $ **FLOATING
C3082 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1240 GND 0.03fF $ **FLOATING
C3083 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1241 GND 0.06fF $ **FLOATING
C3084 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1242 GND 0.02fF $ **FLOATING
C3085 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1243 GND 0.04fF $ **FLOATING
C3086 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1244 GND 0.06fF $ **FLOATING
C3087 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1245 GND 0.02fF $ **FLOATING
C3088 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1246 GND 0.05fF $ **FLOATING
C3089 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1247 GND 0.06fF $ **FLOATING
C3090 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t22 GND 0.01fF
C3091 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t119 GND 0.01fF
C3092 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1248 GND 0.04fF $ **FLOATING
C3093 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1249 GND 0.05fF $ **FLOATING
C3094 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1250 GND 0.02fF $ **FLOATING
C3095 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1251 GND 0.03fF $ **FLOATING
C3096 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1252 GND 0.06fF $ **FLOATING
C3097 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1253 GND 0.02fF $ **FLOATING
C3098 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1254 GND 0.05fF $ **FLOATING
C3099 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1255 GND 0.06fF $ **FLOATING
C3100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1256 GND 0.02fF $ **FLOATING
C3101 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1257 GND 0.05fF $ **FLOATING
C3102 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1258 GND 0.06fF $ **FLOATING
C3103 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t59 GND 0.02fF
C3104 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t128 GND 0.01fF
C3105 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1259 GND 0.10fF $ **FLOATING
C3106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1260 GND 0.04fF $ **FLOATING
C3107 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1261 GND 0.02fF $ **FLOATING
C3108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1262 GND 0.03fF $ **FLOATING
C3109 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1263 GND 0.06fF $ **FLOATING
C3110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1264 GND 0.02fF $ **FLOATING
C3111 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1265 GND 0.05fF $ **FLOATING
C3112 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1266 GND 0.06fF $ **FLOATING
C3113 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1267 GND 0.02fF $ **FLOATING
C3114 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1268 GND 0.05fF $ **FLOATING
C3115 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1269 GND 0.06fF $ **FLOATING
C3116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1270 GND 0.02fF $ **FLOATING
C3117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1271 GND 0.04fF $ **FLOATING
C3118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1272 GND 0.06fF $ **FLOATING
C3119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t60 GND 0.02fF
C3120 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1273 GND 0.06fF $ **FLOATING
C3121 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1274 GND 0.05fF $ **FLOATING
C3122 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t13 GND 0.01fF
C3123 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1275 GND 0.03fF $ **FLOATING
C3124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1276 GND 0.05fF $ **FLOATING
C3125 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1277 GND 0.02fF $ **FLOATING
C3126 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1278 GND 0.04fF $ **FLOATING
C3127 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1279 GND 0.06fF $ **FLOATING
C3128 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1280 GND 0.02fF $ **FLOATING
C3129 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1281 GND 0.04fF $ **FLOATING
C3130 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1282 GND 0.06fF $ **FLOATING
C3131 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t158 GND 0.01fF
C3132 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t58 GND 0.02fF
C3133 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1283 GND 0.04fF $ **FLOATING
C3134 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1284 GND 0.04fF $ **FLOATING
C3135 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1285 GND 0.02fF $ **FLOATING
C3136 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1286 GND 0.03fF $ **FLOATING
C3137 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1287 GND 0.06fF $ **FLOATING
C3138 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1288 GND 0.02fF $ **FLOATING
C3139 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1289 GND 0.05fF $ **FLOATING
C3140 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1290 GND 0.06fF $ **FLOATING
C3141 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1291 GND 0.02fF $ **FLOATING
C3142 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1292 GND 0.05fF $ **FLOATING
C3143 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1293 GND 0.06fF $ **FLOATING
C3144 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1294 GND 0.02fF $ **FLOATING
C3145 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1295 GND 0.05fF $ **FLOATING
C3146 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1296 GND 0.06fF $ **FLOATING
C3147 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t44 GND 0.04fF
C3148 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1297 GND 0.09fF $ **FLOATING
C3149 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1298 GND 0.02fF $ **FLOATING
C3150 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1299 GND 0.03fF $ **FLOATING
C3151 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1300 GND 0.06fF $ **FLOATING
C3152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1301 GND 0.02fF $ **FLOATING
C3153 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1302 GND 0.04fF $ **FLOATING
C3154 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1303 GND 0.06fF $ **FLOATING
C3155 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t184 GND 0.01fF
C3156 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t21 GND 0.01fF
C3157 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1304 GND 0.04fF $ **FLOATING
C3158 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1305 GND 0.05fF $ **FLOATING
C3159 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1306 GND 0.02fF $ **FLOATING
C3160 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1307 GND 0.04fF $ **FLOATING
C3161 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1308 GND 0.06fF $ **FLOATING
C3162 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1309 GND 0.02fF $ **FLOATING
C3163 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1310 GND 0.04fF $ **FLOATING
C3164 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1311 GND 0.06fF $ **FLOATING
C3165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1312 GND 0.02fF $ **FLOATING
C3166 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1313 GND 0.05fF $ **FLOATING
C3167 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1314 GND 0.06fF $ **FLOATING
C3168 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1315 GND 0.02fF $ **FLOATING
C3169 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1316 GND 0.05fF $ **FLOATING
C3170 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1317 GND 0.06fF $ **FLOATING
C3171 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1318 GND 0.02fF $ **FLOATING
C3172 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1319 GND 0.05fF $ **FLOATING
C3173 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1320 GND 0.06fF $ **FLOATING
C3174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t118 GND 0.02fF
C3175 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1321 GND 0.07fF $ **FLOATING
C3176 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1322 GND 0.02fF $ **FLOATING
C3177 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1323 GND 0.03fF $ **FLOATING
C3178 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1324 GND 0.06fF $ **FLOATING
C3179 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1325 GND 0.02fF $ **FLOATING
C3180 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1326 GND 0.04fF $ **FLOATING
C3181 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1327 GND 0.06fF $ **FLOATING
C3182 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1328 GND 0.02fF $ **FLOATING
C3183 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1329 GND 0.05fF $ **FLOATING
C3184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1330 GND 0.06fF $ **FLOATING
C3185 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t233 GND 0.01fF
C3186 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t149 GND 0.01fF
C3187 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1331 GND 0.04fF $ **FLOATING
C3188 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1332 GND 0.05fF $ **FLOATING
C3189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1333 GND 0.02fF $ **FLOATING
C3190 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1334 GND 0.03fF $ **FLOATING
C3191 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1335 GND 0.06fF $ **FLOATING
C3192 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1336 GND 0.02fF $ **FLOATING
C3193 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1337 GND 0.05fF $ **FLOATING
C3194 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1338 GND 0.06fF $ **FLOATING
C3195 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1339 GND 0.02fF $ **FLOATING
C3196 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1340 GND 0.05fF $ **FLOATING
C3197 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1341 GND 0.06fF $ **FLOATING
C3198 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t33 GND 0.02fF
C3199 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t77 GND 0.01fF
C3200 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1342 GND 0.10fF $ **FLOATING
C3201 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1343 GND 0.04fF $ **FLOATING
C3202 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1344 GND 0.02fF $ **FLOATING
C3203 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1345 GND 0.03fF $ **FLOATING
C3204 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1346 GND 0.06fF $ **FLOATING
C3205 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1347 GND 0.02fF $ **FLOATING
C3206 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1348 GND 0.05fF $ **FLOATING
C3207 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1349 GND 0.06fF $ **FLOATING
C3208 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1350 GND 0.02fF $ **FLOATING
C3209 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1351 GND 0.05fF $ **FLOATING
C3210 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1352 GND 0.06fF $ **FLOATING
C3211 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1353 GND 0.02fF $ **FLOATING
C3212 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1354 GND 0.04fF $ **FLOATING
C3213 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1355 GND 0.06fF $ **FLOATING
C3214 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t34 GND 0.02fF
C3215 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1356 GND 0.06fF $ **FLOATING
C3216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1357 GND 0.05fF $ **FLOATING
C3217 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t203 GND 0.01fF
C3218 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1358 GND 0.03fF $ **FLOATING
C3219 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1359 GND 0.05fF $ **FLOATING
C3220 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1360 GND 0.02fF $ **FLOATING
C3221 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1361 GND 0.04fF $ **FLOATING
C3222 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1362 GND 0.06fF $ **FLOATING
C3223 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1363 GND 0.02fF $ **FLOATING
C3224 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1364 GND 0.04fF $ **FLOATING
C3225 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1365 GND 0.06fF $ **FLOATING
C3226 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t166 GND 0.01fF
C3227 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t32 GND 0.02fF
C3228 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1366 GND 0.04fF $ **FLOATING
C3229 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1367 GND 0.04fF $ **FLOATING
C3230 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1368 GND 0.02fF $ **FLOATING
C3231 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1369 GND 0.03fF $ **FLOATING
C3232 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1370 GND 0.06fF $ **FLOATING
C3233 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1371 GND 0.02fF $ **FLOATING
C3234 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1372 GND 0.05fF $ **FLOATING
C3235 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1373 GND 0.06fF $ **FLOATING
C3236 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1374 GND 0.02fF $ **FLOATING
C3237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1375 GND 0.05fF $ **FLOATING
C3238 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1376 GND 0.06fF $ **FLOATING
C3239 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1377 GND 0.02fF $ **FLOATING
C3240 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1378 GND 0.05fF $ **FLOATING
C3241 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1379 GND 0.06fF $ **FLOATING
C3242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t86 GND 0.04fF
C3243 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1380 GND 0.09fF $ **FLOATING
C3244 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1381 GND 0.02fF $ **FLOATING
C3245 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1382 GND 0.03fF $ **FLOATING
C3246 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1383 GND 0.06fF $ **FLOATING
C3247 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1384 GND 0.02fF $ **FLOATING
C3248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1385 GND 0.04fF $ **FLOATING
C3249 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1386 GND 0.06fF $ **FLOATING
C3250 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t182 GND 0.01fF
C3251 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t41 GND 0.01fF
C3252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1387 GND 0.04fF $ **FLOATING
C3253 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1388 GND 0.05fF $ **FLOATING
C3254 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1389 GND 0.02fF $ **FLOATING
C3255 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1390 GND 0.04fF $ **FLOATING
C3256 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1391 GND 0.06fF $ **FLOATING
C3257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1392 GND 0.02fF $ **FLOATING
C3258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1393 GND 0.04fF $ **FLOATING
C3259 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1394 GND 0.06fF $ **FLOATING
C3260 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1395 GND 0.02fF $ **FLOATING
C3261 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1396 GND 0.05fF $ **FLOATING
C3262 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1397 GND 0.06fF $ **FLOATING
C3263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1398 GND 0.02fF $ **FLOATING
C3264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1399 GND 0.05fF $ **FLOATING
C3265 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1400 GND 0.06fF $ **FLOATING
C3266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1401 GND 0.02fF $ **FLOATING
C3267 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1402 GND 0.05fF $ **FLOATING
C3268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1403 GND 0.06fF $ **FLOATING
C3269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t148 GND 0.02fF
C3270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1404 GND 0.07fF $ **FLOATING
C3271 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1405 GND 0.02fF $ **FLOATING
C3272 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1406 GND 0.03fF $ **FLOATING
C3273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1407 GND 0.06fF $ **FLOATING
C3274 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1408 GND 0.02fF $ **FLOATING
C3275 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1409 GND 0.04fF $ **FLOATING
C3276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1410 GND 0.06fF $ **FLOATING
C3277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1411 GND 0.02fF $ **FLOATING
C3278 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1412 GND 0.05fF $ **FLOATING
C3279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1413 GND 0.06fF $ **FLOATING
C3280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t210 GND 0.01fF
C3281 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t202 GND 0.01fF
C3282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1414 GND 0.04fF $ **FLOATING
C3283 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1415 GND 0.05fF $ **FLOATING
C3284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1416 GND 0.02fF $ **FLOATING
C3285 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1417 GND 0.03fF $ **FLOATING
C3286 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1418 GND 0.06fF $ **FLOATING
C3287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1419 GND 0.02fF $ **FLOATING
C3288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1420 GND 0.05fF $ **FLOATING
C3289 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1421 GND 0.06fF $ **FLOATING
C3290 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1422 GND 0.02fF $ **FLOATING
C3291 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1423 GND 0.05fF $ **FLOATING
C3292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1424 GND 0.06fF $ **FLOATING
C3293 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t236 GND 0.02fF
C3294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t14 GND 0.01fF
C3295 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1425 GND 0.10fF $ **FLOATING
C3296 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1426 GND 0.04fF $ **FLOATING
C3297 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1427 GND 0.02fF $ **FLOATING
C3298 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1428 GND 0.03fF $ **FLOATING
C3299 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1429 GND 0.06fF $ **FLOATING
C3300 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1430 GND 0.02fF $ **FLOATING
C3301 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1431 GND 0.05fF $ **FLOATING
C3302 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1432 GND 0.06fF $ **FLOATING
C3303 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1433 GND 0.02fF $ **FLOATING
C3304 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1434 GND 0.05fF $ **FLOATING
C3305 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1435 GND 0.06fF $ **FLOATING
C3306 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1436 GND 0.02fF $ **FLOATING
C3307 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1437 GND 0.04fF $ **FLOATING
C3308 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1438 GND 0.06fF $ **FLOATING
C3309 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t235 GND 0.02fF
C3310 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1439 GND 0.06fF $ **FLOATING
C3311 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1440 GND 0.05fF $ **FLOATING
C3312 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t117 GND 0.01fF
C3313 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1441 GND 0.03fF $ **FLOATING
C3314 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1442 GND 0.05fF $ **FLOATING
C3315 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1443 GND 0.02fF $ **FLOATING
C3316 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1444 GND 0.04fF $ **FLOATING
C3317 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1445 GND 0.06fF $ **FLOATING
C3318 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1446 GND 0.02fF $ **FLOATING
C3319 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1447 GND 0.04fF $ **FLOATING
C3320 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1448 GND 0.06fF $ **FLOATING
C3321 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t162 GND 0.01fF
C3322 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t234 GND 0.02fF
C3323 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1449 GND 0.04fF $ **FLOATING
C3324 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1450 GND 0.04fF $ **FLOATING
C3325 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1451 GND 0.02fF $ **FLOATING
C3326 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1452 GND 0.03fF $ **FLOATING
C3327 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1453 GND 0.06fF $ **FLOATING
C3328 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1454 GND 0.02fF $ **FLOATING
C3329 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1455 GND 0.05fF $ **FLOATING
C3330 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1456 GND 0.06fF $ **FLOATING
C3331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1457 GND 0.02fF $ **FLOATING
C3332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1458 GND 0.05fF $ **FLOATING
C3333 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1459 GND 0.06fF $ **FLOATING
C3334 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1460 GND 0.02fF $ **FLOATING
C3335 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1461 GND 0.05fF $ **FLOATING
C3336 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1462 GND 0.06fF $ **FLOATING
C3337 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t215 GND 0.04fF
C3338 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1463 GND 0.09fF $ **FLOATING
C3339 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1464 GND 0.02fF $ **FLOATING
C3340 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1465 GND 0.03fF $ **FLOATING
C3341 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1466 GND 0.06fF $ **FLOATING
C3342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1467 GND 0.02fF $ **FLOATING
C3343 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1468 GND 0.04fF $ **FLOATING
C3344 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1469 GND 0.06fF $ **FLOATING
C3345 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t194 GND 0.01fF
C3346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t31 GND 0.01fF
C3347 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1470 GND 0.04fF $ **FLOATING
C3348 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1471 GND 0.05fF $ **FLOATING
C3349 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1472 GND 0.02fF $ **FLOATING
C3350 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1473 GND 0.04fF $ **FLOATING
C3351 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1474 GND 0.06fF $ **FLOATING
C3352 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1475 GND 0.02fF $ **FLOATING
C3353 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1476 GND 0.04fF $ **FLOATING
C3354 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1477 GND 0.06fF $ **FLOATING
C3355 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1478 GND 0.02fF $ **FLOATING
C3356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1479 GND 0.05fF $ **FLOATING
C3357 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1480 GND 0.06fF $ **FLOATING
C3358 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1481 GND 0.02fF $ **FLOATING
C3359 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1482 GND 0.05fF $ **FLOATING
C3360 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1483 GND 0.06fF $ **FLOATING
C3361 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1484 GND 0.02fF $ **FLOATING
C3362 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1485 GND 0.05fF $ **FLOATING
C3363 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1486 GND 0.06fF $ **FLOATING
C3364 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1487 GND 0.06fF $ **FLOATING
C3365 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1488 GND 0.06fF $ **FLOATING
C3366 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1489 GND 0.06fF $ **FLOATING
C3367 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1490 GND 0.06fF $ **FLOATING
C3368 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1491 GND 0.06fF $ **FLOATING
C3369 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1492 GND 0.06fF $ **FLOATING
C3370 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1493 GND 0.07fF $ **FLOATING
C3371 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t85 GND 0.01fF
C3372 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t217 GND 0.01fF
C3373 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1494 GND 0.04fF $ **FLOATING
C3374 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1495 GND 0.05fF $ **FLOATING
C3375 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1496 GND 0.02fF $ **FLOATING
C3376 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1497 GND 0.03fF $ **FLOATING
C3377 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1498 GND 0.13fF $ **FLOATING
C3378 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1499 GND 0.02fF $ **FLOATING
C3379 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1500 GND 0.05fF $ **FLOATING
C3380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1501 GND 0.06fF $ **FLOATING
C3381 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1502 GND 0.02fF $ **FLOATING
C3382 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1503 GND 0.04fF $ **FLOATING
C3383 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1504 GND 0.06fF $ **FLOATING
C3384 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t130 GND 0.02fF
C3385 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1505 GND 0.07fF $ **FLOATING
C3386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1506 GND 0.02fF $ **FLOATING
C3387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1507 GND 0.03fF $ **FLOATING
C3388 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1508 GND 0.06fF $ **FLOATING
C3389 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1509 GND 0.02fF $ **FLOATING
C3390 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1510 GND 0.05fF $ **FLOATING
C3391 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1511 GND 0.06fF $ **FLOATING
C3392 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1512 GND 0.02fF $ **FLOATING
C3393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1513 GND 0.05fF $ **FLOATING
C3394 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1514 GND 0.06fF $ **FLOATING
C3395 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1515 GND 0.02fF $ **FLOATING
C3396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1516 GND 0.05fF $ **FLOATING
C3397 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1517 GND 0.06fF $ **FLOATING
C3398 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1518 GND 0.02fF $ **FLOATING
C3399 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1519 GND 0.04fF $ **FLOATING
C3400 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1520 GND 0.06fF $ **FLOATING
C3401 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t156 GND 0.01fF
C3402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t9 GND 0.01fF
C3403 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1521 GND 0.04fF $ **FLOATING
C3404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1522 GND 0.05fF $ **FLOATING
C3405 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1523 GND 0.02fF $ **FLOATING
C3406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1524 GND 0.04fF $ **FLOATING
C3407 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1525 GND 0.06fF $ **FLOATING
C3408 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1526 GND 0.02fF $ **FLOATING
C3409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1527 GND 0.04fF $ **FLOATING
C3410 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1528 GND 0.06fF $ **FLOATING
C3411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t205 GND 0.04fF
C3412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1529 GND 0.09fF $ **FLOATING
C3413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1530 GND 0.02fF $ **FLOATING
C3414 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1531 GND 0.03fF $ **FLOATING
C3415 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1532 GND 0.06fF $ **FLOATING
C3416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1533 GND 0.02fF $ **FLOATING
C3417 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1534 GND 0.05fF $ **FLOATING
C3418 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1535 GND 0.06fF $ **FLOATING
C3419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1536 GND 0.02fF $ **FLOATING
C3420 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1537 GND 0.05fF $ **FLOATING
C3421 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1538 GND 0.06fF $ **FLOATING
C3422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1539 GND 0.02fF $ **FLOATING
C3423 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1540 GND 0.05fF $ **FLOATING
C3424 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1541 GND 0.06fF $ **FLOATING
C3425 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t167 GND 0.01fF
C3426 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t46 GND 0.02fF
C3427 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1542 GND 0.04fF $ **FLOATING
C3428 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1543 GND 0.04fF $ **FLOATING
C3429 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1544 GND 0.02fF $ **FLOATING
C3430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1545 GND 0.03fF $ **FLOATING
C3431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1546 GND 0.06fF $ **FLOATING
C3432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1547 GND 0.02fF $ **FLOATING
C3433 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1548 GND 0.04fF $ **FLOATING
C3434 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1549 GND 0.06fF $ **FLOATING
C3435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t45 GND 0.02fF
C3436 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1550 GND 0.06fF $ **FLOATING
C3437 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1551 GND 0.05fF $ **FLOATING
C3438 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t137 GND 0.01fF
C3439 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1552 GND 0.03fF $ **FLOATING
C3440 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1553 GND 0.05fF $ **FLOATING
C3441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1554 GND 0.02fF $ **FLOATING
C3442 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1555 GND 0.04fF $ **FLOATING
C3443 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1556 GND 0.06fF $ **FLOATING
C3444 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1557 GND 0.02fF $ **FLOATING
C3445 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1558 GND 0.04fF $ **FLOATING
C3446 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1559 GND 0.06fF $ **FLOATING
C3447 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1560 GND 0.02fF $ **FLOATING
C3448 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1561 GND 0.05fF $ **FLOATING
C3449 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1562 GND 0.06fF $ **FLOATING
C3450 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1563 GND 0.02fF $ **FLOATING
C3451 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1564 GND 0.05fF $ **FLOATING
C3452 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1565 GND 0.06fF $ **FLOATING
C3453 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t47 GND 0.02fF
C3454 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t211 GND 0.01fF
C3455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1566 GND 0.10fF $ **FLOATING
C3456 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1567 GND 0.04fF $ **FLOATING
C3457 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1568 GND 0.02fF $ **FLOATING
C3458 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1569 GND 0.03fF $ **FLOATING
C3459 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1570 GND 0.06fF $ **FLOATING
C3460 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1571 GND 0.02fF $ **FLOATING
C3461 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1572 GND 0.05fF $ **FLOATING
C3462 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1573 GND 0.06fF $ **FLOATING
C3463 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1574 GND 0.02fF $ **FLOATING
C3464 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1575 GND 0.05fF $ **FLOATING
C3465 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1576 GND 0.06fF $ **FLOATING
C3466 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t95 GND 0.01fF
C3467 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t131 GND 0.01fF
C3468 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1577 GND 0.04fF $ **FLOATING
C3469 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1578 GND 0.05fF $ **FLOATING
C3470 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1579 GND 0.02fF $ **FLOATING
C3471 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1580 GND 0.03fF $ **FLOATING
C3472 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1581 GND 0.06fF $ **FLOATING
C3473 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1582 GND 0.02fF $ **FLOATING
C3474 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1583 GND 0.05fF $ **FLOATING
C3475 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1584 GND 0.06fF $ **FLOATING
C3476 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1585 GND 0.02fF $ **FLOATING
C3477 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1586 GND 0.04fF $ **FLOATING
C3478 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1587 GND 0.06fF $ **FLOATING
C3479 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t4 GND 0.02fF
C3480 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1588 GND 0.07fF $ **FLOATING
C3481 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1589 GND 0.02fF $ **FLOATING
C3482 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1590 GND 0.03fF $ **FLOATING
C3483 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1591 GND 0.06fF $ **FLOATING
C3484 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1592 GND 0.02fF $ **FLOATING
C3485 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1593 GND 0.05fF $ **FLOATING
C3486 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1594 GND 0.06fF $ **FLOATING
C3487 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1595 GND 0.02fF $ **FLOATING
C3488 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1596 GND 0.05fF $ **FLOATING
C3489 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1597 GND 0.06fF $ **FLOATING
C3490 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1598 GND 0.02fF $ **FLOATING
C3491 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1599 GND 0.05fF $ **FLOATING
C3492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1600 GND 0.06fF $ **FLOATING
C3493 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1601 GND 0.02fF $ **FLOATING
C3494 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1602 GND 0.04fF $ **FLOATING
C3495 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1603 GND 0.06fF $ **FLOATING
C3496 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t187 GND 0.01fF
C3497 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t132 GND 0.01fF
C3498 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1604 GND 0.04fF $ **FLOATING
C3499 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1605 GND 0.05fF $ **FLOATING
C3500 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1606 GND 0.02fF $ **FLOATING
C3501 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1607 GND 0.04fF $ **FLOATING
C3502 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1608 GND 0.06fF $ **FLOATING
C3503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1609 GND 0.02fF $ **FLOATING
C3504 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1610 GND 0.04fF $ **FLOATING
C3505 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1611 GND 0.06fF $ **FLOATING
C3506 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t84 GND 0.04fF
C3507 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1612 GND 0.09fF $ **FLOATING
C3508 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1613 GND 0.02fF $ **FLOATING
C3509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1614 GND 0.03fF $ **FLOATING
C3510 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1615 GND 0.06fF $ **FLOATING
C3511 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1616 GND 0.02fF $ **FLOATING
C3512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1617 GND 0.05fF $ **FLOATING
C3513 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1618 GND 0.06fF $ **FLOATING
C3514 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1619 GND 0.02fF $ **FLOATING
C3515 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1620 GND 0.05fF $ **FLOATING
C3516 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1621 GND 0.06fF $ **FLOATING
C3517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1622 GND 0.06fF $ **FLOATING
C3518 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1623 GND 0.06fF $ **FLOATING
C3519 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1624 GND 0.06fF $ **FLOATING
C3520 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1625 GND 0.06fF $ **FLOATING
C3521 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1626 GND 0.06fF $ **FLOATING
C3522 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1627 GND 0.06fF $ **FLOATING
C3523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1628 GND 0.06fF $ **FLOATING
C3524 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1629 GND 0.06fF $ **FLOATING
C3525 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1630 GND 0.03fF $ **FLOATING
C3526 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t125 GND 0.01fF
C3527 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1631 GND 0.03fF $ **FLOATING
C3528 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t159 GND 0.01fF
C3529 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t225 GND 0.02fF
C3530 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1632 GND 0.04fF $ **FLOATING
C3531 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1633 GND 0.02fF $ **FLOATING
C3532 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1634 GND 0.05fF $ **FLOATING
C3533 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1635 GND 0.04fF $ **FLOATING
C3534 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1636 GND 0.02fF $ **FLOATING
C3535 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1637 GND 0.03fF $ **FLOATING
C3536 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1638 GND 0.02fF $ **FLOATING
C3537 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1639 GND 0.04fF $ **FLOATING
C3538 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1640 GND 0.05fF $ **FLOATING
C3539 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1641 GND 0.02fF $ **FLOATING
C3540 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1642 GND 0.04fF $ **FLOATING
C3541 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t227 GND 0.02fF
C3542 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1643 GND 0.06fF $ **FLOATING
C3543 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1644 GND 0.05fF $ **FLOATING
C3544 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1645 GND 0.02fF $ **FLOATING
C3545 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1646 GND 0.04fF $ **FLOATING
C3546 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1647 GND 0.02fF $ **FLOATING
C3547 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1648 GND 0.05fF $ **FLOATING
C3548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1649 GND 0.02fF $ **FLOATING
C3549 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1650 GND 0.05fF $ **FLOATING
C3550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1651 GND 0.03fF $ **FLOATING
C3551 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t3 GND 0.01fF
C3552 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1652 GND 0.02fF $ **FLOATING
C3553 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.t226 GND 0.02fF
C3554 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1653 GND 0.02fF $ **FLOATING
C3555 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1654 GND 0.03fF $ **FLOATING
C3556 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB.n1655 GND 0.03fF $ **FLOATING
.end

