* SPICE3 file created from wb_flat.ext - technology: sky130A

X0 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X2 Top_1 Bot_1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X3 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X4 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X5 Top_1 Bot_1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X6 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X7 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X8 vinp1 Bot_2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X9 Top_2 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X10 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X11 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X12 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X13 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X14 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X15 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.416e+07u w=2.4e+07u
X16 Top_2 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X17 Top_2 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X18 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X19 vinp2 Bot_1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X20 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X21 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X22 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X23 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X24 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X25 Bot_1 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X26 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X27 Top_1 vbias1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X28 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X29 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X30 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X31 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X32 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X33 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X34 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X35 Top_2 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X36 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X37 Top_1 Bot_1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X38 Top_2 vbias2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X39 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X40 Top_1 Bot_1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X41 Bot_1 Bot_2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X42 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X43 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
