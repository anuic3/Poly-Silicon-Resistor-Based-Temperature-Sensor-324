* SPICE3 file created from 20bitCounter_flat.ext - technology: sky130A

X0 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41487_21# a_41474_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20327_21# a_20314_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_9681_47# a_8491_47# a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22268_47# a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_15617_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_32379_47# a_31933_47# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9747_21# a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30907_21# a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_24384_47# a_23469_47# a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_30167_47# a_29651_47# a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_19237_47# a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_805_47# a_761_289# a_639_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_38631_47# a_38115_47# a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5515_21# a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37255_21# a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_11219_47# a_10773_47# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X23 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28616_47# a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_24081_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 sky130_fd_sc_hd__dfrbp_1_0[18]/D a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_19683_47# a_19237_47# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X28 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_16095_21# a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 sky130_fd_sc_hd__dfrbp_1_0[16]/Q a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_17471_47# a_16955_47# a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X37 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3399_21# a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13979_21# a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35139_21# a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1283_21# a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 a_28791_21# a_28616_47# a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X43 a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_1108_47# a_193_47# a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X45 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11863_21# a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X46 a_15005_47# a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33023_21# a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X48 a_9572_47# a_8657_47# a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X49 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 a_1283_21# a_1108_47# a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_17121_47# a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X53 a_38281_47# a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X54 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 a_4425_47# a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X56 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7631_21# a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X57 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39371_21# a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X58 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_37255_21# a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X59 a_36165_47# a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X60 a_2309_47# a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X61 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_9269_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X62 a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X63 a_34049_47# a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X64 a_24384_47# a_23303_47# a_24037_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X65 a_41474_413# a_40397_47# a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X66 a_20314_413# a_19237_47# a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X67 a_30841_47# a_29651_47# a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X68 a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X69 a_26609_47# a_25419_47# a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X70 a_22268_47# a_21187_47# a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X71 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_11863_21# a_11797_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X72 a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X73 a_651_413# a_27_47# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_37255_21# a_37189_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X75 a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 a_28616_47# a_27535_47# a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X77 a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X78 a_35073_47# a_33883_47# a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X79 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X80 a_34617_289# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X81 a_26500_47# a_25419_47# a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X82 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_16095_21# a_16029_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X83 a_32545_47# a_32501_289# a_32379_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X84 a_13457_289# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X85 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X86 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11341_289# a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 a_38849_289# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X88 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32501_289# a_32391_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X89 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X90 a_11385_47# a_11341_289# a_11219_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X92 a_30732_47# a_29817_47# a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X93 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_4993_289# a_4883_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X95 a_26675_21# a_26500_47# a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X96 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15573_289# a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_36733_289# a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X99 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X100 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_2877_289# a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X101 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_26197_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X102 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_18211_21# a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_19587_47# a_19071_47# a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X105 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X106 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13457_289# a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X107 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X108 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34617_289# a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9225_289# a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X111 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_805_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 a_28051_47# a_27535_47# a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X115 a_3399_21# a_3224_47# a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7109_289# a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X117 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_17689_289# a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X118 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[17]/D a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X119 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_38849_289# a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X120 a_2755_47# a_2309_47# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X121 a_25585_47# a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X122 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X123 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_39371_21# a_39935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X124 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X125 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_30429_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X126 a_32391_413# a_31767_47# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_3399_21# a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X128 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X129 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_30275_413# a_29651_47# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X131 a_32957_47# a_31767_47# a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X132 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_26675_21# a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X133 a_2309_47# a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_36623_413# a_35999_47# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_13979_21# a_13913_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 a_11797_47# a_10607_47# a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X138 a_37189_47# a_35999_47# a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X139 a_34507_413# a_33883_47# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_22443_21# a_22377_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X141 a_9115_413# a_8491_47# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 a_13457_289# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X143 a_34617_289# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X144 a_20261_47# a_19071_47# a_20152_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X145 a_11341_289# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X146 a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 a_7109_289# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_32848_47# a_31933_47# a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X149 a_24037_289# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X150 a_17689_289# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X151 a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24559_21# a_24546_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_11688_47# a_10773_47# a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X154 a_15573_289# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X155 a_41421_47# a_40231_47# a_41312_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X156 a_28970_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X157 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_7631_21# a_7565_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X159 a_25935_47# a_25419_47# a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X160 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_11385_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X162 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[11]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X164 a_20152_47# a_19237_47# a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X165 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28791_21# a_28778_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 a_9225_289# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X167 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_28791_21# a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X168 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X169 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_16095_21# a_15920_47# a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_9225_289# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X173 sky130_fd_sc_hd__dfrbp_1_0[2]/Q a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26675_21# a_26662_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X175 a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X176 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 a_15451_47# a_15005_47# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X178 a_31933_47# a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X179 sky130_fd_sc_hd__dfrbp_1_0[14]/Q a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 a_7153_47# a_7109_289# a_6987_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X182 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X183 a_2659_47# a_2143_47# a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X184 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16095_21# a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X185 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 a_21703_47# a_21353_47# a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 sky130_fd_sc_hd__dfrbp_1_0[4]/Q a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X188 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_32545_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26500_47# a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X190 a_10773_47# a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 a_41312_47# a_40397_47# a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X192 a_10773_47# a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X193 a_36165_47# a_35999_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 a_40747_47# a_40397_47# a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 a_31933_47# a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X196 a_5340_47# a_4425_47# a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X197 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X198 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 a_37255_21# a_37080_47# a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X200 a_28051_47# a_27701_47# a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X201 a_6541_47# a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X202 a_15463_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_41009_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X204 a_36623_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_2767_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_19849_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X207 a_2921_47# a_2877_289# a_2755_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_36611_47# a_36165_47# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X209 a_13347_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X210 a_34507_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X211 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X212 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_15005_47# a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X214 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 a_23819_47# a_23469_47# a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X216 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18211_21# a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X217 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_1283_21# a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_9115_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 a_11231_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 a_12889_47# a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X221 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_24559_21# a_24493_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 a_22377_47# a_21187_47# a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X223 a_22430_413# a_21353_47# a_22268_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 a_6999_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 a_8657_47# a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X226 a_17579_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X227 a_38739_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X228 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_33023_21# a_32957_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 a_19237_47# a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X230 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 a_30385_289# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X232 a_26662_413# a_25585_47# a_26500_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X233 sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X234 a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X235 a_19805_289# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X236 a_40965_289# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X237 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30732_47# a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X238 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X239 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X240 a_24546_413# a_23469_47# a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_9747_21# a_9681_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X242 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_35139_21# a_35126_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 a_7565_47# a_6375_47# a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X245 a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X246 a_761_289# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X247 a_41009_47# a_40965_289# a_40843_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X248 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_33023_21# a_33010_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X249 a_22268_47# a_21353_47# a_21921_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X250 a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X251 a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X252 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_34964_47# a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X254 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X255 a_28778_413# a_27701_47# a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X256 sky130_fd_sc_hd__dfrbp_1_0[19]/Q a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11688_47# a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X258 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_32848_47# a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X259 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_21965_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X260 a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[16]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X262 a_17567_47# a_17121_47# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X263 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X264 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X265 a_15355_47# a_14839_47# a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X266 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37255_21# a_37242_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X267 a_9269_47# a_9225_289# a_9103_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X268 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41487_21# a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X269 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X270 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X271 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_12889_47# a_12723_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X273 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26675_21# a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X274 a_26031_47# a_25585_47# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X275 sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X276 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_37080_47# a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X277 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X278 a_7456_47# a_6541_47# a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X279 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X280 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X281 a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24559_21# a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X283 a_21353_47# a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X284 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_19805_289# a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_35139_21# a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X286 a_38727_47# a_38281_47# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X287 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X288 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X289 a_22443_21# a_22268_47# a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X290 a_36515_47# a_35999_47# a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X291 a_40397_47# a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X292 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22443_21# a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X293 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_13979_21# a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X294 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[7]/D a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X295 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X297 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_30907_21# a_30841_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_3224_47# a_2143_47# a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X299 a_11231_413# a_10607_47# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X300 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_2921_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 a_6541_47# a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X302 a_193_47# a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 a_4883_413# a_4259_47# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X304 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_35139_21# a_35073_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X305 a_34964_47# a_33883_47# a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X306 a_1108_47# a_27_47# a_761_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 a_7631_21# a_7456_47# a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 a_32848_47# a_31767_47# a_32501_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X309 a_32501_289# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X310 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_7153_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X311 a_15463_413# a_14839_47# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X312 a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X313 a_2767_413# a_2143_47# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X314 a_30732_47# a_29651_47# a_30385_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X315 a_11341_289# a_11123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X316 a_39196_47# a_38115_47# a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 a_18036_47# a_16955_47# a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 a_13347_413# a_12723_47# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X319 a_30907_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X320 a_5340_47# a_4259_47# a_4993_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 a_35126_413# a_34049_47# a_34964_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X322 a_19695_413# a_19071_47# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_6999_413# a_6375_47# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X324 a_37080_47# a_35999_47# a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X325 a_19805_289# a_19587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X326 a_17733_47# a_17689_289# a_17567_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X327 a_17579_413# a_16955_47# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 a_38739_413# a_38115_47# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 a_35139_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X330 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X331 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X332 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_40965_289# a_40855_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X333 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X334 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31767_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 a_30429_47# a_30385_289# a_30263_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X336 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10607_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 a_38893_47# a_38849_289# a_38727_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 a_40965_289# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X339 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X340 a_28147_47# a_27701_47# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X341 sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_26153_289# a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X343 a_11863_21# a_11688_47# a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X344 a_4993_289# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X345 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X346 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24037_289# a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X347 a_1462_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X348 a_23469_47# a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X349 a_24559_21# a_24384_47# a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X350 a_543_47# a_27_47# a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X351 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_20327_21# a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X352 a_15920_47# a_15005_47# a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X353 a_23915_47# a_23469_47# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X354 a_21703_47# a_21187_47# a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X355 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X356 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28269_289# a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X357 a_33023_21# a_32848_47# a_33202_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X358 sky130_fd_sc_hd__dfrbp_1_0[1]/Q a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_24559_21# a_25123_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[18]/D a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X361 sky130_fd_sc_hd__dfrbp_1_0[3]/Q a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[1]/D a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X363 a_8657_47# a_8491_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X364 a_25935_47# a_25585_47# a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X365 a_9747_21# a_9572_47# a_9926_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X366 sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_20327_21# a_20261_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X368 a_543_47# a_193_47# a_448_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X369 a_6891_47# a_6375_47# a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X370 a_19695_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X371 a_21921_289# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X372 a_24037_289# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X373 a_19849_47# a_19805_289# a_19683_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_41487_21# a_41421_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_26854_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X376 a_21921_289# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X377 a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[5]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X378 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_5515_21# a_5449_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 a_3333_47# a_2143_47# a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X380 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3399_21# a_3386_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X381 a_28269_289# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X382 a_448_47# sky130_fd_sc_hd__dfrbp_1_0[0]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X383 a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[2]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X384 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_28791_21# a_28725_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X385 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X386 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13979_21# a_13966_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1283_21# a_1270_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X388 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X389 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X390 a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[17]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X391 a_26153_289# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X392 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_3224_47# a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_13979_21# a_13804_47# a_14158_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 a_7109_289# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X396 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7631_21# a_7618_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 a_13335_47# a_12889_47# a_13239_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X398 a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[14]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X399 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 a_3578_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X401 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X402 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30907_21# a_30894_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[4]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X404 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9572_47# a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X405 a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[6]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X406 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_13804_47# a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X407 sky130_fd_sc_hd__dfrbp_1_0[19]/D a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X409 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_1108_47# a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X410 a_5037_47# a_4993_289# a_4871_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X411 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39371_21# a_39358_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X412 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18211_21# a_18198_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X413 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5515_21# a_5502_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X414 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[13]/D a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X415 sky130_fd_sc_hd__dfrbp_1_0[9]/Q a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20327_21# a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X417 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X419 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_7456_47# a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 a_28313_47# a_28269_289# a_28147_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X421 sky130_fd_sc_hd__dfrbp_1_0[9]/D a_20891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X422 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_16095_21# a_16082_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X423 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_38893_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X424 a_34049_47# a_33883_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X425 a_23819_47# a_23303_47# a_23724_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X426 sky130_fd_sc_hd__dfrbp_1_0[7]/Q a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X427 a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[3]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X428 a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[8]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X429 a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[18]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X430 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_39196_47# a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_18036_47# a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X432 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_5340_47# a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 a_35139_21# a_34964_47# a_35318_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X434 a_32283_47# a_31933_47# a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_9747_21# a_9734_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X436 a_34495_47# a_34049_47# a_34399_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X437 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_30907_21# a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X438 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_17733_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X440 a_26500_47# a_25585_47# a_26153_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X441 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_15920_47# a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X442 a_32283_47# a_31767_47# a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X443 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6375_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_9747_21# a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 a_30167_47# a_29817_47# a_30072_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X446 a_21353_47# a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X447 a_11123_47# a_10607_47# a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X448 a_36515_47# a_36165_47# a_36420_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X449 a_27701_47# a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X450 a_26043_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 sky130_fd_sc_hd__dfrbp_1_0[17]/Q a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X452 a_9007_47# a_8491_47# a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X453 a_34399_47# a_34049_47# a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_23927_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X455 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_28791_21# a_29355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X456 a_25585_47# a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X457 a_3224_47# a_2309_47# a_2877_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X458 a_1270_413# a_193_47# a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 a_33010_413# a_31933_47# a_32848_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X460 a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X461 a_193_47# a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X462 a_23469_47# a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X463 a_13804_47# a_12723_47# a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X464 a_30894_413# a_29817_47# a_30732_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X465 a_29817_47# a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X466 a_28159_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X467 a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X468 a_11688_47# a_10607_47# a_11341_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X469 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_18211_21# a_18145_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X470 a_5502_413# a_4425_47# a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X471 a_7631_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X472 a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X473 a_5449_47# a_4259_47# a_5340_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X474 a_7456_47# a_6375_47# a_7109_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X475 a_16082_413# a_15005_47# a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X476 a_37242_413# a_36165_47# a_37080_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X477 a_3386_413# a_2309_47# a_3224_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X478 a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X479 a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X480 a_5515_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 a_37434_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X482 a_15920_47# a_14839_47# a_15573_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X483 a_28725_47# a_27535_47# a_28616_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X484 a_16095_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 a_37255_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X486 a_16274_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X487 a_3399_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_39371_21# a_39305_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X489 a_32188_47# sky130_fd_sc_hd__dfrbp_1_0[15]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 a_7618_413# a_6541_47# a_7456_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X491 a_13239_47# a_12723_47# a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X492 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_21921_289# a_21811_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X493 a_9747_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X494 a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X495 a_36733_289# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X496 a_9572_47# a_8491_47# a_9225_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X497 a_39358_413# a_38281_47# a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X498 a_18198_413# a_17121_47# a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 a_34661_47# a_34617_289# a_34495_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X501 a_15573_289# a_15355_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X502 a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X503 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X504 sky130_fd_sc_hd__dfrbp_1_0[8]/Q a_18211_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X505 a_41487_21# a_41312_47# a_41666_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 a_13501_47# a_13457_289# a_13335_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X507 a_40843_47# a_40397_47# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X508 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_33023_21# a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X509 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_761_289# a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X510 a_34399_47# a_33883_47# a_34304_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X511 a_28616_47# a_27701_47# a_28269_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X512 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[10]/D a_23303_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X513 a_20327_21# a_20152_47# a_20506_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 sky130_fd_sc_hd__dfrbp_1_0[12]/Q a_26675_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X515 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[8]/D a_19071_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X516 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_11863_21# a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X517 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/D a_21187_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X518 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_41487_21# a_42051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X519 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_28313_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X520 a_37080_47# a_36165_47# a_36733_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X521 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X522 sky130_fd_sc_hd__dfrbp_1_0[18]/Q a_39371_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X523 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[12]/D a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X524 a_40397_47# a_40231_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X525 sky130_fd_sc_hd__dfrbp_1_0[10]/Q a_22443_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X526 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14839_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 a_21811_413# a_21187_47# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X528 a_5515_21# a_5340_47# a_5694_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X529 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_5037_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X530 a_27701_47# a_27535_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X531 a_4871_47# a_4425_47# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X532 a_40855_413# a_40231_47# a_40747_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X533 a_18145_47# a_16955_47# a_18036_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X534 a_17689_289# a_17471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X535 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_5515_21# a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 a_9103_47# a_8657_47# a_9007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X537 a_26043_413# a_25419_47# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 a_23927_413# a_23303_47# a_23819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 a_41312_47# a_40231_47# a_40965_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X540 a_20152_47# a_19071_47# a_19805_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X541 a_4425_47# a_4259_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 a_13913_47# a_12723_47# a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X543 a_39305_47# a_38115_47# a_39196_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X544 a_28159_413# a_27535_47# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X545 a_36777_47# a_36733_289# a_36611_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X546 a_25840_47# sky130_fd_sc_hd__dfrbp_1_0[12]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X547 a_18036_47# a_17121_47# a_17689_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X548 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_30385_289# a_30275_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X549 a_15617_47# a_15573_289# a_15451_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X550 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_11863_21# a_11850_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X551 a_34964_47# a_34049_47# a_34617_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X552 a_26153_289# a_25935_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X553 a_40747_47# a_40231_47# a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X554 sky130_fd_sc_hd__dfrbp_1_0[13]/Q a_28791_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X555 a_639_47# a_193_47# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X556 a_22622_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X557 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_1283_21# a_1217_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 a_24081_47# a_24037_289# a_23915_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X559 sky130_fd_sc_hd__dfrbp_1_0[4]/D a_10311_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X560 a_13804_47# a_12889_47# a_13457_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X561 sky130_fd_sc_hd__dfrbp_1_0[14]/D a_31471_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_21799_47# a_21353_47# a_21703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X563 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_34661_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X564 a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[1]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X565 a_39196_47# a_38281_47# a_38849_289# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X566 a_30907_21# a_30732_47# a_31086_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X567 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_13501_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 a_39371_21# a_39196_47# a_39550_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X569 a_30263_47# a_29817_47# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X570 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_22443_21# a_23007_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 sky130_fd_sc_hd__dfrbp_1_0[1]/D a_3963_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 sky130_fd_sc_hd__dfrbp_1_0[6]/D a_14543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 sky130_fd_sc_hd__dfrbp_1_0[11]/Q a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_2877_289# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X575 sky130_fd_sc_hd__dfrbp_1_0[16]/D a_35703_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X576 sky130_fd_sc_hd__dfrbp_1_0[0]/D a_1847_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X577 a_18211_21# a_18036_47# a_18390_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X578 a_6891_47# a_6541_47# a_6796_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X579 a_11123_47# a_10773_47# a_11028_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X580 sky130_fd_sc_hd__dfrbp_1_0[5]/D a_12427_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 sky130_fd_sc_hd__dfrbp_1_0[15]/D a_33587_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 a_7810_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X583 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X584 a_6987_47# a_6541_47# a_6891_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X585 a_17471_47# a_17121_47# a_17376_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 a_38631_47# a_38281_47# a_38536_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X587 a_29817_47# a_29651_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[11]/D a_25419_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X589 a_4775_47# a_4425_47# a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X590 a_4775_47# a_4259_47# a_4680_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X591 sky130_fd_sc_hd__dfrbp_1_0[3]/D a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X593 a_15355_47# a_15005_47# a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 a_2659_47# a_2309_47# a_2564_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X595 sky130_fd_sc_hd__dfrbp_1_0[2]/D a_6079_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_38281_47# a_38115_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_7631_21# a_8195_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X598 sky130_fd_sc_hd__dfrbp_1_0[17]/D a_37819_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 a_9007_47# a_8657_47# a_8912_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X600 a_13239_47# a_12889_47# a_13144_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X601 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[0]/CLK a_27_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X602 a_17121_47# a_16955_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[0]/D a_2143_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X604 a_11850_413# a_10773_47# a_11688_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 a_19587_47# a_19237_47# a_19492_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 a_2877_289# a_2659_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X607 a_24738_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X608 a_16029_47# a_14839_47# a_15920_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X609 a_761_289# a_543_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X610 a_32501_289# a_32283_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X611 a_21608_47# sky130_fd_sc_hd__dfrbp_1_0[10]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X612 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_26675_21# a_26609_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X613 a_24493_47# a_23303_47# a_24384_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X614 a_651_413# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X615 a_27956_47# sky130_fd_sc_hd__dfrbp_1_0[13]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X616 a_30385_289# a_30167_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X617 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_20152_47# a_20327_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X618 a_40652_47# sky130_fd_sc_hd__dfrbp_1_0[19]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X619 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_41312_47# a_41487_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X620 a_12042_47# sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X621 a_13966_413# a_12889_47# a_13804_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 a_38849_289# a_38631_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X623 a_21965_47# a_21921_289# a_21799_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_4993_289# a_4775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X625 a_9734_413# a_8657_47# a_9572_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X626 a_28269_289# a_28051_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X627 sky130_fd_sc_hd__dfrbp_1_0[8]/D a_18775_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X628 sky130_fd_sc_hd__dfrbp_1_0[0]/Q a_1283_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 a_36733_289# a_36515_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X630 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_22443_21# a_22430_413# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB a_24384_47# a_24559_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB a_3399_21# a_3333_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X633 a_15260_47# sky130_fd_sc_hd__dfrbp_1_0[7]/D sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X634 a_26197_47# a_26153_289# a_26031_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X635 a_1217_47# a_27_47# a_1108_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X636 sky130_fd_sc_hd__dfrbp_1_0[5]/Q a_11863_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B a_36777_47# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X638 sky130_fd_sc_hd__dfrbp_1_0[15]/Q a_33023_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X639 sky130_fd_sc_hd__dfrbp_1_0[6]/Q a_13979_21# sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 sky130_fd_sc_hd__dfrbp_1_0[9]/RESET_B sky130_fd_sc_hd__dfrbp_1_0[9]/VPB 8.78fF
C1 sky130_fd_sc_hd__dfrbp_1_0[9]/VPB sky130_fd_sc_hd__dfrbp_1_0[9]/VNB 69.06fF
