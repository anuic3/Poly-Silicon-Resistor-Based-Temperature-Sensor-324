magic
tech sky130A
magscale 1 2
timestamp 1634810165
<< nwell >>
rect 4886 8958 12402 8960
rect 4886 8311 12814 8958
rect 4886 8288 12836 8311
rect 4899 6905 12836 8288
rect 4900 6842 12836 6905
rect 12090 6840 12836 6842
rect 4872 1232 12844 2484
rect 12486 -3214 12948 -3212
rect 4647 -3243 5109 -3230
rect 12486 -3243 13368 -3214
rect 4647 -4008 13368 -3243
rect 4647 -4656 12518 -4008
rect 4894 -4659 12518 -4656
<< pwell >>
rect 247 8653 259 8659
rect 247 -9670 3897 8653
rect 13868 8654 13880 8660
rect 12864 -4026 12950 -4008
rect 12536 -4504 13340 -4026
rect 12536 -4526 12950 -4504
rect 12536 -4530 13380 -4526
rect 13868 -9669 17518 8654
<< nmos >>
rect 443 7150 2043 8550
rect 2101 7150 3701 8550
rect 443 5640 2043 7040
rect 2101 5640 3701 7040
rect 443 4130 2043 5530
rect 2101 4130 3701 5530
rect 443 2620 2043 4020
rect 2101 2620 3701 4020
rect 443 1110 2043 2510
rect 2101 1110 3701 2510
rect 443 -400 2043 1000
rect 2101 -400 3701 1000
rect 443 -1910 2043 -510
rect 2101 -1910 3701 -510
rect 443 -3420 2043 -2020
rect 2101 -3420 3701 -2020
rect 443 -4930 2043 -3530
rect 2101 -4930 3701 -3530
rect 443 -6440 2043 -5040
rect 2101 -6440 3701 -5040
rect 443 -7950 2043 -6550
rect 2101 -7950 3701 -6550
rect 443 -9460 2043 -8060
rect 2101 -9460 3701 -8060
rect 12732 -4320 12762 -4236
rect 13122 -4320 13152 -4236
rect 14064 7151 15664 8551
rect 15722 7151 17322 8551
rect 14064 5641 15664 7041
rect 15722 5641 17322 7041
rect 14064 4131 15664 5531
rect 15722 4131 17322 5531
rect 14064 2621 15664 4021
rect 15722 2621 17322 4021
rect 14064 1111 15664 2511
rect 15722 1111 17322 2511
rect 14064 -399 15664 1001
rect 15722 -399 17322 1001
rect 14064 -1909 15664 -509
rect 15722 -1909 17322 -509
rect 14064 -3419 15664 -2019
rect 15722 -3419 17322 -2019
rect 14064 -4929 15664 -3529
rect 15722 -4929 17322 -3529
rect 14064 -6439 15664 -5039
rect 15722 -6439 17322 -5039
rect 14064 -7949 15664 -6549
rect 15722 -7949 17322 -6549
rect 14064 -9459 15664 -8059
rect 15722 -9459 17322 -8059
<< pmos >>
rect 5412 7414 5528 7524
rect 6798 7414 6914 7524
rect 7168 7414 7284 7524
rect 7590 7414 7706 7524
rect 8012 7414 8128 7524
rect 9512 7414 9628 7524
rect 9882 7414 9998 7524
rect 10304 7414 10420 7524
rect 10726 7414 10842 7524
rect 12166 7414 12282 7524
rect 5412 1732 5528 1842
rect 6798 1731 6914 1841
rect 7168 1731 7284 1841
rect 7590 1731 7706 1841
rect 8012 1731 8128 1841
rect 9512 1735 9628 1845
rect 9882 1735 9998 1845
rect 10304 1735 10420 1845
rect 10726 1735 10842 1845
rect 12110 1732 12226 1842
rect 5457 -4192 5573 -4082
rect 6798 -4194 6914 -4084
rect 7168 -4194 7284 -4084
rect 7590 -4194 7706 -4084
rect 8012 -4194 8128 -4084
rect 9499 -4194 9615 -4084
rect 9869 -4194 9985 -4084
rect 10291 -4194 10407 -4084
rect 10713 -4194 10829 -4084
rect 12728 -3785 12758 -3449
rect 13118 -3787 13148 -3451
<< pmoslvt >>
rect 5461 8298 5661 8498
rect 6121 8298 6321 8498
rect 6591 8298 6791 8498
rect 7194 8297 7394 8497
rect 7452 8297 7652 8497
rect 7710 8297 7910 8497
rect 7968 8297 8168 8497
rect 8226 8297 8426 8497
rect 9009 8297 9209 8497
rect 9267 8297 9467 8497
rect 9525 8297 9725 8497
rect 9783 8297 9983 8497
rect 10041 8297 10241 8497
rect 10815 8297 11015 8497
rect 11073 8297 11273 8497
rect 11331 8297 11531 8497
rect 11589 8297 11789 8497
rect 11847 8297 12047 8497
rect 5765 7414 6565 7524
rect 8435 7414 9235 7524
rect 11098 7415 11898 7525
rect 5757 1732 6557 1842
rect 8434 1732 9234 1842
rect 11098 1733 11898 1843
rect 5765 -4193 6565 -4083
rect 8435 -4193 9235 -4083
rect 11098 -4192 11898 -4082
<< nmoslvt >>
rect 5187 6337 5387 6537
rect 5445 6337 5645 6537
rect 5703 6337 5903 6537
rect 5961 6337 6161 6537
rect 6219 6337 6419 6537
rect 6477 6337 6677 6537
rect 6735 6337 6935 6537
rect 6993 6337 7193 6537
rect 7857 6337 8057 6537
rect 8115 6337 8315 6537
rect 8373 6337 8573 6537
rect 8631 6337 8831 6537
rect 8889 6337 9089 6537
rect 9147 6337 9347 6537
rect 9405 6337 9605 6537
rect 9663 6337 9863 6537
rect 10520 6338 10720 6538
rect 10778 6338 10978 6538
rect 11036 6338 11236 6538
rect 11294 6338 11494 6538
rect 11552 6338 11752 6538
rect 11810 6338 12010 6538
rect 12068 6338 12268 6538
rect 12326 6338 12526 6538
rect 5187 5919 5387 6119
rect 5445 5919 5645 6119
rect 5703 5919 5903 6119
rect 5961 5919 6161 6119
rect 6219 5919 6419 6119
rect 6477 5919 6677 6119
rect 6735 5919 6935 6119
rect 6993 5919 7193 6119
rect 7857 5919 8057 6119
rect 8115 5919 8315 6119
rect 8373 5919 8573 6119
rect 8631 5919 8831 6119
rect 8889 5919 9089 6119
rect 9147 5919 9347 6119
rect 9405 5919 9605 6119
rect 9663 5919 9863 6119
rect 10520 5920 10720 6120
rect 10778 5920 10978 6120
rect 11036 5920 11236 6120
rect 11294 5920 11494 6120
rect 11552 5920 11752 6120
rect 11810 5920 12010 6120
rect 12068 5920 12268 6120
rect 12326 5920 12526 6120
rect 5187 5501 5387 5701
rect 5445 5501 5645 5701
rect 5703 5501 5903 5701
rect 5961 5501 6161 5701
rect 6219 5501 6419 5701
rect 6477 5501 6677 5701
rect 6735 5501 6935 5701
rect 6993 5501 7193 5701
rect 7857 5501 8057 5701
rect 8115 5501 8315 5701
rect 8373 5501 8573 5701
rect 8631 5501 8831 5701
rect 8889 5501 9089 5701
rect 9147 5501 9347 5701
rect 9405 5501 9605 5701
rect 9663 5501 9863 5701
rect 10520 5502 10720 5702
rect 10778 5502 10978 5702
rect 11036 5502 11236 5702
rect 11294 5502 11494 5702
rect 11552 5502 11752 5702
rect 11810 5502 12010 5702
rect 12068 5502 12268 5702
rect 12326 5502 12526 5702
rect 5187 5083 5387 5283
rect 5445 5083 5645 5283
rect 5703 5083 5903 5283
rect 5961 5083 6161 5283
rect 6219 5083 6419 5283
rect 6477 5083 6677 5283
rect 6735 5083 6935 5283
rect 6993 5083 7193 5283
rect 7857 5083 8057 5283
rect 8115 5083 8315 5283
rect 8373 5083 8573 5283
rect 8631 5083 8831 5283
rect 8889 5083 9089 5283
rect 9147 5083 9347 5283
rect 9405 5083 9605 5283
rect 9663 5083 9863 5283
rect 10520 5084 10720 5284
rect 10778 5084 10978 5284
rect 11036 5084 11236 5284
rect 11294 5084 11494 5284
rect 11552 5084 11752 5284
rect 11810 5084 12010 5284
rect 12068 5084 12268 5284
rect 12326 5084 12526 5284
rect 5187 4665 5387 4865
rect 5445 4665 5645 4865
rect 5703 4665 5903 4865
rect 5961 4665 6161 4865
rect 6219 4665 6419 4865
rect 6477 4665 6677 4865
rect 6735 4665 6935 4865
rect 6993 4665 7193 4865
rect 7857 4665 8057 4865
rect 8115 4665 8315 4865
rect 8373 4665 8573 4865
rect 8631 4665 8831 4865
rect 8889 4665 9089 4865
rect 9147 4665 9347 4865
rect 9405 4665 9605 4865
rect 9663 4665 9863 4865
rect 10520 4666 10720 4866
rect 10778 4666 10978 4866
rect 11036 4666 11236 4866
rect 11294 4666 11494 4866
rect 11552 4666 11752 4866
rect 11810 4666 12010 4866
rect 12068 4666 12268 4866
rect 12326 4666 12526 4866
rect 5187 4247 5387 4447
rect 5445 4247 5645 4447
rect 5703 4247 5903 4447
rect 5961 4247 6161 4447
rect 6219 4247 6419 4447
rect 6477 4247 6677 4447
rect 6735 4247 6935 4447
rect 6993 4247 7193 4447
rect 7857 4247 8057 4447
rect 8115 4247 8315 4447
rect 8373 4247 8573 4447
rect 8631 4247 8831 4447
rect 8889 4247 9089 4447
rect 9147 4247 9347 4447
rect 9405 4247 9605 4447
rect 9663 4247 9863 4447
rect 10520 4248 10720 4448
rect 10778 4248 10978 4448
rect 11036 4248 11236 4448
rect 11294 4248 11494 4448
rect 11552 4248 11752 4448
rect 11810 4248 12010 4448
rect 12068 4248 12268 4448
rect 12326 4248 12526 4448
rect 5187 3829 5387 4029
rect 5445 3829 5645 4029
rect 5703 3829 5903 4029
rect 5961 3829 6161 4029
rect 6219 3829 6419 4029
rect 6477 3829 6677 4029
rect 6735 3829 6935 4029
rect 6993 3829 7193 4029
rect 7857 3829 8057 4029
rect 8115 3829 8315 4029
rect 8373 3829 8573 4029
rect 8631 3829 8831 4029
rect 8889 3829 9089 4029
rect 9147 3829 9347 4029
rect 9405 3829 9605 4029
rect 9663 3829 9863 4029
rect 10520 3830 10720 4030
rect 10778 3830 10978 4030
rect 11036 3830 11236 4030
rect 11294 3830 11494 4030
rect 11552 3830 11752 4030
rect 11810 3830 12010 4030
rect 12068 3830 12268 4030
rect 12326 3830 12526 4030
rect 5067 3177 5267 3377
rect 5607 3177 5807 3377
rect 6087 3177 6287 3377
rect 6590 3179 6790 3379
rect 7100 3189 7300 3389
rect 7737 3177 7937 3377
rect 8277 3177 8477 3377
rect 8757 3177 8957 3377
rect 9260 3179 9460 3379
rect 9770 3189 9970 3389
rect 10400 3178 10600 3378
rect 10940 3178 11140 3378
rect 11420 3178 11620 3378
rect 11923 3180 12123 3380
rect 12433 3190 12633 3390
rect 5187 620 5387 820
rect 5445 620 5645 820
rect 5703 620 5903 820
rect 5961 620 6161 820
rect 6219 620 6419 820
rect 6477 620 6677 820
rect 6735 620 6935 820
rect 6993 620 7193 820
rect 7857 620 8057 820
rect 8115 620 8315 820
rect 8373 620 8573 820
rect 8631 620 8831 820
rect 8889 620 9089 820
rect 9147 620 9347 820
rect 9405 620 9605 820
rect 9663 620 9863 820
rect 10520 621 10720 821
rect 10778 621 10978 821
rect 11036 621 11236 821
rect 11294 621 11494 821
rect 11552 621 11752 821
rect 11810 621 12010 821
rect 12068 621 12268 821
rect 12326 621 12526 821
rect 5187 202 5387 402
rect 5445 202 5645 402
rect 5703 202 5903 402
rect 5961 202 6161 402
rect 6219 202 6419 402
rect 6477 202 6677 402
rect 6735 202 6935 402
rect 6993 202 7193 402
rect 7857 202 8057 402
rect 8115 202 8315 402
rect 8373 202 8573 402
rect 8631 202 8831 402
rect 8889 202 9089 402
rect 9147 202 9347 402
rect 9405 202 9605 402
rect 9663 202 9863 402
rect 10520 203 10720 403
rect 10778 203 10978 403
rect 11036 203 11236 403
rect 11294 203 11494 403
rect 11552 203 11752 403
rect 11810 203 12010 403
rect 12068 203 12268 403
rect 12326 203 12526 403
rect 5187 -216 5387 -16
rect 5445 -216 5645 -16
rect 5703 -216 5903 -16
rect 5961 -216 6161 -16
rect 6219 -216 6419 -16
rect 6477 -216 6677 -16
rect 6735 -216 6935 -16
rect 6993 -216 7193 -16
rect 7857 -216 8057 -16
rect 8115 -216 8315 -16
rect 8373 -216 8573 -16
rect 8631 -216 8831 -16
rect 8889 -216 9089 -16
rect 9147 -216 9347 -16
rect 9405 -216 9605 -16
rect 9663 -216 9863 -16
rect 10520 -215 10720 -15
rect 10778 -215 10978 -15
rect 11036 -215 11236 -15
rect 11294 -215 11494 -15
rect 11552 -215 11752 -15
rect 11810 -215 12010 -15
rect 12068 -215 12268 -15
rect 12326 -215 12526 -15
rect 5187 -634 5387 -434
rect 5445 -634 5645 -434
rect 5703 -634 5903 -434
rect 5961 -634 6161 -434
rect 6219 -634 6419 -434
rect 6477 -634 6677 -434
rect 6735 -634 6935 -434
rect 6993 -634 7193 -434
rect 7857 -634 8057 -434
rect 8115 -634 8315 -434
rect 8373 -634 8573 -434
rect 8631 -634 8831 -434
rect 8889 -634 9089 -434
rect 9147 -634 9347 -434
rect 9405 -634 9605 -434
rect 9663 -634 9863 -434
rect 10520 -633 10720 -433
rect 10778 -633 10978 -433
rect 11036 -633 11236 -433
rect 11294 -633 11494 -433
rect 11552 -633 11752 -433
rect 11810 -633 12010 -433
rect 12068 -633 12268 -433
rect 12326 -633 12526 -433
rect 5187 -1052 5387 -852
rect 5445 -1052 5645 -852
rect 5703 -1052 5903 -852
rect 5961 -1052 6161 -852
rect 6219 -1052 6419 -852
rect 6477 -1052 6677 -852
rect 6735 -1052 6935 -852
rect 6993 -1052 7193 -852
rect 7857 -1052 8057 -852
rect 8115 -1052 8315 -852
rect 8373 -1052 8573 -852
rect 8631 -1052 8831 -852
rect 8889 -1052 9089 -852
rect 9147 -1052 9347 -852
rect 9405 -1052 9605 -852
rect 9663 -1052 9863 -852
rect 10520 -1051 10720 -851
rect 10778 -1051 10978 -851
rect 11036 -1051 11236 -851
rect 11294 -1051 11494 -851
rect 11552 -1051 11752 -851
rect 11810 -1051 12010 -851
rect 12068 -1051 12268 -851
rect 12326 -1051 12526 -851
rect 5187 -1470 5387 -1270
rect 5445 -1470 5645 -1270
rect 5703 -1470 5903 -1270
rect 5961 -1470 6161 -1270
rect 6219 -1470 6419 -1270
rect 6477 -1470 6677 -1270
rect 6735 -1470 6935 -1270
rect 6993 -1470 7193 -1270
rect 7857 -1470 8057 -1270
rect 8115 -1470 8315 -1270
rect 8373 -1470 8573 -1270
rect 8631 -1470 8831 -1270
rect 8889 -1470 9089 -1270
rect 9147 -1470 9347 -1270
rect 9405 -1470 9605 -1270
rect 9663 -1470 9863 -1270
rect 10520 -1469 10720 -1269
rect 10778 -1469 10978 -1269
rect 11036 -1469 11236 -1269
rect 11294 -1469 11494 -1269
rect 11552 -1469 11752 -1269
rect 11810 -1469 12010 -1269
rect 12068 -1469 12268 -1269
rect 12326 -1469 12526 -1269
rect 5187 -1888 5387 -1688
rect 5445 -1888 5645 -1688
rect 5703 -1888 5903 -1688
rect 5961 -1888 6161 -1688
rect 6219 -1888 6419 -1688
rect 6477 -1888 6677 -1688
rect 6735 -1888 6935 -1688
rect 6993 -1888 7193 -1688
rect 7857 -1888 8057 -1688
rect 8115 -1888 8315 -1688
rect 8373 -1888 8573 -1688
rect 8631 -1888 8831 -1688
rect 8889 -1888 9089 -1688
rect 9147 -1888 9347 -1688
rect 9405 -1888 9605 -1688
rect 9663 -1888 9863 -1688
rect 10520 -1887 10720 -1687
rect 10778 -1887 10978 -1687
rect 11036 -1887 11236 -1687
rect 11294 -1887 11494 -1687
rect 11552 -1887 11752 -1687
rect 11810 -1887 12010 -1687
rect 12068 -1887 12268 -1687
rect 12326 -1887 12526 -1687
rect 5067 -2540 5267 -2340
rect 5607 -2540 5807 -2340
rect 6087 -2540 6287 -2340
rect 6590 -2538 6790 -2338
rect 7100 -2528 7300 -2328
rect 7737 -2540 7937 -2340
rect 8277 -2540 8477 -2340
rect 8757 -2540 8957 -2340
rect 9260 -2538 9460 -2338
rect 9770 -2528 9970 -2328
rect 10400 -2539 10600 -2339
rect 10940 -2539 11140 -2339
rect 11420 -2539 11620 -2339
rect 11923 -2537 12123 -2337
rect 12433 -2527 12633 -2327
rect 5187 -5284 5387 -5084
rect 5445 -5284 5645 -5084
rect 5703 -5284 5903 -5084
rect 5961 -5284 6161 -5084
rect 6219 -5284 6419 -5084
rect 6477 -5284 6677 -5084
rect 6735 -5284 6935 -5084
rect 6993 -5284 7193 -5084
rect 7857 -5284 8057 -5084
rect 8115 -5284 8315 -5084
rect 8373 -5284 8573 -5084
rect 8631 -5284 8831 -5084
rect 8889 -5284 9089 -5084
rect 9147 -5284 9347 -5084
rect 9405 -5284 9605 -5084
rect 9663 -5284 9863 -5084
rect 10520 -5283 10720 -5083
rect 10778 -5283 10978 -5083
rect 11036 -5283 11236 -5083
rect 11294 -5283 11494 -5083
rect 11552 -5283 11752 -5083
rect 11810 -5283 12010 -5083
rect 12068 -5283 12268 -5083
rect 12326 -5283 12526 -5083
rect 5187 -5702 5387 -5502
rect 5445 -5702 5645 -5502
rect 5703 -5702 5903 -5502
rect 5961 -5702 6161 -5502
rect 6219 -5702 6419 -5502
rect 6477 -5702 6677 -5502
rect 6735 -5702 6935 -5502
rect 6993 -5702 7193 -5502
rect 7857 -5702 8057 -5502
rect 8115 -5702 8315 -5502
rect 8373 -5702 8573 -5502
rect 8631 -5702 8831 -5502
rect 8889 -5702 9089 -5502
rect 9147 -5702 9347 -5502
rect 9405 -5702 9605 -5502
rect 9663 -5702 9863 -5502
rect 10520 -5701 10720 -5501
rect 10778 -5701 10978 -5501
rect 11036 -5701 11236 -5501
rect 11294 -5701 11494 -5501
rect 11552 -5701 11752 -5501
rect 11810 -5701 12010 -5501
rect 12068 -5701 12268 -5501
rect 12326 -5701 12526 -5501
rect 5187 -6120 5387 -5920
rect 5445 -6120 5645 -5920
rect 5703 -6120 5903 -5920
rect 5961 -6120 6161 -5920
rect 6219 -6120 6419 -5920
rect 6477 -6120 6677 -5920
rect 6735 -6120 6935 -5920
rect 6993 -6120 7193 -5920
rect 7857 -6120 8057 -5920
rect 8115 -6120 8315 -5920
rect 8373 -6120 8573 -5920
rect 8631 -6120 8831 -5920
rect 8889 -6120 9089 -5920
rect 9147 -6120 9347 -5920
rect 9405 -6120 9605 -5920
rect 9663 -6120 9863 -5920
rect 10520 -6119 10720 -5919
rect 10778 -6119 10978 -5919
rect 11036 -6119 11236 -5919
rect 11294 -6119 11494 -5919
rect 11552 -6119 11752 -5919
rect 11810 -6119 12010 -5919
rect 12068 -6119 12268 -5919
rect 12326 -6119 12526 -5919
rect 5187 -6538 5387 -6338
rect 5445 -6538 5645 -6338
rect 5703 -6538 5903 -6338
rect 5961 -6538 6161 -6338
rect 6219 -6538 6419 -6338
rect 6477 -6538 6677 -6338
rect 6735 -6538 6935 -6338
rect 6993 -6538 7193 -6338
rect 7857 -6538 8057 -6338
rect 8115 -6538 8315 -6338
rect 8373 -6538 8573 -6338
rect 8631 -6538 8831 -6338
rect 8889 -6538 9089 -6338
rect 9147 -6538 9347 -6338
rect 9405 -6538 9605 -6338
rect 9663 -6538 9863 -6338
rect 10520 -6537 10720 -6337
rect 10778 -6537 10978 -6337
rect 11036 -6537 11236 -6337
rect 11294 -6537 11494 -6337
rect 11552 -6537 11752 -6337
rect 11810 -6537 12010 -6337
rect 12068 -6537 12268 -6337
rect 12326 -6537 12526 -6337
rect 5187 -6956 5387 -6756
rect 5445 -6956 5645 -6756
rect 5703 -6956 5903 -6756
rect 5961 -6956 6161 -6756
rect 6219 -6956 6419 -6756
rect 6477 -6956 6677 -6756
rect 6735 -6956 6935 -6756
rect 6993 -6956 7193 -6756
rect 7857 -6956 8057 -6756
rect 8115 -6956 8315 -6756
rect 8373 -6956 8573 -6756
rect 8631 -6956 8831 -6756
rect 8889 -6956 9089 -6756
rect 9147 -6956 9347 -6756
rect 9405 -6956 9605 -6756
rect 9663 -6956 9863 -6756
rect 10520 -6955 10720 -6755
rect 10778 -6955 10978 -6755
rect 11036 -6955 11236 -6755
rect 11294 -6955 11494 -6755
rect 11552 -6955 11752 -6755
rect 11810 -6955 12010 -6755
rect 12068 -6955 12268 -6755
rect 12326 -6955 12526 -6755
rect 5187 -7374 5387 -7174
rect 5445 -7374 5645 -7174
rect 5703 -7374 5903 -7174
rect 5961 -7374 6161 -7174
rect 6219 -7374 6419 -7174
rect 6477 -7374 6677 -7174
rect 6735 -7374 6935 -7174
rect 6993 -7374 7193 -7174
rect 7857 -7374 8057 -7174
rect 8115 -7374 8315 -7174
rect 8373 -7374 8573 -7174
rect 8631 -7374 8831 -7174
rect 8889 -7374 9089 -7174
rect 9147 -7374 9347 -7174
rect 9405 -7374 9605 -7174
rect 9663 -7374 9863 -7174
rect 10520 -7373 10720 -7173
rect 10778 -7373 10978 -7173
rect 11036 -7373 11236 -7173
rect 11294 -7373 11494 -7173
rect 11552 -7373 11752 -7173
rect 11810 -7373 12010 -7173
rect 12068 -7373 12268 -7173
rect 12326 -7373 12526 -7173
rect 5187 -7792 5387 -7592
rect 5445 -7792 5645 -7592
rect 5703 -7792 5903 -7592
rect 5961 -7792 6161 -7592
rect 6219 -7792 6419 -7592
rect 6477 -7792 6677 -7592
rect 6735 -7792 6935 -7592
rect 6993 -7792 7193 -7592
rect 7857 -7792 8057 -7592
rect 8115 -7792 8315 -7592
rect 8373 -7792 8573 -7592
rect 8631 -7792 8831 -7592
rect 8889 -7792 9089 -7592
rect 9147 -7792 9347 -7592
rect 9405 -7792 9605 -7592
rect 9663 -7792 9863 -7592
rect 10520 -7791 10720 -7591
rect 10778 -7791 10978 -7591
rect 11036 -7791 11236 -7591
rect 11294 -7791 11494 -7591
rect 11552 -7791 11752 -7591
rect 11810 -7791 12010 -7591
rect 12068 -7791 12268 -7591
rect 12326 -7791 12526 -7591
rect 5067 -8444 5267 -8244
rect 5607 -8444 5807 -8244
rect 6087 -8444 6287 -8244
rect 6590 -8442 6790 -8242
rect 7100 -8432 7300 -8232
rect 7737 -8444 7937 -8244
rect 8277 -8444 8477 -8244
rect 8757 -8444 8957 -8244
rect 9260 -8442 9460 -8242
rect 9770 -8432 9970 -8232
rect 10400 -8443 10600 -8243
rect 10940 -8443 11140 -8243
rect 11420 -8443 11620 -8243
rect 11923 -8441 12123 -8241
rect 12433 -8431 12633 -8231
<< ndiff >>
rect 385 8538 443 8550
rect 385 7162 397 8538
rect 431 7162 443 8538
rect 385 7150 443 7162
rect 2043 8538 2101 8550
rect 2043 7162 2055 8538
rect 2089 7162 2101 8538
rect 2043 7150 2101 7162
rect 3701 8538 3759 8550
rect 3701 7162 3713 8538
rect 3747 7162 3759 8538
rect 3701 7150 3759 7162
rect 385 7028 443 7040
rect 385 5652 397 7028
rect 431 5652 443 7028
rect 385 5640 443 5652
rect 2043 7028 2101 7040
rect 2043 5652 2055 7028
rect 2089 5652 2101 7028
rect 2043 5640 2101 5652
rect 3701 7028 3759 7040
rect 3701 5652 3713 7028
rect 3747 5652 3759 7028
rect 3701 5640 3759 5652
rect 385 5518 443 5530
rect 385 4142 397 5518
rect 431 4142 443 5518
rect 385 4130 443 4142
rect 2043 5518 2101 5530
rect 2043 4142 2055 5518
rect 2089 4142 2101 5518
rect 2043 4130 2101 4142
rect 3701 5518 3759 5530
rect 3701 4142 3713 5518
rect 3747 4142 3759 5518
rect 3701 4130 3759 4142
rect 385 4008 443 4020
rect 385 2632 397 4008
rect 431 2632 443 4008
rect 385 2620 443 2632
rect 2043 4008 2101 4020
rect 2043 2632 2055 4008
rect 2089 2632 2101 4008
rect 2043 2620 2101 2632
rect 3701 4008 3759 4020
rect 3701 2632 3713 4008
rect 3747 2632 3759 4008
rect 3701 2620 3759 2632
rect 385 2498 443 2510
rect 385 1122 397 2498
rect 431 1122 443 2498
rect 385 1110 443 1122
rect 2043 2498 2101 2510
rect 2043 1122 2055 2498
rect 2089 1122 2101 2498
rect 2043 1110 2101 1122
rect 3701 2498 3759 2510
rect 3701 1122 3713 2498
rect 3747 1122 3759 2498
rect 3701 1110 3759 1122
rect 385 988 443 1000
rect 385 -388 397 988
rect 431 -388 443 988
rect 385 -400 443 -388
rect 2043 988 2101 1000
rect 2043 -388 2055 988
rect 2089 -388 2101 988
rect 2043 -400 2101 -388
rect 3701 988 3759 1000
rect 3701 -388 3713 988
rect 3747 -388 3759 988
rect 3701 -400 3759 -388
rect 385 -522 443 -510
rect 385 -1898 397 -522
rect 431 -1898 443 -522
rect 385 -1910 443 -1898
rect 2043 -522 2101 -510
rect 2043 -1898 2055 -522
rect 2089 -1898 2101 -522
rect 2043 -1910 2101 -1898
rect 3701 -522 3759 -510
rect 3701 -1898 3713 -522
rect 3747 -1898 3759 -522
rect 3701 -1910 3759 -1898
rect 385 -2032 443 -2020
rect 385 -3408 397 -2032
rect 431 -3408 443 -2032
rect 385 -3420 443 -3408
rect 2043 -2032 2101 -2020
rect 2043 -3408 2055 -2032
rect 2089 -3408 2101 -2032
rect 2043 -3420 2101 -3408
rect 3701 -2032 3759 -2020
rect 3701 -3408 3713 -2032
rect 3747 -3408 3759 -2032
rect 3701 -3420 3759 -3408
rect 385 -3542 443 -3530
rect 385 -4918 397 -3542
rect 431 -4918 443 -3542
rect 385 -4930 443 -4918
rect 2043 -3542 2101 -3530
rect 2043 -4918 2055 -3542
rect 2089 -4918 2101 -3542
rect 2043 -4930 2101 -4918
rect 3701 -3542 3759 -3530
rect 3701 -4918 3713 -3542
rect 3747 -4918 3759 -3542
rect 3701 -4930 3759 -4918
rect 385 -5052 443 -5040
rect 385 -6428 397 -5052
rect 431 -6428 443 -5052
rect 385 -6440 443 -6428
rect 2043 -5052 2101 -5040
rect 2043 -6428 2055 -5052
rect 2089 -6428 2101 -5052
rect 2043 -6440 2101 -6428
rect 3701 -5052 3759 -5040
rect 3701 -6428 3713 -5052
rect 3747 -6428 3759 -5052
rect 3701 -6440 3759 -6428
rect 385 -6562 443 -6550
rect 385 -7938 397 -6562
rect 431 -7938 443 -6562
rect 385 -7950 443 -7938
rect 2043 -6562 2101 -6550
rect 2043 -7938 2055 -6562
rect 2089 -7938 2101 -6562
rect 2043 -7950 2101 -7938
rect 3701 -6562 3759 -6550
rect 3701 -7938 3713 -6562
rect 3747 -7938 3759 -6562
rect 3701 -7950 3759 -7938
rect 385 -8072 443 -8060
rect 385 -9448 397 -8072
rect 431 -9448 443 -8072
rect 385 -9460 443 -9448
rect 2043 -8072 2101 -8060
rect 2043 -9448 2055 -8072
rect 2089 -9448 2101 -8072
rect 2043 -9460 2101 -9448
rect 3701 -8072 3759 -8060
rect 3701 -9448 3713 -8072
rect 3747 -9448 3759 -8072
rect 3701 -9460 3759 -9448
rect 5129 6525 5187 6537
rect 5129 6489 5141 6525
rect 5175 6489 5187 6525
rect 5129 6455 5187 6489
rect 5129 6419 5141 6455
rect 5175 6419 5187 6455
rect 5129 6385 5187 6419
rect 5129 6349 5141 6385
rect 5175 6349 5187 6385
rect 5129 6337 5187 6349
rect 5387 6525 5445 6537
rect 5387 6489 5399 6525
rect 5433 6489 5445 6525
rect 5387 6455 5445 6489
rect 5387 6419 5399 6455
rect 5433 6419 5445 6455
rect 5387 6385 5445 6419
rect 5387 6349 5399 6385
rect 5433 6349 5445 6385
rect 5387 6337 5445 6349
rect 5645 6525 5703 6537
rect 5645 6489 5657 6525
rect 5691 6489 5703 6525
rect 5645 6455 5703 6489
rect 5645 6419 5657 6455
rect 5691 6419 5703 6455
rect 5645 6384 5703 6419
rect 5645 6348 5657 6384
rect 5691 6348 5703 6384
rect 5645 6337 5703 6348
rect 5903 6525 5961 6537
rect 5903 6489 5915 6525
rect 5949 6489 5961 6525
rect 5903 6455 5961 6489
rect 5903 6419 5915 6455
rect 5949 6419 5961 6455
rect 5903 6385 5961 6419
rect 5903 6349 5915 6385
rect 5949 6349 5961 6385
rect 5903 6337 5961 6349
rect 6161 6525 6219 6537
rect 6161 6489 6173 6525
rect 6207 6489 6219 6525
rect 6161 6455 6219 6489
rect 6161 6419 6173 6455
rect 6207 6419 6219 6455
rect 6161 6385 6219 6419
rect 6161 6349 6173 6385
rect 6207 6349 6219 6385
rect 6161 6337 6219 6349
rect 6419 6525 6477 6537
rect 6419 6489 6431 6525
rect 6465 6489 6477 6525
rect 6419 6455 6477 6489
rect 6419 6419 6431 6455
rect 6465 6419 6477 6455
rect 6419 6385 6477 6419
rect 6419 6349 6431 6385
rect 6465 6349 6477 6385
rect 6419 6337 6477 6349
rect 6677 6525 6735 6537
rect 6677 6489 6689 6525
rect 6723 6489 6735 6525
rect 6677 6455 6735 6489
rect 6677 6419 6689 6455
rect 6723 6419 6735 6455
rect 6677 6385 6735 6419
rect 6677 6349 6689 6385
rect 6723 6349 6735 6385
rect 6677 6337 6735 6349
rect 6935 6525 6993 6537
rect 6935 6489 6947 6525
rect 6981 6489 6993 6525
rect 6935 6455 6993 6489
rect 6935 6419 6947 6455
rect 6981 6419 6993 6455
rect 6935 6385 6993 6419
rect 6935 6349 6947 6385
rect 6981 6349 6993 6385
rect 6935 6337 6993 6349
rect 7193 6525 7251 6537
rect 7193 6489 7205 6525
rect 7239 6489 7251 6525
rect 7193 6455 7251 6489
rect 7193 6419 7205 6455
rect 7239 6419 7251 6455
rect 7193 6385 7251 6419
rect 7193 6349 7205 6385
rect 7239 6349 7251 6385
rect 7193 6337 7251 6349
rect 7799 6525 7857 6537
rect 7799 6489 7811 6525
rect 7845 6489 7857 6525
rect 7799 6455 7857 6489
rect 7799 6419 7811 6455
rect 7845 6419 7857 6455
rect 7799 6385 7857 6419
rect 7799 6349 7811 6385
rect 7845 6349 7857 6385
rect 7799 6337 7857 6349
rect 8057 6525 8115 6537
rect 8057 6489 8069 6525
rect 8103 6489 8115 6525
rect 8057 6455 8115 6489
rect 8057 6419 8069 6455
rect 8103 6419 8115 6455
rect 8057 6385 8115 6419
rect 8057 6349 8069 6385
rect 8103 6349 8115 6385
rect 8057 6337 8115 6349
rect 8315 6525 8373 6537
rect 8315 6489 8327 6525
rect 8361 6489 8373 6525
rect 8315 6455 8373 6489
rect 8315 6419 8327 6455
rect 8361 6419 8373 6455
rect 8315 6384 8373 6419
rect 8315 6348 8327 6384
rect 8361 6348 8373 6384
rect 8315 6337 8373 6348
rect 8573 6525 8631 6537
rect 8573 6489 8585 6525
rect 8619 6489 8631 6525
rect 8573 6455 8631 6489
rect 8573 6419 8585 6455
rect 8619 6419 8631 6455
rect 8573 6385 8631 6419
rect 8573 6349 8585 6385
rect 8619 6349 8631 6385
rect 8573 6337 8631 6349
rect 8831 6525 8889 6537
rect 8831 6489 8843 6525
rect 8877 6489 8889 6525
rect 8831 6455 8889 6489
rect 8831 6419 8843 6455
rect 8877 6419 8889 6455
rect 8831 6385 8889 6419
rect 8831 6349 8843 6385
rect 8877 6349 8889 6385
rect 8831 6337 8889 6349
rect 9089 6525 9147 6537
rect 9089 6489 9101 6525
rect 9135 6489 9147 6525
rect 9089 6455 9147 6489
rect 9089 6419 9101 6455
rect 9135 6419 9147 6455
rect 9089 6385 9147 6419
rect 9089 6349 9101 6385
rect 9135 6349 9147 6385
rect 9089 6337 9147 6349
rect 9347 6525 9405 6537
rect 9347 6489 9359 6525
rect 9393 6489 9405 6525
rect 9347 6455 9405 6489
rect 9347 6419 9359 6455
rect 9393 6419 9405 6455
rect 9347 6385 9405 6419
rect 9347 6349 9359 6385
rect 9393 6349 9405 6385
rect 9347 6337 9405 6349
rect 9605 6525 9663 6537
rect 9605 6489 9617 6525
rect 9651 6489 9663 6525
rect 9605 6455 9663 6489
rect 9605 6419 9617 6455
rect 9651 6419 9663 6455
rect 9605 6385 9663 6419
rect 9605 6349 9617 6385
rect 9651 6349 9663 6385
rect 9605 6337 9663 6349
rect 9863 6525 9921 6537
rect 9863 6489 9875 6525
rect 9909 6489 9921 6525
rect 9863 6455 9921 6489
rect 9863 6419 9875 6455
rect 9909 6419 9921 6455
rect 9863 6385 9921 6419
rect 9863 6349 9875 6385
rect 9909 6349 9921 6385
rect 9863 6337 9921 6349
rect 10462 6526 10520 6538
rect 10462 6490 10474 6526
rect 10508 6490 10520 6526
rect 10462 6456 10520 6490
rect 10462 6420 10474 6456
rect 10508 6420 10520 6456
rect 10462 6386 10520 6420
rect 10462 6350 10474 6386
rect 10508 6350 10520 6386
rect 10462 6338 10520 6350
rect 10720 6526 10778 6538
rect 10720 6490 10732 6526
rect 10766 6490 10778 6526
rect 10720 6456 10778 6490
rect 10720 6420 10732 6456
rect 10766 6420 10778 6456
rect 10720 6386 10778 6420
rect 10720 6350 10732 6386
rect 10766 6350 10778 6386
rect 10720 6338 10778 6350
rect 10978 6526 11036 6538
rect 10978 6490 10990 6526
rect 11024 6490 11036 6526
rect 10978 6456 11036 6490
rect 10978 6420 10990 6456
rect 11024 6420 11036 6456
rect 10978 6385 11036 6420
rect 10978 6349 10990 6385
rect 11024 6349 11036 6385
rect 10978 6338 11036 6349
rect 11236 6526 11294 6538
rect 11236 6490 11248 6526
rect 11282 6490 11294 6526
rect 11236 6456 11294 6490
rect 11236 6420 11248 6456
rect 11282 6420 11294 6456
rect 11236 6386 11294 6420
rect 11236 6350 11248 6386
rect 11282 6350 11294 6386
rect 11236 6338 11294 6350
rect 11494 6526 11552 6538
rect 11494 6490 11506 6526
rect 11540 6490 11552 6526
rect 11494 6456 11552 6490
rect 11494 6420 11506 6456
rect 11540 6420 11552 6456
rect 11494 6386 11552 6420
rect 11494 6350 11506 6386
rect 11540 6350 11552 6386
rect 11494 6338 11552 6350
rect 11752 6526 11810 6538
rect 11752 6490 11764 6526
rect 11798 6490 11810 6526
rect 11752 6456 11810 6490
rect 11752 6420 11764 6456
rect 11798 6420 11810 6456
rect 11752 6386 11810 6420
rect 11752 6350 11764 6386
rect 11798 6350 11810 6386
rect 11752 6338 11810 6350
rect 12010 6526 12068 6538
rect 12010 6490 12022 6526
rect 12056 6490 12068 6526
rect 12010 6456 12068 6490
rect 12010 6420 12022 6456
rect 12056 6420 12068 6456
rect 12010 6386 12068 6420
rect 12010 6350 12022 6386
rect 12056 6350 12068 6386
rect 12010 6338 12068 6350
rect 12268 6526 12326 6538
rect 12268 6490 12280 6526
rect 12314 6490 12326 6526
rect 12268 6456 12326 6490
rect 12268 6420 12280 6456
rect 12314 6420 12326 6456
rect 12268 6386 12326 6420
rect 12268 6350 12280 6386
rect 12314 6350 12326 6386
rect 12268 6338 12326 6350
rect 12526 6526 12584 6538
rect 12526 6490 12538 6526
rect 12572 6490 12584 6526
rect 12526 6456 12584 6490
rect 12526 6420 12538 6456
rect 12572 6420 12584 6456
rect 12526 6386 12584 6420
rect 12526 6350 12538 6386
rect 12572 6350 12584 6386
rect 12526 6338 12584 6350
rect 5129 6107 5187 6119
rect 5129 6071 5141 6107
rect 5175 6071 5187 6107
rect 5129 6037 5187 6071
rect 5129 6001 5141 6037
rect 5175 6001 5187 6037
rect 5129 5967 5187 6001
rect 5129 5931 5141 5967
rect 5175 5931 5187 5967
rect 5129 5919 5187 5931
rect 5387 6107 5445 6119
rect 5387 6071 5399 6107
rect 5433 6071 5445 6107
rect 5387 6037 5445 6071
rect 5387 6001 5399 6037
rect 5433 6001 5445 6037
rect 5387 5967 5445 6001
rect 5387 5931 5399 5967
rect 5433 5931 5445 5967
rect 5387 5919 5445 5931
rect 5645 6107 5703 6119
rect 5645 6071 5657 6107
rect 5691 6071 5703 6107
rect 5645 6037 5703 6071
rect 5645 6001 5657 6037
rect 5691 6001 5703 6037
rect 5645 5966 5703 6001
rect 5645 5930 5657 5966
rect 5691 5930 5703 5966
rect 5645 5919 5703 5930
rect 5903 6107 5961 6119
rect 5903 6071 5915 6107
rect 5949 6071 5961 6107
rect 5903 6037 5961 6071
rect 5903 6001 5915 6037
rect 5949 6001 5961 6037
rect 5903 5967 5961 6001
rect 5903 5931 5915 5967
rect 5949 5931 5961 5967
rect 5903 5919 5961 5931
rect 6161 6107 6219 6119
rect 6161 6071 6173 6107
rect 6207 6071 6219 6107
rect 6161 6037 6219 6071
rect 6161 6001 6173 6037
rect 6207 6001 6219 6037
rect 6161 5967 6219 6001
rect 6161 5931 6173 5967
rect 6207 5931 6219 5967
rect 6161 5919 6219 5931
rect 6419 6107 6477 6119
rect 6419 6071 6431 6107
rect 6465 6071 6477 6107
rect 6419 6037 6477 6071
rect 6419 6001 6431 6037
rect 6465 6001 6477 6037
rect 6419 5967 6477 6001
rect 6419 5931 6431 5967
rect 6465 5931 6477 5967
rect 6419 5919 6477 5931
rect 6677 6107 6735 6119
rect 6677 6071 6689 6107
rect 6723 6071 6735 6107
rect 6677 6037 6735 6071
rect 6677 6001 6689 6037
rect 6723 6001 6735 6037
rect 6677 5967 6735 6001
rect 6677 5931 6689 5967
rect 6723 5931 6735 5967
rect 6677 5919 6735 5931
rect 6935 6107 6993 6119
rect 6935 6071 6947 6107
rect 6981 6071 6993 6107
rect 6935 6037 6993 6071
rect 6935 6001 6947 6037
rect 6981 6001 6993 6037
rect 6935 5967 6993 6001
rect 6935 5931 6947 5967
rect 6981 5931 6993 5967
rect 6935 5919 6993 5931
rect 7193 6107 7251 6119
rect 7193 6071 7205 6107
rect 7239 6071 7251 6107
rect 7193 6037 7251 6071
rect 7193 6001 7205 6037
rect 7239 6001 7251 6037
rect 7193 5967 7251 6001
rect 7193 5931 7205 5967
rect 7239 5931 7251 5967
rect 7193 5919 7251 5931
rect 7799 6107 7857 6119
rect 7799 6071 7811 6107
rect 7845 6071 7857 6107
rect 7799 6037 7857 6071
rect 7799 6001 7811 6037
rect 7845 6001 7857 6037
rect 7799 5967 7857 6001
rect 7799 5931 7811 5967
rect 7845 5931 7857 5967
rect 7799 5919 7857 5931
rect 8057 6107 8115 6119
rect 8057 6071 8069 6107
rect 8103 6071 8115 6107
rect 8057 6037 8115 6071
rect 8057 6001 8069 6037
rect 8103 6001 8115 6037
rect 8057 5967 8115 6001
rect 8057 5931 8069 5967
rect 8103 5931 8115 5967
rect 8057 5919 8115 5931
rect 8315 6107 8373 6119
rect 8315 6071 8327 6107
rect 8361 6071 8373 6107
rect 8315 6037 8373 6071
rect 8315 6001 8327 6037
rect 8361 6001 8373 6037
rect 8315 5966 8373 6001
rect 8315 5930 8327 5966
rect 8361 5930 8373 5966
rect 8315 5919 8373 5930
rect 8573 6107 8631 6119
rect 8573 6071 8585 6107
rect 8619 6071 8631 6107
rect 8573 6037 8631 6071
rect 8573 6001 8585 6037
rect 8619 6001 8631 6037
rect 8573 5967 8631 6001
rect 8573 5931 8585 5967
rect 8619 5931 8631 5967
rect 8573 5919 8631 5931
rect 8831 6107 8889 6119
rect 8831 6071 8843 6107
rect 8877 6071 8889 6107
rect 8831 6037 8889 6071
rect 8831 6001 8843 6037
rect 8877 6001 8889 6037
rect 8831 5967 8889 6001
rect 8831 5931 8843 5967
rect 8877 5931 8889 5967
rect 8831 5919 8889 5931
rect 9089 6107 9147 6119
rect 9089 6071 9101 6107
rect 9135 6071 9147 6107
rect 9089 6037 9147 6071
rect 9089 6001 9101 6037
rect 9135 6001 9147 6037
rect 9089 5967 9147 6001
rect 9089 5931 9101 5967
rect 9135 5931 9147 5967
rect 9089 5919 9147 5931
rect 9347 6107 9405 6119
rect 9347 6071 9359 6107
rect 9393 6071 9405 6107
rect 9347 6037 9405 6071
rect 9347 6001 9359 6037
rect 9393 6001 9405 6037
rect 9347 5967 9405 6001
rect 9347 5931 9359 5967
rect 9393 5931 9405 5967
rect 9347 5919 9405 5931
rect 9605 6107 9663 6119
rect 9605 6071 9617 6107
rect 9651 6071 9663 6107
rect 9605 6037 9663 6071
rect 9605 6001 9617 6037
rect 9651 6001 9663 6037
rect 9605 5967 9663 6001
rect 9605 5931 9617 5967
rect 9651 5931 9663 5967
rect 9605 5919 9663 5931
rect 9863 6107 9921 6119
rect 9863 6071 9875 6107
rect 9909 6071 9921 6107
rect 9863 6037 9921 6071
rect 9863 6001 9875 6037
rect 9909 6001 9921 6037
rect 9863 5967 9921 6001
rect 9863 5931 9875 5967
rect 9909 5931 9921 5967
rect 9863 5919 9921 5931
rect 10462 6108 10520 6120
rect 10462 6072 10474 6108
rect 10508 6072 10520 6108
rect 10462 6038 10520 6072
rect 10462 6002 10474 6038
rect 10508 6002 10520 6038
rect 10462 5968 10520 6002
rect 10462 5932 10474 5968
rect 10508 5932 10520 5968
rect 10462 5920 10520 5932
rect 10720 6108 10778 6120
rect 10720 6072 10732 6108
rect 10766 6072 10778 6108
rect 10720 6038 10778 6072
rect 10720 6002 10732 6038
rect 10766 6002 10778 6038
rect 10720 5968 10778 6002
rect 10720 5932 10732 5968
rect 10766 5932 10778 5968
rect 10720 5920 10778 5932
rect 10978 6108 11036 6120
rect 10978 6072 10990 6108
rect 11024 6072 11036 6108
rect 10978 6038 11036 6072
rect 10978 6002 10990 6038
rect 11024 6002 11036 6038
rect 10978 5967 11036 6002
rect 10978 5931 10990 5967
rect 11024 5931 11036 5967
rect 10978 5920 11036 5931
rect 11236 6108 11294 6120
rect 11236 6072 11248 6108
rect 11282 6072 11294 6108
rect 11236 6038 11294 6072
rect 11236 6002 11248 6038
rect 11282 6002 11294 6038
rect 11236 5968 11294 6002
rect 11236 5932 11248 5968
rect 11282 5932 11294 5968
rect 11236 5920 11294 5932
rect 11494 6108 11552 6120
rect 11494 6072 11506 6108
rect 11540 6072 11552 6108
rect 11494 6038 11552 6072
rect 11494 6002 11506 6038
rect 11540 6002 11552 6038
rect 11494 5968 11552 6002
rect 11494 5932 11506 5968
rect 11540 5932 11552 5968
rect 11494 5920 11552 5932
rect 11752 6108 11810 6120
rect 11752 6072 11764 6108
rect 11798 6072 11810 6108
rect 11752 6038 11810 6072
rect 11752 6002 11764 6038
rect 11798 6002 11810 6038
rect 11752 5968 11810 6002
rect 11752 5932 11764 5968
rect 11798 5932 11810 5968
rect 11752 5920 11810 5932
rect 12010 6108 12068 6120
rect 12010 6072 12022 6108
rect 12056 6072 12068 6108
rect 12010 6038 12068 6072
rect 12010 6002 12022 6038
rect 12056 6002 12068 6038
rect 12010 5968 12068 6002
rect 12010 5932 12022 5968
rect 12056 5932 12068 5968
rect 12010 5920 12068 5932
rect 12268 6108 12326 6120
rect 12268 6072 12280 6108
rect 12314 6072 12326 6108
rect 12268 6038 12326 6072
rect 12268 6002 12280 6038
rect 12314 6002 12326 6038
rect 12268 5968 12326 6002
rect 12268 5932 12280 5968
rect 12314 5932 12326 5968
rect 12268 5920 12326 5932
rect 12526 6108 12584 6120
rect 12526 6072 12538 6108
rect 12572 6072 12584 6108
rect 12526 6038 12584 6072
rect 12526 6002 12538 6038
rect 12572 6002 12584 6038
rect 12526 5968 12584 6002
rect 12526 5932 12538 5968
rect 12572 5932 12584 5968
rect 12526 5920 12584 5932
rect 5129 5689 5187 5701
rect 5129 5653 5141 5689
rect 5175 5653 5187 5689
rect 5129 5619 5187 5653
rect 5129 5583 5141 5619
rect 5175 5583 5187 5619
rect 5129 5549 5187 5583
rect 5129 5513 5141 5549
rect 5175 5513 5187 5549
rect 5129 5501 5187 5513
rect 5387 5689 5445 5701
rect 5387 5653 5399 5689
rect 5433 5653 5445 5689
rect 5387 5619 5445 5653
rect 5387 5583 5399 5619
rect 5433 5583 5445 5619
rect 5387 5549 5445 5583
rect 5387 5513 5399 5549
rect 5433 5513 5445 5549
rect 5387 5501 5445 5513
rect 5645 5689 5703 5701
rect 5645 5653 5657 5689
rect 5691 5653 5703 5689
rect 5645 5619 5703 5653
rect 5645 5583 5657 5619
rect 5691 5583 5703 5619
rect 5645 5548 5703 5583
rect 5645 5512 5657 5548
rect 5691 5512 5703 5548
rect 5645 5501 5703 5512
rect 5903 5689 5961 5701
rect 5903 5653 5915 5689
rect 5949 5653 5961 5689
rect 5903 5619 5961 5653
rect 5903 5583 5915 5619
rect 5949 5583 5961 5619
rect 5903 5549 5961 5583
rect 5903 5513 5915 5549
rect 5949 5513 5961 5549
rect 5903 5501 5961 5513
rect 6161 5689 6219 5701
rect 6161 5653 6173 5689
rect 6207 5653 6219 5689
rect 6161 5619 6219 5653
rect 6161 5583 6173 5619
rect 6207 5583 6219 5619
rect 6161 5549 6219 5583
rect 6161 5513 6173 5549
rect 6207 5513 6219 5549
rect 6161 5501 6219 5513
rect 6419 5689 6477 5701
rect 6419 5653 6431 5689
rect 6465 5653 6477 5689
rect 6419 5619 6477 5653
rect 6419 5583 6431 5619
rect 6465 5583 6477 5619
rect 6419 5549 6477 5583
rect 6419 5513 6431 5549
rect 6465 5513 6477 5549
rect 6419 5501 6477 5513
rect 6677 5689 6735 5701
rect 6677 5653 6689 5689
rect 6723 5653 6735 5689
rect 6677 5619 6735 5653
rect 6677 5583 6689 5619
rect 6723 5583 6735 5619
rect 6677 5549 6735 5583
rect 6677 5513 6689 5549
rect 6723 5513 6735 5549
rect 6677 5501 6735 5513
rect 6935 5689 6993 5701
rect 6935 5653 6947 5689
rect 6981 5653 6993 5689
rect 6935 5619 6993 5653
rect 6935 5583 6947 5619
rect 6981 5583 6993 5619
rect 6935 5549 6993 5583
rect 6935 5513 6947 5549
rect 6981 5513 6993 5549
rect 6935 5501 6993 5513
rect 7193 5689 7251 5701
rect 7193 5653 7205 5689
rect 7239 5653 7251 5689
rect 7193 5619 7251 5653
rect 7193 5583 7205 5619
rect 7239 5583 7251 5619
rect 7193 5549 7251 5583
rect 7193 5513 7205 5549
rect 7239 5513 7251 5549
rect 7193 5501 7251 5513
rect 7799 5689 7857 5701
rect 7799 5653 7811 5689
rect 7845 5653 7857 5689
rect 7799 5619 7857 5653
rect 7799 5583 7811 5619
rect 7845 5583 7857 5619
rect 7799 5549 7857 5583
rect 7799 5513 7811 5549
rect 7845 5513 7857 5549
rect 7799 5501 7857 5513
rect 8057 5689 8115 5701
rect 8057 5653 8069 5689
rect 8103 5653 8115 5689
rect 8057 5619 8115 5653
rect 8057 5583 8069 5619
rect 8103 5583 8115 5619
rect 8057 5549 8115 5583
rect 8057 5513 8069 5549
rect 8103 5513 8115 5549
rect 8057 5501 8115 5513
rect 8315 5689 8373 5701
rect 8315 5653 8327 5689
rect 8361 5653 8373 5689
rect 8315 5619 8373 5653
rect 8315 5583 8327 5619
rect 8361 5583 8373 5619
rect 8315 5548 8373 5583
rect 8315 5512 8327 5548
rect 8361 5512 8373 5548
rect 8315 5501 8373 5512
rect 8573 5689 8631 5701
rect 8573 5653 8585 5689
rect 8619 5653 8631 5689
rect 8573 5619 8631 5653
rect 8573 5583 8585 5619
rect 8619 5583 8631 5619
rect 8573 5549 8631 5583
rect 8573 5513 8585 5549
rect 8619 5513 8631 5549
rect 8573 5501 8631 5513
rect 8831 5689 8889 5701
rect 8831 5653 8843 5689
rect 8877 5653 8889 5689
rect 8831 5619 8889 5653
rect 8831 5583 8843 5619
rect 8877 5583 8889 5619
rect 8831 5549 8889 5583
rect 8831 5513 8843 5549
rect 8877 5513 8889 5549
rect 8831 5501 8889 5513
rect 9089 5689 9147 5701
rect 9089 5653 9101 5689
rect 9135 5653 9147 5689
rect 9089 5619 9147 5653
rect 9089 5583 9101 5619
rect 9135 5583 9147 5619
rect 9089 5549 9147 5583
rect 9089 5513 9101 5549
rect 9135 5513 9147 5549
rect 9089 5501 9147 5513
rect 9347 5689 9405 5701
rect 9347 5653 9359 5689
rect 9393 5653 9405 5689
rect 9347 5619 9405 5653
rect 9347 5583 9359 5619
rect 9393 5583 9405 5619
rect 9347 5549 9405 5583
rect 9347 5513 9359 5549
rect 9393 5513 9405 5549
rect 9347 5501 9405 5513
rect 9605 5689 9663 5701
rect 9605 5653 9617 5689
rect 9651 5653 9663 5689
rect 9605 5619 9663 5653
rect 9605 5583 9617 5619
rect 9651 5583 9663 5619
rect 9605 5549 9663 5583
rect 9605 5513 9617 5549
rect 9651 5513 9663 5549
rect 9605 5501 9663 5513
rect 9863 5689 9921 5701
rect 9863 5653 9875 5689
rect 9909 5653 9921 5689
rect 9863 5619 9921 5653
rect 9863 5583 9875 5619
rect 9909 5583 9921 5619
rect 9863 5549 9921 5583
rect 9863 5513 9875 5549
rect 9909 5513 9921 5549
rect 9863 5501 9921 5513
rect 10462 5690 10520 5702
rect 10462 5654 10474 5690
rect 10508 5654 10520 5690
rect 10462 5620 10520 5654
rect 10462 5584 10474 5620
rect 10508 5584 10520 5620
rect 10462 5550 10520 5584
rect 10462 5514 10474 5550
rect 10508 5514 10520 5550
rect 10462 5502 10520 5514
rect 10720 5690 10778 5702
rect 10720 5654 10732 5690
rect 10766 5654 10778 5690
rect 10720 5620 10778 5654
rect 10720 5584 10732 5620
rect 10766 5584 10778 5620
rect 10720 5550 10778 5584
rect 10720 5514 10732 5550
rect 10766 5514 10778 5550
rect 10720 5502 10778 5514
rect 10978 5690 11036 5702
rect 10978 5654 10990 5690
rect 11024 5654 11036 5690
rect 10978 5620 11036 5654
rect 10978 5584 10990 5620
rect 11024 5584 11036 5620
rect 10978 5549 11036 5584
rect 10978 5513 10990 5549
rect 11024 5513 11036 5549
rect 10978 5502 11036 5513
rect 11236 5690 11294 5702
rect 11236 5654 11248 5690
rect 11282 5654 11294 5690
rect 11236 5620 11294 5654
rect 11236 5584 11248 5620
rect 11282 5584 11294 5620
rect 11236 5550 11294 5584
rect 11236 5514 11248 5550
rect 11282 5514 11294 5550
rect 11236 5502 11294 5514
rect 11494 5690 11552 5702
rect 11494 5654 11506 5690
rect 11540 5654 11552 5690
rect 11494 5620 11552 5654
rect 11494 5584 11506 5620
rect 11540 5584 11552 5620
rect 11494 5550 11552 5584
rect 11494 5514 11506 5550
rect 11540 5514 11552 5550
rect 11494 5502 11552 5514
rect 11752 5690 11810 5702
rect 11752 5654 11764 5690
rect 11798 5654 11810 5690
rect 11752 5620 11810 5654
rect 11752 5584 11764 5620
rect 11798 5584 11810 5620
rect 11752 5550 11810 5584
rect 11752 5514 11764 5550
rect 11798 5514 11810 5550
rect 11752 5502 11810 5514
rect 12010 5690 12068 5702
rect 12010 5654 12022 5690
rect 12056 5654 12068 5690
rect 12010 5620 12068 5654
rect 12010 5584 12022 5620
rect 12056 5584 12068 5620
rect 12010 5550 12068 5584
rect 12010 5514 12022 5550
rect 12056 5514 12068 5550
rect 12010 5502 12068 5514
rect 12268 5690 12326 5702
rect 12268 5654 12280 5690
rect 12314 5654 12326 5690
rect 12268 5620 12326 5654
rect 12268 5584 12280 5620
rect 12314 5584 12326 5620
rect 12268 5550 12326 5584
rect 12268 5514 12280 5550
rect 12314 5514 12326 5550
rect 12268 5502 12326 5514
rect 12526 5690 12584 5702
rect 12526 5654 12538 5690
rect 12572 5654 12584 5690
rect 12526 5620 12584 5654
rect 12526 5584 12538 5620
rect 12572 5584 12584 5620
rect 12526 5550 12584 5584
rect 12526 5514 12538 5550
rect 12572 5514 12584 5550
rect 12526 5502 12584 5514
rect 5129 5271 5187 5283
rect 5129 5235 5141 5271
rect 5175 5235 5187 5271
rect 5129 5201 5187 5235
rect 5129 5165 5141 5201
rect 5175 5165 5187 5201
rect 5129 5131 5187 5165
rect 5129 5095 5141 5131
rect 5175 5095 5187 5131
rect 5129 5083 5187 5095
rect 5387 5271 5445 5283
rect 5387 5235 5399 5271
rect 5433 5235 5445 5271
rect 5387 5201 5445 5235
rect 5387 5165 5399 5201
rect 5433 5165 5445 5201
rect 5387 5131 5445 5165
rect 5387 5095 5399 5131
rect 5433 5095 5445 5131
rect 5387 5083 5445 5095
rect 5645 5271 5703 5283
rect 5645 5235 5657 5271
rect 5691 5235 5703 5271
rect 5645 5201 5703 5235
rect 5645 5165 5657 5201
rect 5691 5165 5703 5201
rect 5645 5130 5703 5165
rect 5645 5094 5657 5130
rect 5691 5094 5703 5130
rect 5645 5083 5703 5094
rect 5903 5271 5961 5283
rect 5903 5235 5915 5271
rect 5949 5235 5961 5271
rect 5903 5201 5961 5235
rect 5903 5165 5915 5201
rect 5949 5165 5961 5201
rect 5903 5131 5961 5165
rect 5903 5095 5915 5131
rect 5949 5095 5961 5131
rect 5903 5083 5961 5095
rect 6161 5271 6219 5283
rect 6161 5235 6173 5271
rect 6207 5235 6219 5271
rect 6161 5201 6219 5235
rect 6161 5165 6173 5201
rect 6207 5165 6219 5201
rect 6161 5131 6219 5165
rect 6161 5095 6173 5131
rect 6207 5095 6219 5131
rect 6161 5083 6219 5095
rect 6419 5271 6477 5283
rect 6419 5235 6431 5271
rect 6465 5235 6477 5271
rect 6419 5201 6477 5235
rect 6419 5165 6431 5201
rect 6465 5165 6477 5201
rect 6419 5131 6477 5165
rect 6419 5095 6431 5131
rect 6465 5095 6477 5131
rect 6419 5083 6477 5095
rect 6677 5271 6735 5283
rect 6677 5235 6689 5271
rect 6723 5235 6735 5271
rect 6677 5201 6735 5235
rect 6677 5165 6689 5201
rect 6723 5165 6735 5201
rect 6677 5131 6735 5165
rect 6677 5095 6689 5131
rect 6723 5095 6735 5131
rect 6677 5083 6735 5095
rect 6935 5271 6993 5283
rect 6935 5235 6947 5271
rect 6981 5235 6993 5271
rect 6935 5201 6993 5235
rect 6935 5165 6947 5201
rect 6981 5165 6993 5201
rect 6935 5131 6993 5165
rect 6935 5095 6947 5131
rect 6981 5095 6993 5131
rect 6935 5083 6993 5095
rect 7193 5271 7251 5283
rect 7193 5235 7205 5271
rect 7239 5235 7251 5271
rect 7193 5201 7251 5235
rect 7193 5165 7205 5201
rect 7239 5165 7251 5201
rect 7193 5131 7251 5165
rect 7193 5095 7205 5131
rect 7239 5095 7251 5131
rect 7193 5083 7251 5095
rect 7799 5271 7857 5283
rect 7799 5235 7811 5271
rect 7845 5235 7857 5271
rect 7799 5201 7857 5235
rect 7799 5165 7811 5201
rect 7845 5165 7857 5201
rect 7799 5131 7857 5165
rect 7799 5095 7811 5131
rect 7845 5095 7857 5131
rect 7799 5083 7857 5095
rect 8057 5271 8115 5283
rect 8057 5235 8069 5271
rect 8103 5235 8115 5271
rect 8057 5201 8115 5235
rect 8057 5165 8069 5201
rect 8103 5165 8115 5201
rect 8057 5131 8115 5165
rect 8057 5095 8069 5131
rect 8103 5095 8115 5131
rect 8057 5083 8115 5095
rect 8315 5271 8373 5283
rect 8315 5235 8327 5271
rect 8361 5235 8373 5271
rect 8315 5201 8373 5235
rect 8315 5165 8327 5201
rect 8361 5165 8373 5201
rect 8315 5130 8373 5165
rect 8315 5094 8327 5130
rect 8361 5094 8373 5130
rect 8315 5083 8373 5094
rect 8573 5271 8631 5283
rect 8573 5235 8585 5271
rect 8619 5235 8631 5271
rect 8573 5201 8631 5235
rect 8573 5165 8585 5201
rect 8619 5165 8631 5201
rect 8573 5131 8631 5165
rect 8573 5095 8585 5131
rect 8619 5095 8631 5131
rect 8573 5083 8631 5095
rect 8831 5271 8889 5283
rect 8831 5235 8843 5271
rect 8877 5235 8889 5271
rect 8831 5201 8889 5235
rect 8831 5165 8843 5201
rect 8877 5165 8889 5201
rect 8831 5131 8889 5165
rect 8831 5095 8843 5131
rect 8877 5095 8889 5131
rect 8831 5083 8889 5095
rect 9089 5271 9147 5283
rect 9089 5235 9101 5271
rect 9135 5235 9147 5271
rect 9089 5201 9147 5235
rect 9089 5165 9101 5201
rect 9135 5165 9147 5201
rect 9089 5131 9147 5165
rect 9089 5095 9101 5131
rect 9135 5095 9147 5131
rect 9089 5083 9147 5095
rect 9347 5271 9405 5283
rect 9347 5235 9359 5271
rect 9393 5235 9405 5271
rect 9347 5201 9405 5235
rect 9347 5165 9359 5201
rect 9393 5165 9405 5201
rect 9347 5131 9405 5165
rect 9347 5095 9359 5131
rect 9393 5095 9405 5131
rect 9347 5083 9405 5095
rect 9605 5271 9663 5283
rect 9605 5235 9617 5271
rect 9651 5235 9663 5271
rect 9605 5201 9663 5235
rect 9605 5165 9617 5201
rect 9651 5165 9663 5201
rect 9605 5131 9663 5165
rect 9605 5095 9617 5131
rect 9651 5095 9663 5131
rect 9605 5083 9663 5095
rect 9863 5271 9921 5283
rect 9863 5235 9875 5271
rect 9909 5235 9921 5271
rect 9863 5201 9921 5235
rect 9863 5165 9875 5201
rect 9909 5165 9921 5201
rect 9863 5131 9921 5165
rect 9863 5095 9875 5131
rect 9909 5095 9921 5131
rect 9863 5083 9921 5095
rect 10462 5272 10520 5284
rect 10462 5236 10474 5272
rect 10508 5236 10520 5272
rect 10462 5202 10520 5236
rect 10462 5166 10474 5202
rect 10508 5166 10520 5202
rect 10462 5132 10520 5166
rect 10462 5096 10474 5132
rect 10508 5096 10520 5132
rect 10462 5084 10520 5096
rect 10720 5272 10778 5284
rect 10720 5236 10732 5272
rect 10766 5236 10778 5272
rect 10720 5202 10778 5236
rect 10720 5166 10732 5202
rect 10766 5166 10778 5202
rect 10720 5132 10778 5166
rect 10720 5096 10732 5132
rect 10766 5096 10778 5132
rect 10720 5084 10778 5096
rect 10978 5272 11036 5284
rect 10978 5236 10990 5272
rect 11024 5236 11036 5272
rect 10978 5202 11036 5236
rect 10978 5166 10990 5202
rect 11024 5166 11036 5202
rect 10978 5131 11036 5166
rect 10978 5095 10990 5131
rect 11024 5095 11036 5131
rect 10978 5084 11036 5095
rect 11236 5272 11294 5284
rect 11236 5236 11248 5272
rect 11282 5236 11294 5272
rect 11236 5202 11294 5236
rect 11236 5166 11248 5202
rect 11282 5166 11294 5202
rect 11236 5132 11294 5166
rect 11236 5096 11248 5132
rect 11282 5096 11294 5132
rect 11236 5084 11294 5096
rect 11494 5272 11552 5284
rect 11494 5236 11506 5272
rect 11540 5236 11552 5272
rect 11494 5202 11552 5236
rect 11494 5166 11506 5202
rect 11540 5166 11552 5202
rect 11494 5132 11552 5166
rect 11494 5096 11506 5132
rect 11540 5096 11552 5132
rect 11494 5084 11552 5096
rect 11752 5272 11810 5284
rect 11752 5236 11764 5272
rect 11798 5236 11810 5272
rect 11752 5202 11810 5236
rect 11752 5166 11764 5202
rect 11798 5166 11810 5202
rect 11752 5132 11810 5166
rect 11752 5096 11764 5132
rect 11798 5096 11810 5132
rect 11752 5084 11810 5096
rect 12010 5272 12068 5284
rect 12010 5236 12022 5272
rect 12056 5236 12068 5272
rect 12010 5202 12068 5236
rect 12010 5166 12022 5202
rect 12056 5166 12068 5202
rect 12010 5132 12068 5166
rect 12010 5096 12022 5132
rect 12056 5096 12068 5132
rect 12010 5084 12068 5096
rect 12268 5272 12326 5284
rect 12268 5236 12280 5272
rect 12314 5236 12326 5272
rect 12268 5202 12326 5236
rect 12268 5166 12280 5202
rect 12314 5166 12326 5202
rect 12268 5132 12326 5166
rect 12268 5096 12280 5132
rect 12314 5096 12326 5132
rect 12268 5084 12326 5096
rect 12526 5272 12584 5284
rect 12526 5236 12538 5272
rect 12572 5236 12584 5272
rect 12526 5202 12584 5236
rect 12526 5166 12538 5202
rect 12572 5166 12584 5202
rect 12526 5132 12584 5166
rect 12526 5096 12538 5132
rect 12572 5096 12584 5132
rect 12526 5084 12584 5096
rect 5129 4853 5187 4865
rect 5129 4817 5141 4853
rect 5175 4817 5187 4853
rect 5129 4783 5187 4817
rect 5129 4747 5141 4783
rect 5175 4747 5187 4783
rect 5129 4713 5187 4747
rect 5129 4677 5141 4713
rect 5175 4677 5187 4713
rect 5129 4665 5187 4677
rect 5387 4853 5445 4865
rect 5387 4817 5399 4853
rect 5433 4817 5445 4853
rect 5387 4783 5445 4817
rect 5387 4747 5399 4783
rect 5433 4747 5445 4783
rect 5387 4713 5445 4747
rect 5387 4677 5399 4713
rect 5433 4677 5445 4713
rect 5387 4665 5445 4677
rect 5645 4853 5703 4865
rect 5645 4817 5657 4853
rect 5691 4817 5703 4853
rect 5645 4783 5703 4817
rect 5645 4747 5657 4783
rect 5691 4747 5703 4783
rect 5645 4712 5703 4747
rect 5645 4676 5657 4712
rect 5691 4676 5703 4712
rect 5645 4665 5703 4676
rect 5903 4853 5961 4865
rect 5903 4817 5915 4853
rect 5949 4817 5961 4853
rect 5903 4783 5961 4817
rect 5903 4747 5915 4783
rect 5949 4747 5961 4783
rect 5903 4713 5961 4747
rect 5903 4677 5915 4713
rect 5949 4677 5961 4713
rect 5903 4665 5961 4677
rect 6161 4853 6219 4865
rect 6161 4817 6173 4853
rect 6207 4817 6219 4853
rect 6161 4783 6219 4817
rect 6161 4747 6173 4783
rect 6207 4747 6219 4783
rect 6161 4713 6219 4747
rect 6161 4677 6173 4713
rect 6207 4677 6219 4713
rect 6161 4665 6219 4677
rect 6419 4853 6477 4865
rect 6419 4817 6431 4853
rect 6465 4817 6477 4853
rect 6419 4783 6477 4817
rect 6419 4747 6431 4783
rect 6465 4747 6477 4783
rect 6419 4713 6477 4747
rect 6419 4677 6431 4713
rect 6465 4677 6477 4713
rect 6419 4665 6477 4677
rect 6677 4853 6735 4865
rect 6677 4817 6689 4853
rect 6723 4817 6735 4853
rect 6677 4783 6735 4817
rect 6677 4747 6689 4783
rect 6723 4747 6735 4783
rect 6677 4713 6735 4747
rect 6677 4677 6689 4713
rect 6723 4677 6735 4713
rect 6677 4665 6735 4677
rect 6935 4853 6993 4865
rect 6935 4817 6947 4853
rect 6981 4817 6993 4853
rect 6935 4783 6993 4817
rect 6935 4747 6947 4783
rect 6981 4747 6993 4783
rect 6935 4713 6993 4747
rect 6935 4677 6947 4713
rect 6981 4677 6993 4713
rect 6935 4665 6993 4677
rect 7193 4853 7251 4865
rect 7193 4817 7205 4853
rect 7239 4817 7251 4853
rect 7193 4783 7251 4817
rect 7193 4747 7205 4783
rect 7239 4747 7251 4783
rect 7193 4713 7251 4747
rect 7193 4677 7205 4713
rect 7239 4677 7251 4713
rect 7193 4665 7251 4677
rect 7799 4853 7857 4865
rect 7799 4817 7811 4853
rect 7845 4817 7857 4853
rect 7799 4783 7857 4817
rect 7799 4747 7811 4783
rect 7845 4747 7857 4783
rect 7799 4713 7857 4747
rect 7799 4677 7811 4713
rect 7845 4677 7857 4713
rect 7799 4665 7857 4677
rect 8057 4853 8115 4865
rect 8057 4817 8069 4853
rect 8103 4817 8115 4853
rect 8057 4783 8115 4817
rect 8057 4747 8069 4783
rect 8103 4747 8115 4783
rect 8057 4713 8115 4747
rect 8057 4677 8069 4713
rect 8103 4677 8115 4713
rect 8057 4665 8115 4677
rect 8315 4853 8373 4865
rect 8315 4817 8327 4853
rect 8361 4817 8373 4853
rect 8315 4783 8373 4817
rect 8315 4747 8327 4783
rect 8361 4747 8373 4783
rect 8315 4712 8373 4747
rect 8315 4676 8327 4712
rect 8361 4676 8373 4712
rect 8315 4665 8373 4676
rect 8573 4853 8631 4865
rect 8573 4817 8585 4853
rect 8619 4817 8631 4853
rect 8573 4783 8631 4817
rect 8573 4747 8585 4783
rect 8619 4747 8631 4783
rect 8573 4713 8631 4747
rect 8573 4677 8585 4713
rect 8619 4677 8631 4713
rect 8573 4665 8631 4677
rect 8831 4853 8889 4865
rect 8831 4817 8843 4853
rect 8877 4817 8889 4853
rect 8831 4783 8889 4817
rect 8831 4747 8843 4783
rect 8877 4747 8889 4783
rect 8831 4713 8889 4747
rect 8831 4677 8843 4713
rect 8877 4677 8889 4713
rect 8831 4665 8889 4677
rect 9089 4853 9147 4865
rect 9089 4817 9101 4853
rect 9135 4817 9147 4853
rect 9089 4783 9147 4817
rect 9089 4747 9101 4783
rect 9135 4747 9147 4783
rect 9089 4713 9147 4747
rect 9089 4677 9101 4713
rect 9135 4677 9147 4713
rect 9089 4665 9147 4677
rect 9347 4853 9405 4865
rect 9347 4817 9359 4853
rect 9393 4817 9405 4853
rect 9347 4783 9405 4817
rect 9347 4747 9359 4783
rect 9393 4747 9405 4783
rect 9347 4713 9405 4747
rect 9347 4677 9359 4713
rect 9393 4677 9405 4713
rect 9347 4665 9405 4677
rect 9605 4853 9663 4865
rect 9605 4817 9617 4853
rect 9651 4817 9663 4853
rect 9605 4783 9663 4817
rect 9605 4747 9617 4783
rect 9651 4747 9663 4783
rect 9605 4713 9663 4747
rect 9605 4677 9617 4713
rect 9651 4677 9663 4713
rect 9605 4665 9663 4677
rect 9863 4853 9921 4865
rect 9863 4817 9875 4853
rect 9909 4817 9921 4853
rect 9863 4783 9921 4817
rect 9863 4747 9875 4783
rect 9909 4747 9921 4783
rect 9863 4713 9921 4747
rect 9863 4677 9875 4713
rect 9909 4677 9921 4713
rect 9863 4665 9921 4677
rect 10462 4854 10520 4866
rect 10462 4818 10474 4854
rect 10508 4818 10520 4854
rect 10462 4784 10520 4818
rect 10462 4748 10474 4784
rect 10508 4748 10520 4784
rect 10462 4714 10520 4748
rect 10462 4678 10474 4714
rect 10508 4678 10520 4714
rect 10462 4666 10520 4678
rect 10720 4854 10778 4866
rect 10720 4818 10732 4854
rect 10766 4818 10778 4854
rect 10720 4784 10778 4818
rect 10720 4748 10732 4784
rect 10766 4748 10778 4784
rect 10720 4714 10778 4748
rect 10720 4678 10732 4714
rect 10766 4678 10778 4714
rect 10720 4666 10778 4678
rect 10978 4854 11036 4866
rect 10978 4818 10990 4854
rect 11024 4818 11036 4854
rect 10978 4784 11036 4818
rect 10978 4748 10990 4784
rect 11024 4748 11036 4784
rect 10978 4713 11036 4748
rect 10978 4677 10990 4713
rect 11024 4677 11036 4713
rect 10978 4666 11036 4677
rect 11236 4854 11294 4866
rect 11236 4818 11248 4854
rect 11282 4818 11294 4854
rect 11236 4784 11294 4818
rect 11236 4748 11248 4784
rect 11282 4748 11294 4784
rect 11236 4714 11294 4748
rect 11236 4678 11248 4714
rect 11282 4678 11294 4714
rect 11236 4666 11294 4678
rect 11494 4854 11552 4866
rect 11494 4818 11506 4854
rect 11540 4818 11552 4854
rect 11494 4784 11552 4818
rect 11494 4748 11506 4784
rect 11540 4748 11552 4784
rect 11494 4714 11552 4748
rect 11494 4678 11506 4714
rect 11540 4678 11552 4714
rect 11494 4666 11552 4678
rect 11752 4854 11810 4866
rect 11752 4818 11764 4854
rect 11798 4818 11810 4854
rect 11752 4784 11810 4818
rect 11752 4748 11764 4784
rect 11798 4748 11810 4784
rect 11752 4714 11810 4748
rect 11752 4678 11764 4714
rect 11798 4678 11810 4714
rect 11752 4666 11810 4678
rect 12010 4854 12068 4866
rect 12010 4818 12022 4854
rect 12056 4818 12068 4854
rect 12010 4784 12068 4818
rect 12010 4748 12022 4784
rect 12056 4748 12068 4784
rect 12010 4714 12068 4748
rect 12010 4678 12022 4714
rect 12056 4678 12068 4714
rect 12010 4666 12068 4678
rect 12268 4854 12326 4866
rect 12268 4818 12280 4854
rect 12314 4818 12326 4854
rect 12268 4784 12326 4818
rect 12268 4748 12280 4784
rect 12314 4748 12326 4784
rect 12268 4714 12326 4748
rect 12268 4678 12280 4714
rect 12314 4678 12326 4714
rect 12268 4666 12326 4678
rect 12526 4854 12584 4866
rect 12526 4818 12538 4854
rect 12572 4818 12584 4854
rect 12526 4784 12584 4818
rect 12526 4748 12538 4784
rect 12572 4748 12584 4784
rect 12526 4714 12584 4748
rect 12526 4678 12538 4714
rect 12572 4678 12584 4714
rect 12526 4666 12584 4678
rect 5129 4435 5187 4447
rect 5129 4399 5141 4435
rect 5175 4399 5187 4435
rect 5129 4365 5187 4399
rect 5129 4329 5141 4365
rect 5175 4329 5187 4365
rect 5129 4295 5187 4329
rect 5129 4259 5141 4295
rect 5175 4259 5187 4295
rect 5129 4247 5187 4259
rect 5387 4435 5445 4447
rect 5387 4399 5399 4435
rect 5433 4399 5445 4435
rect 5387 4365 5445 4399
rect 5387 4329 5399 4365
rect 5433 4329 5445 4365
rect 5387 4295 5445 4329
rect 5387 4259 5399 4295
rect 5433 4259 5445 4295
rect 5387 4247 5445 4259
rect 5645 4435 5703 4447
rect 5645 4399 5657 4435
rect 5691 4399 5703 4435
rect 5645 4365 5703 4399
rect 5645 4329 5657 4365
rect 5691 4329 5703 4365
rect 5645 4294 5703 4329
rect 5645 4258 5657 4294
rect 5691 4258 5703 4294
rect 5645 4247 5703 4258
rect 5903 4435 5961 4447
rect 5903 4399 5915 4435
rect 5949 4399 5961 4435
rect 5903 4365 5961 4399
rect 5903 4329 5915 4365
rect 5949 4329 5961 4365
rect 5903 4295 5961 4329
rect 5903 4259 5915 4295
rect 5949 4259 5961 4295
rect 5903 4247 5961 4259
rect 6161 4435 6219 4447
rect 6161 4399 6173 4435
rect 6207 4399 6219 4435
rect 6161 4365 6219 4399
rect 6161 4329 6173 4365
rect 6207 4329 6219 4365
rect 6161 4295 6219 4329
rect 6161 4259 6173 4295
rect 6207 4259 6219 4295
rect 6161 4247 6219 4259
rect 6419 4435 6477 4447
rect 6419 4399 6431 4435
rect 6465 4399 6477 4435
rect 6419 4365 6477 4399
rect 6419 4329 6431 4365
rect 6465 4329 6477 4365
rect 6419 4295 6477 4329
rect 6419 4259 6431 4295
rect 6465 4259 6477 4295
rect 6419 4247 6477 4259
rect 6677 4435 6735 4447
rect 6677 4399 6689 4435
rect 6723 4399 6735 4435
rect 6677 4365 6735 4399
rect 6677 4329 6689 4365
rect 6723 4329 6735 4365
rect 6677 4295 6735 4329
rect 6677 4259 6689 4295
rect 6723 4259 6735 4295
rect 6677 4247 6735 4259
rect 6935 4435 6993 4447
rect 6935 4399 6947 4435
rect 6981 4399 6993 4435
rect 6935 4365 6993 4399
rect 6935 4329 6947 4365
rect 6981 4329 6993 4365
rect 6935 4295 6993 4329
rect 6935 4259 6947 4295
rect 6981 4259 6993 4295
rect 6935 4247 6993 4259
rect 7193 4435 7251 4447
rect 7193 4399 7205 4435
rect 7239 4399 7251 4435
rect 7193 4365 7251 4399
rect 7193 4329 7205 4365
rect 7239 4329 7251 4365
rect 7193 4295 7251 4329
rect 7193 4259 7205 4295
rect 7239 4259 7251 4295
rect 7193 4247 7251 4259
rect 7799 4435 7857 4447
rect 7799 4399 7811 4435
rect 7845 4399 7857 4435
rect 7799 4365 7857 4399
rect 7799 4329 7811 4365
rect 7845 4329 7857 4365
rect 7799 4295 7857 4329
rect 7799 4259 7811 4295
rect 7845 4259 7857 4295
rect 7799 4247 7857 4259
rect 8057 4435 8115 4447
rect 8057 4399 8069 4435
rect 8103 4399 8115 4435
rect 8057 4365 8115 4399
rect 8057 4329 8069 4365
rect 8103 4329 8115 4365
rect 8057 4295 8115 4329
rect 8057 4259 8069 4295
rect 8103 4259 8115 4295
rect 8057 4247 8115 4259
rect 8315 4435 8373 4447
rect 8315 4399 8327 4435
rect 8361 4399 8373 4435
rect 8315 4365 8373 4399
rect 8315 4329 8327 4365
rect 8361 4329 8373 4365
rect 8315 4294 8373 4329
rect 8315 4258 8327 4294
rect 8361 4258 8373 4294
rect 8315 4247 8373 4258
rect 8573 4435 8631 4447
rect 8573 4399 8585 4435
rect 8619 4399 8631 4435
rect 8573 4365 8631 4399
rect 8573 4329 8585 4365
rect 8619 4329 8631 4365
rect 8573 4295 8631 4329
rect 8573 4259 8585 4295
rect 8619 4259 8631 4295
rect 8573 4247 8631 4259
rect 8831 4435 8889 4447
rect 8831 4399 8843 4435
rect 8877 4399 8889 4435
rect 8831 4365 8889 4399
rect 8831 4329 8843 4365
rect 8877 4329 8889 4365
rect 8831 4295 8889 4329
rect 8831 4259 8843 4295
rect 8877 4259 8889 4295
rect 8831 4247 8889 4259
rect 9089 4435 9147 4447
rect 9089 4399 9101 4435
rect 9135 4399 9147 4435
rect 9089 4365 9147 4399
rect 9089 4329 9101 4365
rect 9135 4329 9147 4365
rect 9089 4295 9147 4329
rect 9089 4259 9101 4295
rect 9135 4259 9147 4295
rect 9089 4247 9147 4259
rect 9347 4435 9405 4447
rect 9347 4399 9359 4435
rect 9393 4399 9405 4435
rect 9347 4365 9405 4399
rect 9347 4329 9359 4365
rect 9393 4329 9405 4365
rect 9347 4295 9405 4329
rect 9347 4259 9359 4295
rect 9393 4259 9405 4295
rect 9347 4247 9405 4259
rect 9605 4435 9663 4447
rect 9605 4399 9617 4435
rect 9651 4399 9663 4435
rect 9605 4365 9663 4399
rect 9605 4329 9617 4365
rect 9651 4329 9663 4365
rect 9605 4295 9663 4329
rect 9605 4259 9617 4295
rect 9651 4259 9663 4295
rect 9605 4247 9663 4259
rect 9863 4435 9921 4447
rect 9863 4399 9875 4435
rect 9909 4399 9921 4435
rect 9863 4365 9921 4399
rect 9863 4329 9875 4365
rect 9909 4329 9921 4365
rect 9863 4295 9921 4329
rect 9863 4259 9875 4295
rect 9909 4259 9921 4295
rect 9863 4247 9921 4259
rect 10462 4436 10520 4448
rect 10462 4400 10474 4436
rect 10508 4400 10520 4436
rect 10462 4366 10520 4400
rect 10462 4330 10474 4366
rect 10508 4330 10520 4366
rect 10462 4296 10520 4330
rect 10462 4260 10474 4296
rect 10508 4260 10520 4296
rect 10462 4248 10520 4260
rect 10720 4436 10778 4448
rect 10720 4400 10732 4436
rect 10766 4400 10778 4436
rect 10720 4366 10778 4400
rect 10720 4330 10732 4366
rect 10766 4330 10778 4366
rect 10720 4296 10778 4330
rect 10720 4260 10732 4296
rect 10766 4260 10778 4296
rect 10720 4248 10778 4260
rect 10978 4436 11036 4448
rect 10978 4400 10990 4436
rect 11024 4400 11036 4436
rect 10978 4366 11036 4400
rect 10978 4330 10990 4366
rect 11024 4330 11036 4366
rect 10978 4295 11036 4330
rect 10978 4259 10990 4295
rect 11024 4259 11036 4295
rect 10978 4248 11036 4259
rect 11236 4436 11294 4448
rect 11236 4400 11248 4436
rect 11282 4400 11294 4436
rect 11236 4366 11294 4400
rect 11236 4330 11248 4366
rect 11282 4330 11294 4366
rect 11236 4296 11294 4330
rect 11236 4260 11248 4296
rect 11282 4260 11294 4296
rect 11236 4248 11294 4260
rect 11494 4436 11552 4448
rect 11494 4400 11506 4436
rect 11540 4400 11552 4436
rect 11494 4366 11552 4400
rect 11494 4330 11506 4366
rect 11540 4330 11552 4366
rect 11494 4296 11552 4330
rect 11494 4260 11506 4296
rect 11540 4260 11552 4296
rect 11494 4248 11552 4260
rect 11752 4436 11810 4448
rect 11752 4400 11764 4436
rect 11798 4400 11810 4436
rect 11752 4366 11810 4400
rect 11752 4330 11764 4366
rect 11798 4330 11810 4366
rect 11752 4296 11810 4330
rect 11752 4260 11764 4296
rect 11798 4260 11810 4296
rect 11752 4248 11810 4260
rect 12010 4436 12068 4448
rect 12010 4400 12022 4436
rect 12056 4400 12068 4436
rect 12010 4366 12068 4400
rect 12010 4330 12022 4366
rect 12056 4330 12068 4366
rect 12010 4296 12068 4330
rect 12010 4260 12022 4296
rect 12056 4260 12068 4296
rect 12010 4248 12068 4260
rect 12268 4436 12326 4448
rect 12268 4400 12280 4436
rect 12314 4400 12326 4436
rect 12268 4366 12326 4400
rect 12268 4330 12280 4366
rect 12314 4330 12326 4366
rect 12268 4296 12326 4330
rect 12268 4260 12280 4296
rect 12314 4260 12326 4296
rect 12268 4248 12326 4260
rect 12526 4436 12584 4448
rect 12526 4400 12538 4436
rect 12572 4400 12584 4436
rect 12526 4366 12584 4400
rect 12526 4330 12538 4366
rect 12572 4330 12584 4366
rect 12526 4296 12584 4330
rect 12526 4260 12538 4296
rect 12572 4260 12584 4296
rect 12526 4248 12584 4260
rect 5129 4017 5187 4029
rect 5129 3981 5141 4017
rect 5175 3981 5187 4017
rect 5129 3947 5187 3981
rect 5129 3911 5141 3947
rect 5175 3911 5187 3947
rect 5129 3877 5187 3911
rect 5129 3841 5141 3877
rect 5175 3841 5187 3877
rect 5129 3829 5187 3841
rect 5387 4017 5445 4029
rect 5387 3981 5399 4017
rect 5433 3981 5445 4017
rect 5387 3947 5445 3981
rect 5387 3911 5399 3947
rect 5433 3911 5445 3947
rect 5387 3877 5445 3911
rect 5387 3841 5399 3877
rect 5433 3841 5445 3877
rect 5387 3829 5445 3841
rect 5645 4017 5703 4029
rect 5645 3981 5657 4017
rect 5691 3981 5703 4017
rect 5645 3947 5703 3981
rect 5645 3911 5657 3947
rect 5691 3911 5703 3947
rect 5645 3876 5703 3911
rect 5645 3840 5657 3876
rect 5691 3840 5703 3876
rect 5645 3829 5703 3840
rect 5903 4017 5961 4029
rect 5903 3981 5915 4017
rect 5949 3981 5961 4017
rect 5903 3947 5961 3981
rect 5903 3911 5915 3947
rect 5949 3911 5961 3947
rect 5903 3877 5961 3911
rect 5903 3841 5915 3877
rect 5949 3841 5961 3877
rect 5903 3829 5961 3841
rect 6161 4017 6219 4029
rect 6161 3981 6173 4017
rect 6207 3981 6219 4017
rect 6161 3947 6219 3981
rect 6161 3911 6173 3947
rect 6207 3911 6219 3947
rect 6161 3877 6219 3911
rect 6161 3841 6173 3877
rect 6207 3841 6219 3877
rect 6161 3829 6219 3841
rect 6419 4017 6477 4029
rect 6419 3981 6431 4017
rect 6465 3981 6477 4017
rect 6419 3947 6477 3981
rect 6419 3911 6431 3947
rect 6465 3911 6477 3947
rect 6419 3877 6477 3911
rect 6419 3841 6431 3877
rect 6465 3841 6477 3877
rect 6419 3829 6477 3841
rect 6677 4017 6735 4029
rect 6677 3981 6689 4017
rect 6723 3981 6735 4017
rect 6677 3947 6735 3981
rect 6677 3911 6689 3947
rect 6723 3911 6735 3947
rect 6677 3877 6735 3911
rect 6677 3841 6689 3877
rect 6723 3841 6735 3877
rect 6677 3829 6735 3841
rect 6935 4017 6993 4029
rect 6935 3981 6947 4017
rect 6981 3981 6993 4017
rect 6935 3947 6993 3981
rect 6935 3911 6947 3947
rect 6981 3911 6993 3947
rect 6935 3877 6993 3911
rect 6935 3841 6947 3877
rect 6981 3841 6993 3877
rect 6935 3829 6993 3841
rect 7193 4017 7251 4029
rect 7193 3981 7205 4017
rect 7239 3981 7251 4017
rect 7193 3947 7251 3981
rect 7193 3911 7205 3947
rect 7239 3911 7251 3947
rect 7193 3877 7251 3911
rect 7193 3841 7205 3877
rect 7239 3841 7251 3877
rect 7193 3829 7251 3841
rect 7799 4017 7857 4029
rect 7799 3981 7811 4017
rect 7845 3981 7857 4017
rect 7799 3947 7857 3981
rect 7799 3911 7811 3947
rect 7845 3911 7857 3947
rect 7799 3877 7857 3911
rect 7799 3841 7811 3877
rect 7845 3841 7857 3877
rect 7799 3829 7857 3841
rect 8057 4017 8115 4029
rect 8057 3981 8069 4017
rect 8103 3981 8115 4017
rect 8057 3947 8115 3981
rect 8057 3911 8069 3947
rect 8103 3911 8115 3947
rect 8057 3877 8115 3911
rect 8057 3841 8069 3877
rect 8103 3841 8115 3877
rect 8057 3829 8115 3841
rect 8315 4017 8373 4029
rect 8315 3981 8327 4017
rect 8361 3981 8373 4017
rect 8315 3947 8373 3981
rect 8315 3911 8327 3947
rect 8361 3911 8373 3947
rect 8315 3876 8373 3911
rect 8315 3840 8327 3876
rect 8361 3840 8373 3876
rect 8315 3829 8373 3840
rect 8573 4017 8631 4029
rect 8573 3981 8585 4017
rect 8619 3981 8631 4017
rect 8573 3947 8631 3981
rect 8573 3911 8585 3947
rect 8619 3911 8631 3947
rect 8573 3877 8631 3911
rect 8573 3841 8585 3877
rect 8619 3841 8631 3877
rect 8573 3829 8631 3841
rect 8831 4017 8889 4029
rect 8831 3981 8843 4017
rect 8877 3981 8889 4017
rect 8831 3947 8889 3981
rect 8831 3911 8843 3947
rect 8877 3911 8889 3947
rect 8831 3877 8889 3911
rect 8831 3841 8843 3877
rect 8877 3841 8889 3877
rect 8831 3829 8889 3841
rect 9089 4017 9147 4029
rect 9089 3981 9101 4017
rect 9135 3981 9147 4017
rect 9089 3947 9147 3981
rect 9089 3911 9101 3947
rect 9135 3911 9147 3947
rect 9089 3877 9147 3911
rect 9089 3841 9101 3877
rect 9135 3841 9147 3877
rect 9089 3829 9147 3841
rect 9347 4017 9405 4029
rect 9347 3981 9359 4017
rect 9393 3981 9405 4017
rect 9347 3947 9405 3981
rect 9347 3911 9359 3947
rect 9393 3911 9405 3947
rect 9347 3877 9405 3911
rect 9347 3841 9359 3877
rect 9393 3841 9405 3877
rect 9347 3829 9405 3841
rect 9605 4017 9663 4029
rect 9605 3981 9617 4017
rect 9651 3981 9663 4017
rect 9605 3947 9663 3981
rect 9605 3911 9617 3947
rect 9651 3911 9663 3947
rect 9605 3877 9663 3911
rect 9605 3841 9617 3877
rect 9651 3841 9663 3877
rect 9605 3829 9663 3841
rect 9863 4017 9921 4029
rect 9863 3981 9875 4017
rect 9909 3981 9921 4017
rect 9863 3947 9921 3981
rect 9863 3911 9875 3947
rect 9909 3911 9921 3947
rect 9863 3877 9921 3911
rect 9863 3841 9875 3877
rect 9909 3841 9921 3877
rect 9863 3829 9921 3841
rect 10462 4018 10520 4030
rect 10462 3982 10474 4018
rect 10508 3982 10520 4018
rect 10462 3948 10520 3982
rect 10462 3912 10474 3948
rect 10508 3912 10520 3948
rect 10462 3878 10520 3912
rect 10462 3842 10474 3878
rect 10508 3842 10520 3878
rect 10462 3830 10520 3842
rect 10720 4018 10778 4030
rect 10720 3982 10732 4018
rect 10766 3982 10778 4018
rect 10720 3948 10778 3982
rect 10720 3912 10732 3948
rect 10766 3912 10778 3948
rect 10720 3878 10778 3912
rect 10720 3842 10732 3878
rect 10766 3842 10778 3878
rect 10720 3830 10778 3842
rect 10978 4018 11036 4030
rect 10978 3982 10990 4018
rect 11024 3982 11036 4018
rect 10978 3948 11036 3982
rect 10978 3912 10990 3948
rect 11024 3912 11036 3948
rect 10978 3877 11036 3912
rect 10978 3841 10990 3877
rect 11024 3841 11036 3877
rect 10978 3830 11036 3841
rect 11236 4018 11294 4030
rect 11236 3982 11248 4018
rect 11282 3982 11294 4018
rect 11236 3948 11294 3982
rect 11236 3912 11248 3948
rect 11282 3912 11294 3948
rect 11236 3878 11294 3912
rect 11236 3842 11248 3878
rect 11282 3842 11294 3878
rect 11236 3830 11294 3842
rect 11494 4018 11552 4030
rect 11494 3982 11506 4018
rect 11540 3982 11552 4018
rect 11494 3948 11552 3982
rect 11494 3912 11506 3948
rect 11540 3912 11552 3948
rect 11494 3878 11552 3912
rect 11494 3842 11506 3878
rect 11540 3842 11552 3878
rect 11494 3830 11552 3842
rect 11752 4018 11810 4030
rect 11752 3982 11764 4018
rect 11798 3982 11810 4018
rect 11752 3948 11810 3982
rect 11752 3912 11764 3948
rect 11798 3912 11810 3948
rect 11752 3878 11810 3912
rect 11752 3842 11764 3878
rect 11798 3842 11810 3878
rect 11752 3830 11810 3842
rect 12010 4018 12068 4030
rect 12010 3982 12022 4018
rect 12056 3982 12068 4018
rect 12010 3948 12068 3982
rect 12010 3912 12022 3948
rect 12056 3912 12068 3948
rect 12010 3878 12068 3912
rect 12010 3842 12022 3878
rect 12056 3842 12068 3878
rect 12010 3830 12068 3842
rect 12268 4018 12326 4030
rect 12268 3982 12280 4018
rect 12314 3982 12326 4018
rect 12268 3948 12326 3982
rect 12268 3912 12280 3948
rect 12314 3912 12326 3948
rect 12268 3878 12326 3912
rect 12268 3842 12280 3878
rect 12314 3842 12326 3878
rect 12268 3830 12326 3842
rect 12526 4018 12584 4030
rect 12526 3982 12538 4018
rect 12572 3982 12584 4018
rect 12526 3948 12584 3982
rect 12526 3912 12538 3948
rect 12572 3912 12584 3948
rect 12526 3878 12584 3912
rect 12526 3842 12538 3878
rect 12572 3842 12584 3878
rect 12526 3830 12584 3842
rect 5009 3363 5067 3377
rect 5009 3329 5021 3363
rect 5055 3329 5067 3363
rect 5009 3295 5067 3329
rect 5009 3259 5021 3295
rect 5055 3259 5067 3295
rect 5009 3225 5067 3259
rect 5009 3191 5021 3225
rect 5055 3191 5067 3225
rect 5009 3177 5067 3191
rect 5267 3363 5325 3377
rect 5267 3329 5279 3363
rect 5313 3329 5325 3363
rect 5267 3295 5325 3329
rect 5267 3259 5279 3295
rect 5313 3259 5325 3295
rect 5267 3225 5325 3259
rect 5267 3191 5279 3225
rect 5313 3191 5325 3225
rect 5267 3177 5325 3191
rect 5549 3363 5607 3377
rect 5549 3329 5561 3363
rect 5595 3329 5607 3363
rect 5549 3295 5607 3329
rect 5549 3259 5561 3295
rect 5595 3259 5607 3295
rect 5549 3225 5607 3259
rect 5549 3191 5561 3225
rect 5595 3191 5607 3225
rect 5549 3177 5607 3191
rect 5807 3363 5865 3377
rect 5807 3329 5819 3363
rect 5853 3329 5865 3363
rect 5807 3295 5865 3329
rect 5807 3259 5819 3295
rect 5853 3259 5865 3295
rect 5807 3225 5865 3259
rect 5807 3191 5819 3225
rect 5853 3191 5865 3225
rect 5807 3177 5865 3191
rect 6029 3363 6087 3377
rect 6029 3329 6041 3363
rect 6075 3329 6087 3363
rect 6029 3295 6087 3329
rect 6029 3259 6041 3295
rect 6075 3259 6087 3295
rect 6029 3225 6087 3259
rect 6029 3191 6041 3225
rect 6075 3191 6087 3225
rect 6029 3177 6087 3191
rect 6287 3363 6345 3377
rect 6287 3329 6299 3363
rect 6333 3329 6345 3363
rect 6287 3295 6345 3329
rect 6287 3259 6299 3295
rect 6333 3259 6345 3295
rect 6287 3225 6345 3259
rect 6287 3191 6299 3225
rect 6333 3191 6345 3225
rect 6287 3177 6345 3191
rect 6532 3365 6590 3379
rect 6532 3331 6544 3365
rect 6578 3331 6590 3365
rect 6532 3297 6590 3331
rect 6532 3261 6544 3297
rect 6578 3261 6590 3297
rect 6532 3227 6590 3261
rect 6532 3193 6544 3227
rect 6578 3193 6590 3227
rect 6532 3179 6590 3193
rect 6790 3365 6848 3379
rect 6790 3331 6802 3365
rect 6836 3331 6848 3365
rect 6790 3297 6848 3331
rect 6790 3261 6802 3297
rect 6836 3261 6848 3297
rect 6790 3227 6848 3261
rect 6790 3193 6802 3227
rect 6836 3193 6848 3227
rect 6790 3179 6848 3193
rect 7042 3375 7100 3389
rect 7042 3341 7054 3375
rect 7088 3341 7100 3375
rect 7042 3307 7100 3341
rect 7042 3271 7054 3307
rect 7088 3271 7100 3307
rect 7042 3237 7100 3271
rect 7042 3203 7054 3237
rect 7088 3203 7100 3237
rect 7042 3189 7100 3203
rect 7300 3375 7358 3389
rect 7300 3341 7312 3375
rect 7346 3341 7358 3375
rect 7300 3307 7358 3341
rect 7300 3271 7312 3307
rect 7346 3271 7358 3307
rect 7300 3237 7358 3271
rect 7300 3203 7312 3237
rect 7346 3203 7358 3237
rect 7300 3189 7358 3203
rect 7679 3363 7737 3377
rect 7679 3329 7691 3363
rect 7725 3329 7737 3363
rect 7679 3295 7737 3329
rect 7679 3259 7691 3295
rect 7725 3259 7737 3295
rect 7679 3225 7737 3259
rect 7679 3191 7691 3225
rect 7725 3191 7737 3225
rect 7679 3177 7737 3191
rect 7937 3363 7995 3377
rect 7937 3329 7949 3363
rect 7983 3329 7995 3363
rect 7937 3295 7995 3329
rect 7937 3259 7949 3295
rect 7983 3259 7995 3295
rect 7937 3225 7995 3259
rect 7937 3191 7949 3225
rect 7983 3191 7995 3225
rect 7937 3177 7995 3191
rect 8219 3363 8277 3377
rect 8219 3329 8231 3363
rect 8265 3329 8277 3363
rect 8219 3295 8277 3329
rect 8219 3259 8231 3295
rect 8265 3259 8277 3295
rect 8219 3225 8277 3259
rect 8219 3191 8231 3225
rect 8265 3191 8277 3225
rect 8219 3177 8277 3191
rect 8477 3363 8535 3377
rect 8477 3329 8489 3363
rect 8523 3329 8535 3363
rect 8477 3295 8535 3329
rect 8477 3259 8489 3295
rect 8523 3259 8535 3295
rect 8477 3225 8535 3259
rect 8477 3191 8489 3225
rect 8523 3191 8535 3225
rect 8477 3177 8535 3191
rect 8699 3363 8757 3377
rect 8699 3329 8711 3363
rect 8745 3329 8757 3363
rect 8699 3295 8757 3329
rect 8699 3259 8711 3295
rect 8745 3259 8757 3295
rect 8699 3225 8757 3259
rect 8699 3191 8711 3225
rect 8745 3191 8757 3225
rect 8699 3177 8757 3191
rect 8957 3363 9015 3377
rect 8957 3329 8969 3363
rect 9003 3329 9015 3363
rect 8957 3295 9015 3329
rect 8957 3259 8969 3295
rect 9003 3259 9015 3295
rect 8957 3225 9015 3259
rect 8957 3191 8969 3225
rect 9003 3191 9015 3225
rect 8957 3177 9015 3191
rect 9202 3365 9260 3379
rect 9202 3331 9214 3365
rect 9248 3331 9260 3365
rect 9202 3297 9260 3331
rect 9202 3261 9214 3297
rect 9248 3261 9260 3297
rect 9202 3227 9260 3261
rect 9202 3193 9214 3227
rect 9248 3193 9260 3227
rect 9202 3179 9260 3193
rect 9460 3365 9518 3379
rect 9460 3331 9472 3365
rect 9506 3331 9518 3365
rect 9460 3297 9518 3331
rect 9460 3261 9472 3297
rect 9506 3261 9518 3297
rect 9460 3227 9518 3261
rect 9460 3193 9472 3227
rect 9506 3193 9518 3227
rect 9460 3179 9518 3193
rect 9712 3375 9770 3389
rect 9712 3341 9724 3375
rect 9758 3341 9770 3375
rect 9712 3307 9770 3341
rect 9712 3271 9724 3307
rect 9758 3271 9770 3307
rect 9712 3237 9770 3271
rect 9712 3203 9724 3237
rect 9758 3203 9770 3237
rect 9712 3189 9770 3203
rect 9970 3375 10028 3389
rect 9970 3341 9982 3375
rect 10016 3341 10028 3375
rect 9970 3307 10028 3341
rect 9970 3271 9982 3307
rect 10016 3271 10028 3307
rect 9970 3237 10028 3271
rect 9970 3203 9982 3237
rect 10016 3203 10028 3237
rect 9970 3189 10028 3203
rect 10342 3364 10400 3378
rect 10342 3330 10354 3364
rect 10388 3330 10400 3364
rect 10342 3296 10400 3330
rect 10342 3260 10354 3296
rect 10388 3260 10400 3296
rect 10342 3226 10400 3260
rect 10342 3192 10354 3226
rect 10388 3192 10400 3226
rect 10342 3178 10400 3192
rect 10600 3364 10658 3378
rect 10600 3330 10612 3364
rect 10646 3330 10658 3364
rect 10600 3296 10658 3330
rect 10600 3260 10612 3296
rect 10646 3260 10658 3296
rect 10600 3226 10658 3260
rect 10600 3192 10612 3226
rect 10646 3192 10658 3226
rect 10600 3178 10658 3192
rect 10882 3364 10940 3378
rect 10882 3330 10894 3364
rect 10928 3330 10940 3364
rect 10882 3296 10940 3330
rect 10882 3260 10894 3296
rect 10928 3260 10940 3296
rect 10882 3226 10940 3260
rect 10882 3192 10894 3226
rect 10928 3192 10940 3226
rect 10882 3178 10940 3192
rect 11140 3364 11198 3378
rect 11140 3330 11152 3364
rect 11186 3330 11198 3364
rect 11140 3296 11198 3330
rect 11140 3260 11152 3296
rect 11186 3260 11198 3296
rect 11140 3226 11198 3260
rect 11140 3192 11152 3226
rect 11186 3192 11198 3226
rect 11140 3178 11198 3192
rect 11362 3364 11420 3378
rect 11362 3330 11374 3364
rect 11408 3330 11420 3364
rect 11362 3296 11420 3330
rect 11362 3260 11374 3296
rect 11408 3260 11420 3296
rect 11362 3226 11420 3260
rect 11362 3192 11374 3226
rect 11408 3192 11420 3226
rect 11362 3178 11420 3192
rect 11620 3364 11678 3378
rect 11620 3330 11632 3364
rect 11666 3330 11678 3364
rect 11620 3296 11678 3330
rect 11620 3260 11632 3296
rect 11666 3260 11678 3296
rect 11620 3226 11678 3260
rect 11620 3192 11632 3226
rect 11666 3192 11678 3226
rect 11620 3178 11678 3192
rect 11865 3366 11923 3380
rect 11865 3332 11877 3366
rect 11911 3332 11923 3366
rect 11865 3298 11923 3332
rect 11865 3262 11877 3298
rect 11911 3262 11923 3298
rect 11865 3228 11923 3262
rect 11865 3194 11877 3228
rect 11911 3194 11923 3228
rect 11865 3180 11923 3194
rect 12123 3366 12181 3380
rect 12123 3332 12135 3366
rect 12169 3332 12181 3366
rect 12123 3298 12181 3332
rect 12123 3262 12135 3298
rect 12169 3262 12181 3298
rect 12123 3228 12181 3262
rect 12123 3194 12135 3228
rect 12169 3194 12181 3228
rect 12123 3180 12181 3194
rect 12375 3376 12433 3390
rect 12375 3342 12387 3376
rect 12421 3342 12433 3376
rect 12375 3308 12433 3342
rect 12375 3272 12387 3308
rect 12421 3272 12433 3308
rect 12375 3238 12433 3272
rect 12375 3204 12387 3238
rect 12421 3204 12433 3238
rect 12375 3190 12433 3204
rect 12633 3376 12691 3390
rect 12633 3342 12645 3376
rect 12679 3342 12691 3376
rect 12633 3308 12691 3342
rect 12633 3272 12645 3308
rect 12679 3272 12691 3308
rect 12633 3238 12691 3272
rect 12633 3204 12645 3238
rect 12679 3204 12691 3238
rect 12633 3190 12691 3204
rect 5129 808 5187 820
rect 5129 772 5141 808
rect 5175 772 5187 808
rect 5129 738 5187 772
rect 5129 702 5141 738
rect 5175 702 5187 738
rect 5129 668 5187 702
rect 5129 632 5141 668
rect 5175 632 5187 668
rect 5129 620 5187 632
rect 5387 808 5445 820
rect 5387 772 5399 808
rect 5433 772 5445 808
rect 5387 738 5445 772
rect 5387 702 5399 738
rect 5433 702 5445 738
rect 5387 668 5445 702
rect 5387 632 5399 668
rect 5433 632 5445 668
rect 5387 620 5445 632
rect 5645 808 5703 820
rect 5645 772 5657 808
rect 5691 772 5703 808
rect 5645 738 5703 772
rect 5645 702 5657 738
rect 5691 702 5703 738
rect 5645 667 5703 702
rect 5645 631 5657 667
rect 5691 631 5703 667
rect 5645 620 5703 631
rect 5903 808 5961 820
rect 5903 772 5915 808
rect 5949 772 5961 808
rect 5903 738 5961 772
rect 5903 702 5915 738
rect 5949 702 5961 738
rect 5903 668 5961 702
rect 5903 632 5915 668
rect 5949 632 5961 668
rect 5903 620 5961 632
rect 6161 808 6219 820
rect 6161 772 6173 808
rect 6207 772 6219 808
rect 6161 738 6219 772
rect 6161 702 6173 738
rect 6207 702 6219 738
rect 6161 668 6219 702
rect 6161 632 6173 668
rect 6207 632 6219 668
rect 6161 620 6219 632
rect 6419 808 6477 820
rect 6419 772 6431 808
rect 6465 772 6477 808
rect 6419 738 6477 772
rect 6419 702 6431 738
rect 6465 702 6477 738
rect 6419 668 6477 702
rect 6419 632 6431 668
rect 6465 632 6477 668
rect 6419 620 6477 632
rect 6677 808 6735 820
rect 6677 772 6689 808
rect 6723 772 6735 808
rect 6677 738 6735 772
rect 6677 702 6689 738
rect 6723 702 6735 738
rect 6677 668 6735 702
rect 6677 632 6689 668
rect 6723 632 6735 668
rect 6677 620 6735 632
rect 6935 808 6993 820
rect 6935 772 6947 808
rect 6981 772 6993 808
rect 6935 738 6993 772
rect 6935 702 6947 738
rect 6981 702 6993 738
rect 6935 668 6993 702
rect 6935 632 6947 668
rect 6981 632 6993 668
rect 6935 620 6993 632
rect 7193 808 7251 820
rect 7193 772 7205 808
rect 7239 772 7251 808
rect 7193 738 7251 772
rect 7193 702 7205 738
rect 7239 702 7251 738
rect 7193 668 7251 702
rect 7193 632 7205 668
rect 7239 632 7251 668
rect 7193 620 7251 632
rect 7799 808 7857 820
rect 7799 772 7811 808
rect 7845 772 7857 808
rect 7799 738 7857 772
rect 7799 702 7811 738
rect 7845 702 7857 738
rect 7799 668 7857 702
rect 7799 632 7811 668
rect 7845 632 7857 668
rect 7799 620 7857 632
rect 8057 808 8115 820
rect 8057 772 8069 808
rect 8103 772 8115 808
rect 8057 738 8115 772
rect 8057 702 8069 738
rect 8103 702 8115 738
rect 8057 668 8115 702
rect 8057 632 8069 668
rect 8103 632 8115 668
rect 8057 620 8115 632
rect 8315 808 8373 820
rect 8315 772 8327 808
rect 8361 772 8373 808
rect 8315 738 8373 772
rect 8315 702 8327 738
rect 8361 702 8373 738
rect 8315 667 8373 702
rect 8315 631 8327 667
rect 8361 631 8373 667
rect 8315 620 8373 631
rect 8573 808 8631 820
rect 8573 772 8585 808
rect 8619 772 8631 808
rect 8573 738 8631 772
rect 8573 702 8585 738
rect 8619 702 8631 738
rect 8573 668 8631 702
rect 8573 632 8585 668
rect 8619 632 8631 668
rect 8573 620 8631 632
rect 8831 808 8889 820
rect 8831 772 8843 808
rect 8877 772 8889 808
rect 8831 738 8889 772
rect 8831 702 8843 738
rect 8877 702 8889 738
rect 8831 668 8889 702
rect 8831 632 8843 668
rect 8877 632 8889 668
rect 8831 620 8889 632
rect 9089 808 9147 820
rect 9089 772 9101 808
rect 9135 772 9147 808
rect 9089 738 9147 772
rect 9089 702 9101 738
rect 9135 702 9147 738
rect 9089 668 9147 702
rect 9089 632 9101 668
rect 9135 632 9147 668
rect 9089 620 9147 632
rect 9347 808 9405 820
rect 9347 772 9359 808
rect 9393 772 9405 808
rect 9347 738 9405 772
rect 9347 702 9359 738
rect 9393 702 9405 738
rect 9347 668 9405 702
rect 9347 632 9359 668
rect 9393 632 9405 668
rect 9347 620 9405 632
rect 9605 808 9663 820
rect 9605 772 9617 808
rect 9651 772 9663 808
rect 9605 738 9663 772
rect 9605 702 9617 738
rect 9651 702 9663 738
rect 9605 668 9663 702
rect 9605 632 9617 668
rect 9651 632 9663 668
rect 9605 620 9663 632
rect 9863 808 9921 820
rect 9863 772 9875 808
rect 9909 772 9921 808
rect 9863 738 9921 772
rect 9863 702 9875 738
rect 9909 702 9921 738
rect 9863 668 9921 702
rect 9863 632 9875 668
rect 9909 632 9921 668
rect 9863 620 9921 632
rect 10462 809 10520 821
rect 10462 773 10474 809
rect 10508 773 10520 809
rect 10462 739 10520 773
rect 10462 703 10474 739
rect 10508 703 10520 739
rect 10462 669 10520 703
rect 10462 633 10474 669
rect 10508 633 10520 669
rect 10462 621 10520 633
rect 10720 809 10778 821
rect 10720 773 10732 809
rect 10766 773 10778 809
rect 10720 739 10778 773
rect 10720 703 10732 739
rect 10766 703 10778 739
rect 10720 669 10778 703
rect 10720 633 10732 669
rect 10766 633 10778 669
rect 10720 621 10778 633
rect 10978 809 11036 821
rect 10978 773 10990 809
rect 11024 773 11036 809
rect 10978 739 11036 773
rect 10978 703 10990 739
rect 11024 703 11036 739
rect 10978 668 11036 703
rect 10978 632 10990 668
rect 11024 632 11036 668
rect 10978 621 11036 632
rect 11236 809 11294 821
rect 11236 773 11248 809
rect 11282 773 11294 809
rect 11236 739 11294 773
rect 11236 703 11248 739
rect 11282 703 11294 739
rect 11236 669 11294 703
rect 11236 633 11248 669
rect 11282 633 11294 669
rect 11236 621 11294 633
rect 11494 809 11552 821
rect 11494 773 11506 809
rect 11540 773 11552 809
rect 11494 739 11552 773
rect 11494 703 11506 739
rect 11540 703 11552 739
rect 11494 669 11552 703
rect 11494 633 11506 669
rect 11540 633 11552 669
rect 11494 621 11552 633
rect 11752 809 11810 821
rect 11752 773 11764 809
rect 11798 773 11810 809
rect 11752 739 11810 773
rect 11752 703 11764 739
rect 11798 703 11810 739
rect 11752 669 11810 703
rect 11752 633 11764 669
rect 11798 633 11810 669
rect 11752 621 11810 633
rect 12010 809 12068 821
rect 12010 773 12022 809
rect 12056 773 12068 809
rect 12010 739 12068 773
rect 12010 703 12022 739
rect 12056 703 12068 739
rect 12010 669 12068 703
rect 12010 633 12022 669
rect 12056 633 12068 669
rect 12010 621 12068 633
rect 12268 809 12326 821
rect 12268 773 12280 809
rect 12314 773 12326 809
rect 12268 739 12326 773
rect 12268 703 12280 739
rect 12314 703 12326 739
rect 12268 669 12326 703
rect 12268 633 12280 669
rect 12314 633 12326 669
rect 12268 621 12326 633
rect 12526 809 12584 821
rect 12526 773 12538 809
rect 12572 773 12584 809
rect 12526 739 12584 773
rect 12526 703 12538 739
rect 12572 703 12584 739
rect 12526 669 12584 703
rect 12526 633 12538 669
rect 12572 633 12584 669
rect 12526 621 12584 633
rect 5129 390 5187 402
rect 5129 354 5141 390
rect 5175 354 5187 390
rect 5129 320 5187 354
rect 5129 284 5141 320
rect 5175 284 5187 320
rect 5129 250 5187 284
rect 5129 214 5141 250
rect 5175 214 5187 250
rect 5129 202 5187 214
rect 5387 390 5445 402
rect 5387 354 5399 390
rect 5433 354 5445 390
rect 5387 320 5445 354
rect 5387 284 5399 320
rect 5433 284 5445 320
rect 5387 250 5445 284
rect 5387 214 5399 250
rect 5433 214 5445 250
rect 5387 202 5445 214
rect 5645 390 5703 402
rect 5645 354 5657 390
rect 5691 354 5703 390
rect 5645 320 5703 354
rect 5645 284 5657 320
rect 5691 284 5703 320
rect 5645 249 5703 284
rect 5645 213 5657 249
rect 5691 213 5703 249
rect 5645 202 5703 213
rect 5903 390 5961 402
rect 5903 354 5915 390
rect 5949 354 5961 390
rect 5903 320 5961 354
rect 5903 284 5915 320
rect 5949 284 5961 320
rect 5903 250 5961 284
rect 5903 214 5915 250
rect 5949 214 5961 250
rect 5903 202 5961 214
rect 6161 390 6219 402
rect 6161 354 6173 390
rect 6207 354 6219 390
rect 6161 320 6219 354
rect 6161 284 6173 320
rect 6207 284 6219 320
rect 6161 250 6219 284
rect 6161 214 6173 250
rect 6207 214 6219 250
rect 6161 202 6219 214
rect 6419 390 6477 402
rect 6419 354 6431 390
rect 6465 354 6477 390
rect 6419 320 6477 354
rect 6419 284 6431 320
rect 6465 284 6477 320
rect 6419 250 6477 284
rect 6419 214 6431 250
rect 6465 214 6477 250
rect 6419 202 6477 214
rect 6677 390 6735 402
rect 6677 354 6689 390
rect 6723 354 6735 390
rect 6677 320 6735 354
rect 6677 284 6689 320
rect 6723 284 6735 320
rect 6677 250 6735 284
rect 6677 214 6689 250
rect 6723 214 6735 250
rect 6677 202 6735 214
rect 6935 390 6993 402
rect 6935 354 6947 390
rect 6981 354 6993 390
rect 6935 320 6993 354
rect 6935 284 6947 320
rect 6981 284 6993 320
rect 6935 250 6993 284
rect 6935 214 6947 250
rect 6981 214 6993 250
rect 6935 202 6993 214
rect 7193 390 7251 402
rect 7193 354 7205 390
rect 7239 354 7251 390
rect 7193 320 7251 354
rect 7193 284 7205 320
rect 7239 284 7251 320
rect 7193 250 7251 284
rect 7193 214 7205 250
rect 7239 214 7251 250
rect 7193 202 7251 214
rect 7799 390 7857 402
rect 7799 354 7811 390
rect 7845 354 7857 390
rect 7799 320 7857 354
rect 7799 284 7811 320
rect 7845 284 7857 320
rect 7799 250 7857 284
rect 7799 214 7811 250
rect 7845 214 7857 250
rect 7799 202 7857 214
rect 8057 390 8115 402
rect 8057 354 8069 390
rect 8103 354 8115 390
rect 8057 320 8115 354
rect 8057 284 8069 320
rect 8103 284 8115 320
rect 8057 250 8115 284
rect 8057 214 8069 250
rect 8103 214 8115 250
rect 8057 202 8115 214
rect 8315 390 8373 402
rect 8315 354 8327 390
rect 8361 354 8373 390
rect 8315 320 8373 354
rect 8315 284 8327 320
rect 8361 284 8373 320
rect 8315 249 8373 284
rect 8315 213 8327 249
rect 8361 213 8373 249
rect 8315 202 8373 213
rect 8573 390 8631 402
rect 8573 354 8585 390
rect 8619 354 8631 390
rect 8573 320 8631 354
rect 8573 284 8585 320
rect 8619 284 8631 320
rect 8573 250 8631 284
rect 8573 214 8585 250
rect 8619 214 8631 250
rect 8573 202 8631 214
rect 8831 390 8889 402
rect 8831 354 8843 390
rect 8877 354 8889 390
rect 8831 320 8889 354
rect 8831 284 8843 320
rect 8877 284 8889 320
rect 8831 250 8889 284
rect 8831 214 8843 250
rect 8877 214 8889 250
rect 8831 202 8889 214
rect 9089 390 9147 402
rect 9089 354 9101 390
rect 9135 354 9147 390
rect 9089 320 9147 354
rect 9089 284 9101 320
rect 9135 284 9147 320
rect 9089 250 9147 284
rect 9089 214 9101 250
rect 9135 214 9147 250
rect 9089 202 9147 214
rect 9347 390 9405 402
rect 9347 354 9359 390
rect 9393 354 9405 390
rect 9347 320 9405 354
rect 9347 284 9359 320
rect 9393 284 9405 320
rect 9347 250 9405 284
rect 9347 214 9359 250
rect 9393 214 9405 250
rect 9347 202 9405 214
rect 9605 390 9663 402
rect 9605 354 9617 390
rect 9651 354 9663 390
rect 9605 320 9663 354
rect 9605 284 9617 320
rect 9651 284 9663 320
rect 9605 250 9663 284
rect 9605 214 9617 250
rect 9651 214 9663 250
rect 9605 202 9663 214
rect 9863 390 9921 402
rect 9863 354 9875 390
rect 9909 354 9921 390
rect 9863 320 9921 354
rect 9863 284 9875 320
rect 9909 284 9921 320
rect 9863 250 9921 284
rect 9863 214 9875 250
rect 9909 214 9921 250
rect 9863 202 9921 214
rect 10462 391 10520 403
rect 10462 355 10474 391
rect 10508 355 10520 391
rect 10462 321 10520 355
rect 10462 285 10474 321
rect 10508 285 10520 321
rect 10462 251 10520 285
rect 10462 215 10474 251
rect 10508 215 10520 251
rect 10462 203 10520 215
rect 10720 391 10778 403
rect 10720 355 10732 391
rect 10766 355 10778 391
rect 10720 321 10778 355
rect 10720 285 10732 321
rect 10766 285 10778 321
rect 10720 251 10778 285
rect 10720 215 10732 251
rect 10766 215 10778 251
rect 10720 203 10778 215
rect 10978 391 11036 403
rect 10978 355 10990 391
rect 11024 355 11036 391
rect 10978 321 11036 355
rect 10978 285 10990 321
rect 11024 285 11036 321
rect 10978 250 11036 285
rect 10978 214 10990 250
rect 11024 214 11036 250
rect 10978 203 11036 214
rect 11236 391 11294 403
rect 11236 355 11248 391
rect 11282 355 11294 391
rect 11236 321 11294 355
rect 11236 285 11248 321
rect 11282 285 11294 321
rect 11236 251 11294 285
rect 11236 215 11248 251
rect 11282 215 11294 251
rect 11236 203 11294 215
rect 11494 391 11552 403
rect 11494 355 11506 391
rect 11540 355 11552 391
rect 11494 321 11552 355
rect 11494 285 11506 321
rect 11540 285 11552 321
rect 11494 251 11552 285
rect 11494 215 11506 251
rect 11540 215 11552 251
rect 11494 203 11552 215
rect 11752 391 11810 403
rect 11752 355 11764 391
rect 11798 355 11810 391
rect 11752 321 11810 355
rect 11752 285 11764 321
rect 11798 285 11810 321
rect 11752 251 11810 285
rect 11752 215 11764 251
rect 11798 215 11810 251
rect 11752 203 11810 215
rect 12010 391 12068 403
rect 12010 355 12022 391
rect 12056 355 12068 391
rect 12010 321 12068 355
rect 12010 285 12022 321
rect 12056 285 12068 321
rect 12010 251 12068 285
rect 12010 215 12022 251
rect 12056 215 12068 251
rect 12010 203 12068 215
rect 12268 391 12326 403
rect 12268 355 12280 391
rect 12314 355 12326 391
rect 12268 321 12326 355
rect 12268 285 12280 321
rect 12314 285 12326 321
rect 12268 251 12326 285
rect 12268 215 12280 251
rect 12314 215 12326 251
rect 12268 203 12326 215
rect 12526 391 12584 403
rect 12526 355 12538 391
rect 12572 355 12584 391
rect 12526 321 12584 355
rect 12526 285 12538 321
rect 12572 285 12584 321
rect 12526 251 12584 285
rect 12526 215 12538 251
rect 12572 215 12584 251
rect 12526 203 12584 215
rect 5129 -28 5187 -16
rect 5129 -64 5141 -28
rect 5175 -64 5187 -28
rect 5129 -98 5187 -64
rect 5129 -134 5141 -98
rect 5175 -134 5187 -98
rect 5129 -168 5187 -134
rect 5129 -204 5141 -168
rect 5175 -204 5187 -168
rect 5129 -216 5187 -204
rect 5387 -28 5445 -16
rect 5387 -64 5399 -28
rect 5433 -64 5445 -28
rect 5387 -98 5445 -64
rect 5387 -134 5399 -98
rect 5433 -134 5445 -98
rect 5387 -168 5445 -134
rect 5387 -204 5399 -168
rect 5433 -204 5445 -168
rect 5387 -216 5445 -204
rect 5645 -28 5703 -16
rect 5645 -64 5657 -28
rect 5691 -64 5703 -28
rect 5645 -98 5703 -64
rect 5645 -134 5657 -98
rect 5691 -134 5703 -98
rect 5645 -169 5703 -134
rect 5645 -205 5657 -169
rect 5691 -205 5703 -169
rect 5645 -216 5703 -205
rect 5903 -28 5961 -16
rect 5903 -64 5915 -28
rect 5949 -64 5961 -28
rect 5903 -98 5961 -64
rect 5903 -134 5915 -98
rect 5949 -134 5961 -98
rect 5903 -168 5961 -134
rect 5903 -204 5915 -168
rect 5949 -204 5961 -168
rect 5903 -216 5961 -204
rect 6161 -28 6219 -16
rect 6161 -64 6173 -28
rect 6207 -64 6219 -28
rect 6161 -98 6219 -64
rect 6161 -134 6173 -98
rect 6207 -134 6219 -98
rect 6161 -168 6219 -134
rect 6161 -204 6173 -168
rect 6207 -204 6219 -168
rect 6161 -216 6219 -204
rect 6419 -28 6477 -16
rect 6419 -64 6431 -28
rect 6465 -64 6477 -28
rect 6419 -98 6477 -64
rect 6419 -134 6431 -98
rect 6465 -134 6477 -98
rect 6419 -168 6477 -134
rect 6419 -204 6431 -168
rect 6465 -204 6477 -168
rect 6419 -216 6477 -204
rect 6677 -28 6735 -16
rect 6677 -64 6689 -28
rect 6723 -64 6735 -28
rect 6677 -98 6735 -64
rect 6677 -134 6689 -98
rect 6723 -134 6735 -98
rect 6677 -168 6735 -134
rect 6677 -204 6689 -168
rect 6723 -204 6735 -168
rect 6677 -216 6735 -204
rect 6935 -28 6993 -16
rect 6935 -64 6947 -28
rect 6981 -64 6993 -28
rect 6935 -98 6993 -64
rect 6935 -134 6947 -98
rect 6981 -134 6993 -98
rect 6935 -168 6993 -134
rect 6935 -204 6947 -168
rect 6981 -204 6993 -168
rect 6935 -216 6993 -204
rect 7193 -28 7251 -16
rect 7193 -64 7205 -28
rect 7239 -64 7251 -28
rect 7193 -98 7251 -64
rect 7193 -134 7205 -98
rect 7239 -134 7251 -98
rect 7193 -168 7251 -134
rect 7193 -204 7205 -168
rect 7239 -204 7251 -168
rect 7193 -216 7251 -204
rect 7799 -28 7857 -16
rect 7799 -64 7811 -28
rect 7845 -64 7857 -28
rect 7799 -98 7857 -64
rect 7799 -134 7811 -98
rect 7845 -134 7857 -98
rect 7799 -168 7857 -134
rect 7799 -204 7811 -168
rect 7845 -204 7857 -168
rect 7799 -216 7857 -204
rect 8057 -28 8115 -16
rect 8057 -64 8069 -28
rect 8103 -64 8115 -28
rect 8057 -98 8115 -64
rect 8057 -134 8069 -98
rect 8103 -134 8115 -98
rect 8057 -168 8115 -134
rect 8057 -204 8069 -168
rect 8103 -204 8115 -168
rect 8057 -216 8115 -204
rect 8315 -28 8373 -16
rect 8315 -64 8327 -28
rect 8361 -64 8373 -28
rect 8315 -98 8373 -64
rect 8315 -134 8327 -98
rect 8361 -134 8373 -98
rect 8315 -169 8373 -134
rect 8315 -205 8327 -169
rect 8361 -205 8373 -169
rect 8315 -216 8373 -205
rect 8573 -28 8631 -16
rect 8573 -64 8585 -28
rect 8619 -64 8631 -28
rect 8573 -98 8631 -64
rect 8573 -134 8585 -98
rect 8619 -134 8631 -98
rect 8573 -168 8631 -134
rect 8573 -204 8585 -168
rect 8619 -204 8631 -168
rect 8573 -216 8631 -204
rect 8831 -28 8889 -16
rect 8831 -64 8843 -28
rect 8877 -64 8889 -28
rect 8831 -98 8889 -64
rect 8831 -134 8843 -98
rect 8877 -134 8889 -98
rect 8831 -168 8889 -134
rect 8831 -204 8843 -168
rect 8877 -204 8889 -168
rect 8831 -216 8889 -204
rect 9089 -28 9147 -16
rect 9089 -64 9101 -28
rect 9135 -64 9147 -28
rect 9089 -98 9147 -64
rect 9089 -134 9101 -98
rect 9135 -134 9147 -98
rect 9089 -168 9147 -134
rect 9089 -204 9101 -168
rect 9135 -204 9147 -168
rect 9089 -216 9147 -204
rect 9347 -28 9405 -16
rect 9347 -64 9359 -28
rect 9393 -64 9405 -28
rect 9347 -98 9405 -64
rect 9347 -134 9359 -98
rect 9393 -134 9405 -98
rect 9347 -168 9405 -134
rect 9347 -204 9359 -168
rect 9393 -204 9405 -168
rect 9347 -216 9405 -204
rect 9605 -28 9663 -16
rect 9605 -64 9617 -28
rect 9651 -64 9663 -28
rect 9605 -98 9663 -64
rect 9605 -134 9617 -98
rect 9651 -134 9663 -98
rect 9605 -168 9663 -134
rect 9605 -204 9617 -168
rect 9651 -204 9663 -168
rect 9605 -216 9663 -204
rect 9863 -28 9921 -16
rect 9863 -64 9875 -28
rect 9909 -64 9921 -28
rect 9863 -98 9921 -64
rect 9863 -134 9875 -98
rect 9909 -134 9921 -98
rect 9863 -168 9921 -134
rect 9863 -204 9875 -168
rect 9909 -204 9921 -168
rect 9863 -216 9921 -204
rect 10462 -27 10520 -15
rect 10462 -63 10474 -27
rect 10508 -63 10520 -27
rect 10462 -97 10520 -63
rect 10462 -133 10474 -97
rect 10508 -133 10520 -97
rect 10462 -167 10520 -133
rect 10462 -203 10474 -167
rect 10508 -203 10520 -167
rect 10462 -215 10520 -203
rect 10720 -27 10778 -15
rect 10720 -63 10732 -27
rect 10766 -63 10778 -27
rect 10720 -97 10778 -63
rect 10720 -133 10732 -97
rect 10766 -133 10778 -97
rect 10720 -167 10778 -133
rect 10720 -203 10732 -167
rect 10766 -203 10778 -167
rect 10720 -215 10778 -203
rect 10978 -27 11036 -15
rect 10978 -63 10990 -27
rect 11024 -63 11036 -27
rect 10978 -97 11036 -63
rect 10978 -133 10990 -97
rect 11024 -133 11036 -97
rect 10978 -168 11036 -133
rect 10978 -204 10990 -168
rect 11024 -204 11036 -168
rect 10978 -215 11036 -204
rect 11236 -27 11294 -15
rect 11236 -63 11248 -27
rect 11282 -63 11294 -27
rect 11236 -97 11294 -63
rect 11236 -133 11248 -97
rect 11282 -133 11294 -97
rect 11236 -167 11294 -133
rect 11236 -203 11248 -167
rect 11282 -203 11294 -167
rect 11236 -215 11294 -203
rect 11494 -27 11552 -15
rect 11494 -63 11506 -27
rect 11540 -63 11552 -27
rect 11494 -97 11552 -63
rect 11494 -133 11506 -97
rect 11540 -133 11552 -97
rect 11494 -167 11552 -133
rect 11494 -203 11506 -167
rect 11540 -203 11552 -167
rect 11494 -215 11552 -203
rect 11752 -27 11810 -15
rect 11752 -63 11764 -27
rect 11798 -63 11810 -27
rect 11752 -97 11810 -63
rect 11752 -133 11764 -97
rect 11798 -133 11810 -97
rect 11752 -167 11810 -133
rect 11752 -203 11764 -167
rect 11798 -203 11810 -167
rect 11752 -215 11810 -203
rect 12010 -27 12068 -15
rect 12010 -63 12022 -27
rect 12056 -63 12068 -27
rect 12010 -97 12068 -63
rect 12010 -133 12022 -97
rect 12056 -133 12068 -97
rect 12010 -167 12068 -133
rect 12010 -203 12022 -167
rect 12056 -203 12068 -167
rect 12010 -215 12068 -203
rect 12268 -27 12326 -15
rect 12268 -63 12280 -27
rect 12314 -63 12326 -27
rect 12268 -97 12326 -63
rect 12268 -133 12280 -97
rect 12314 -133 12326 -97
rect 12268 -167 12326 -133
rect 12268 -203 12280 -167
rect 12314 -203 12326 -167
rect 12268 -215 12326 -203
rect 12526 -27 12584 -15
rect 12526 -63 12538 -27
rect 12572 -63 12584 -27
rect 12526 -97 12584 -63
rect 12526 -133 12538 -97
rect 12572 -133 12584 -97
rect 12526 -167 12584 -133
rect 12526 -203 12538 -167
rect 12572 -203 12584 -167
rect 12526 -215 12584 -203
rect 5129 -446 5187 -434
rect 5129 -482 5141 -446
rect 5175 -482 5187 -446
rect 5129 -516 5187 -482
rect 5129 -552 5141 -516
rect 5175 -552 5187 -516
rect 5129 -586 5187 -552
rect 5129 -622 5141 -586
rect 5175 -622 5187 -586
rect 5129 -634 5187 -622
rect 5387 -446 5445 -434
rect 5387 -482 5399 -446
rect 5433 -482 5445 -446
rect 5387 -516 5445 -482
rect 5387 -552 5399 -516
rect 5433 -552 5445 -516
rect 5387 -586 5445 -552
rect 5387 -622 5399 -586
rect 5433 -622 5445 -586
rect 5387 -634 5445 -622
rect 5645 -446 5703 -434
rect 5645 -482 5657 -446
rect 5691 -482 5703 -446
rect 5645 -516 5703 -482
rect 5645 -552 5657 -516
rect 5691 -552 5703 -516
rect 5645 -587 5703 -552
rect 5645 -623 5657 -587
rect 5691 -623 5703 -587
rect 5645 -634 5703 -623
rect 5903 -446 5961 -434
rect 5903 -482 5915 -446
rect 5949 -482 5961 -446
rect 5903 -516 5961 -482
rect 5903 -552 5915 -516
rect 5949 -552 5961 -516
rect 5903 -586 5961 -552
rect 5903 -622 5915 -586
rect 5949 -622 5961 -586
rect 5903 -634 5961 -622
rect 6161 -446 6219 -434
rect 6161 -482 6173 -446
rect 6207 -482 6219 -446
rect 6161 -516 6219 -482
rect 6161 -552 6173 -516
rect 6207 -552 6219 -516
rect 6161 -586 6219 -552
rect 6161 -622 6173 -586
rect 6207 -622 6219 -586
rect 6161 -634 6219 -622
rect 6419 -446 6477 -434
rect 6419 -482 6431 -446
rect 6465 -482 6477 -446
rect 6419 -516 6477 -482
rect 6419 -552 6431 -516
rect 6465 -552 6477 -516
rect 6419 -586 6477 -552
rect 6419 -622 6431 -586
rect 6465 -622 6477 -586
rect 6419 -634 6477 -622
rect 6677 -446 6735 -434
rect 6677 -482 6689 -446
rect 6723 -482 6735 -446
rect 6677 -516 6735 -482
rect 6677 -552 6689 -516
rect 6723 -552 6735 -516
rect 6677 -586 6735 -552
rect 6677 -622 6689 -586
rect 6723 -622 6735 -586
rect 6677 -634 6735 -622
rect 6935 -446 6993 -434
rect 6935 -482 6947 -446
rect 6981 -482 6993 -446
rect 6935 -516 6993 -482
rect 6935 -552 6947 -516
rect 6981 -552 6993 -516
rect 6935 -586 6993 -552
rect 6935 -622 6947 -586
rect 6981 -622 6993 -586
rect 6935 -634 6993 -622
rect 7193 -446 7251 -434
rect 7193 -482 7205 -446
rect 7239 -482 7251 -446
rect 7193 -516 7251 -482
rect 7193 -552 7205 -516
rect 7239 -552 7251 -516
rect 7193 -586 7251 -552
rect 7193 -622 7205 -586
rect 7239 -622 7251 -586
rect 7193 -634 7251 -622
rect 7799 -446 7857 -434
rect 7799 -482 7811 -446
rect 7845 -482 7857 -446
rect 7799 -516 7857 -482
rect 7799 -552 7811 -516
rect 7845 -552 7857 -516
rect 7799 -586 7857 -552
rect 7799 -622 7811 -586
rect 7845 -622 7857 -586
rect 7799 -634 7857 -622
rect 8057 -446 8115 -434
rect 8057 -482 8069 -446
rect 8103 -482 8115 -446
rect 8057 -516 8115 -482
rect 8057 -552 8069 -516
rect 8103 -552 8115 -516
rect 8057 -586 8115 -552
rect 8057 -622 8069 -586
rect 8103 -622 8115 -586
rect 8057 -634 8115 -622
rect 8315 -446 8373 -434
rect 8315 -482 8327 -446
rect 8361 -482 8373 -446
rect 8315 -516 8373 -482
rect 8315 -552 8327 -516
rect 8361 -552 8373 -516
rect 8315 -587 8373 -552
rect 8315 -623 8327 -587
rect 8361 -623 8373 -587
rect 8315 -634 8373 -623
rect 8573 -446 8631 -434
rect 8573 -482 8585 -446
rect 8619 -482 8631 -446
rect 8573 -516 8631 -482
rect 8573 -552 8585 -516
rect 8619 -552 8631 -516
rect 8573 -586 8631 -552
rect 8573 -622 8585 -586
rect 8619 -622 8631 -586
rect 8573 -634 8631 -622
rect 8831 -446 8889 -434
rect 8831 -482 8843 -446
rect 8877 -482 8889 -446
rect 8831 -516 8889 -482
rect 8831 -552 8843 -516
rect 8877 -552 8889 -516
rect 8831 -586 8889 -552
rect 8831 -622 8843 -586
rect 8877 -622 8889 -586
rect 8831 -634 8889 -622
rect 9089 -446 9147 -434
rect 9089 -482 9101 -446
rect 9135 -482 9147 -446
rect 9089 -516 9147 -482
rect 9089 -552 9101 -516
rect 9135 -552 9147 -516
rect 9089 -586 9147 -552
rect 9089 -622 9101 -586
rect 9135 -622 9147 -586
rect 9089 -634 9147 -622
rect 9347 -446 9405 -434
rect 9347 -482 9359 -446
rect 9393 -482 9405 -446
rect 9347 -516 9405 -482
rect 9347 -552 9359 -516
rect 9393 -552 9405 -516
rect 9347 -586 9405 -552
rect 9347 -622 9359 -586
rect 9393 -622 9405 -586
rect 9347 -634 9405 -622
rect 9605 -446 9663 -434
rect 9605 -482 9617 -446
rect 9651 -482 9663 -446
rect 9605 -516 9663 -482
rect 9605 -552 9617 -516
rect 9651 -552 9663 -516
rect 9605 -586 9663 -552
rect 9605 -622 9617 -586
rect 9651 -622 9663 -586
rect 9605 -634 9663 -622
rect 9863 -446 9921 -434
rect 9863 -482 9875 -446
rect 9909 -482 9921 -446
rect 9863 -516 9921 -482
rect 9863 -552 9875 -516
rect 9909 -552 9921 -516
rect 9863 -586 9921 -552
rect 9863 -622 9875 -586
rect 9909 -622 9921 -586
rect 9863 -634 9921 -622
rect 10462 -445 10520 -433
rect 10462 -481 10474 -445
rect 10508 -481 10520 -445
rect 10462 -515 10520 -481
rect 10462 -551 10474 -515
rect 10508 -551 10520 -515
rect 10462 -585 10520 -551
rect 10462 -621 10474 -585
rect 10508 -621 10520 -585
rect 10462 -633 10520 -621
rect 10720 -445 10778 -433
rect 10720 -481 10732 -445
rect 10766 -481 10778 -445
rect 10720 -515 10778 -481
rect 10720 -551 10732 -515
rect 10766 -551 10778 -515
rect 10720 -585 10778 -551
rect 10720 -621 10732 -585
rect 10766 -621 10778 -585
rect 10720 -633 10778 -621
rect 10978 -445 11036 -433
rect 10978 -481 10990 -445
rect 11024 -481 11036 -445
rect 10978 -515 11036 -481
rect 10978 -551 10990 -515
rect 11024 -551 11036 -515
rect 10978 -586 11036 -551
rect 10978 -622 10990 -586
rect 11024 -622 11036 -586
rect 10978 -633 11036 -622
rect 11236 -445 11294 -433
rect 11236 -481 11248 -445
rect 11282 -481 11294 -445
rect 11236 -515 11294 -481
rect 11236 -551 11248 -515
rect 11282 -551 11294 -515
rect 11236 -585 11294 -551
rect 11236 -621 11248 -585
rect 11282 -621 11294 -585
rect 11236 -633 11294 -621
rect 11494 -445 11552 -433
rect 11494 -481 11506 -445
rect 11540 -481 11552 -445
rect 11494 -515 11552 -481
rect 11494 -551 11506 -515
rect 11540 -551 11552 -515
rect 11494 -585 11552 -551
rect 11494 -621 11506 -585
rect 11540 -621 11552 -585
rect 11494 -633 11552 -621
rect 11752 -445 11810 -433
rect 11752 -481 11764 -445
rect 11798 -481 11810 -445
rect 11752 -515 11810 -481
rect 11752 -551 11764 -515
rect 11798 -551 11810 -515
rect 11752 -585 11810 -551
rect 11752 -621 11764 -585
rect 11798 -621 11810 -585
rect 11752 -633 11810 -621
rect 12010 -445 12068 -433
rect 12010 -481 12022 -445
rect 12056 -481 12068 -445
rect 12010 -515 12068 -481
rect 12010 -551 12022 -515
rect 12056 -551 12068 -515
rect 12010 -585 12068 -551
rect 12010 -621 12022 -585
rect 12056 -621 12068 -585
rect 12010 -633 12068 -621
rect 12268 -445 12326 -433
rect 12268 -481 12280 -445
rect 12314 -481 12326 -445
rect 12268 -515 12326 -481
rect 12268 -551 12280 -515
rect 12314 -551 12326 -515
rect 12268 -585 12326 -551
rect 12268 -621 12280 -585
rect 12314 -621 12326 -585
rect 12268 -633 12326 -621
rect 12526 -445 12584 -433
rect 12526 -481 12538 -445
rect 12572 -481 12584 -445
rect 12526 -515 12584 -481
rect 12526 -551 12538 -515
rect 12572 -551 12584 -515
rect 12526 -585 12584 -551
rect 12526 -621 12538 -585
rect 12572 -621 12584 -585
rect 12526 -633 12584 -621
rect 5129 -864 5187 -852
rect 5129 -900 5141 -864
rect 5175 -900 5187 -864
rect 5129 -934 5187 -900
rect 5129 -970 5141 -934
rect 5175 -970 5187 -934
rect 5129 -1004 5187 -970
rect 5129 -1040 5141 -1004
rect 5175 -1040 5187 -1004
rect 5129 -1052 5187 -1040
rect 5387 -864 5445 -852
rect 5387 -900 5399 -864
rect 5433 -900 5445 -864
rect 5387 -934 5445 -900
rect 5387 -970 5399 -934
rect 5433 -970 5445 -934
rect 5387 -1004 5445 -970
rect 5387 -1040 5399 -1004
rect 5433 -1040 5445 -1004
rect 5387 -1052 5445 -1040
rect 5645 -864 5703 -852
rect 5645 -900 5657 -864
rect 5691 -900 5703 -864
rect 5645 -934 5703 -900
rect 5645 -970 5657 -934
rect 5691 -970 5703 -934
rect 5645 -1005 5703 -970
rect 5645 -1041 5657 -1005
rect 5691 -1041 5703 -1005
rect 5645 -1052 5703 -1041
rect 5903 -864 5961 -852
rect 5903 -900 5915 -864
rect 5949 -900 5961 -864
rect 5903 -934 5961 -900
rect 5903 -970 5915 -934
rect 5949 -970 5961 -934
rect 5903 -1004 5961 -970
rect 5903 -1040 5915 -1004
rect 5949 -1040 5961 -1004
rect 5903 -1052 5961 -1040
rect 6161 -864 6219 -852
rect 6161 -900 6173 -864
rect 6207 -900 6219 -864
rect 6161 -934 6219 -900
rect 6161 -970 6173 -934
rect 6207 -970 6219 -934
rect 6161 -1004 6219 -970
rect 6161 -1040 6173 -1004
rect 6207 -1040 6219 -1004
rect 6161 -1052 6219 -1040
rect 6419 -864 6477 -852
rect 6419 -900 6431 -864
rect 6465 -900 6477 -864
rect 6419 -934 6477 -900
rect 6419 -970 6431 -934
rect 6465 -970 6477 -934
rect 6419 -1004 6477 -970
rect 6419 -1040 6431 -1004
rect 6465 -1040 6477 -1004
rect 6419 -1052 6477 -1040
rect 6677 -864 6735 -852
rect 6677 -900 6689 -864
rect 6723 -900 6735 -864
rect 6677 -934 6735 -900
rect 6677 -970 6689 -934
rect 6723 -970 6735 -934
rect 6677 -1004 6735 -970
rect 6677 -1040 6689 -1004
rect 6723 -1040 6735 -1004
rect 6677 -1052 6735 -1040
rect 6935 -864 6993 -852
rect 6935 -900 6947 -864
rect 6981 -900 6993 -864
rect 6935 -934 6993 -900
rect 6935 -970 6947 -934
rect 6981 -970 6993 -934
rect 6935 -1004 6993 -970
rect 6935 -1040 6947 -1004
rect 6981 -1040 6993 -1004
rect 6935 -1052 6993 -1040
rect 7193 -864 7251 -852
rect 7193 -900 7205 -864
rect 7239 -900 7251 -864
rect 7193 -934 7251 -900
rect 7193 -970 7205 -934
rect 7239 -970 7251 -934
rect 7193 -1004 7251 -970
rect 7193 -1040 7205 -1004
rect 7239 -1040 7251 -1004
rect 7193 -1052 7251 -1040
rect 7799 -864 7857 -852
rect 7799 -900 7811 -864
rect 7845 -900 7857 -864
rect 7799 -934 7857 -900
rect 7799 -970 7811 -934
rect 7845 -970 7857 -934
rect 7799 -1004 7857 -970
rect 7799 -1040 7811 -1004
rect 7845 -1040 7857 -1004
rect 7799 -1052 7857 -1040
rect 8057 -864 8115 -852
rect 8057 -900 8069 -864
rect 8103 -900 8115 -864
rect 8057 -934 8115 -900
rect 8057 -970 8069 -934
rect 8103 -970 8115 -934
rect 8057 -1004 8115 -970
rect 8057 -1040 8069 -1004
rect 8103 -1040 8115 -1004
rect 8057 -1052 8115 -1040
rect 8315 -864 8373 -852
rect 8315 -900 8327 -864
rect 8361 -900 8373 -864
rect 8315 -934 8373 -900
rect 8315 -970 8327 -934
rect 8361 -970 8373 -934
rect 8315 -1005 8373 -970
rect 8315 -1041 8327 -1005
rect 8361 -1041 8373 -1005
rect 8315 -1052 8373 -1041
rect 8573 -864 8631 -852
rect 8573 -900 8585 -864
rect 8619 -900 8631 -864
rect 8573 -934 8631 -900
rect 8573 -970 8585 -934
rect 8619 -970 8631 -934
rect 8573 -1004 8631 -970
rect 8573 -1040 8585 -1004
rect 8619 -1040 8631 -1004
rect 8573 -1052 8631 -1040
rect 8831 -864 8889 -852
rect 8831 -900 8843 -864
rect 8877 -900 8889 -864
rect 8831 -934 8889 -900
rect 8831 -970 8843 -934
rect 8877 -970 8889 -934
rect 8831 -1004 8889 -970
rect 8831 -1040 8843 -1004
rect 8877 -1040 8889 -1004
rect 8831 -1052 8889 -1040
rect 9089 -864 9147 -852
rect 9089 -900 9101 -864
rect 9135 -900 9147 -864
rect 9089 -934 9147 -900
rect 9089 -970 9101 -934
rect 9135 -970 9147 -934
rect 9089 -1004 9147 -970
rect 9089 -1040 9101 -1004
rect 9135 -1040 9147 -1004
rect 9089 -1052 9147 -1040
rect 9347 -864 9405 -852
rect 9347 -900 9359 -864
rect 9393 -900 9405 -864
rect 9347 -934 9405 -900
rect 9347 -970 9359 -934
rect 9393 -970 9405 -934
rect 9347 -1004 9405 -970
rect 9347 -1040 9359 -1004
rect 9393 -1040 9405 -1004
rect 9347 -1052 9405 -1040
rect 9605 -864 9663 -852
rect 9605 -900 9617 -864
rect 9651 -900 9663 -864
rect 9605 -934 9663 -900
rect 9605 -970 9617 -934
rect 9651 -970 9663 -934
rect 9605 -1004 9663 -970
rect 9605 -1040 9617 -1004
rect 9651 -1040 9663 -1004
rect 9605 -1052 9663 -1040
rect 9863 -864 9921 -852
rect 9863 -900 9875 -864
rect 9909 -900 9921 -864
rect 9863 -934 9921 -900
rect 9863 -970 9875 -934
rect 9909 -970 9921 -934
rect 9863 -1004 9921 -970
rect 9863 -1040 9875 -1004
rect 9909 -1040 9921 -1004
rect 9863 -1052 9921 -1040
rect 10462 -863 10520 -851
rect 10462 -899 10474 -863
rect 10508 -899 10520 -863
rect 10462 -933 10520 -899
rect 10462 -969 10474 -933
rect 10508 -969 10520 -933
rect 10462 -1003 10520 -969
rect 10462 -1039 10474 -1003
rect 10508 -1039 10520 -1003
rect 10462 -1051 10520 -1039
rect 10720 -863 10778 -851
rect 10720 -899 10732 -863
rect 10766 -899 10778 -863
rect 10720 -933 10778 -899
rect 10720 -969 10732 -933
rect 10766 -969 10778 -933
rect 10720 -1003 10778 -969
rect 10720 -1039 10732 -1003
rect 10766 -1039 10778 -1003
rect 10720 -1051 10778 -1039
rect 10978 -863 11036 -851
rect 10978 -899 10990 -863
rect 11024 -899 11036 -863
rect 10978 -933 11036 -899
rect 10978 -969 10990 -933
rect 11024 -969 11036 -933
rect 10978 -1004 11036 -969
rect 10978 -1040 10990 -1004
rect 11024 -1040 11036 -1004
rect 10978 -1051 11036 -1040
rect 11236 -863 11294 -851
rect 11236 -899 11248 -863
rect 11282 -899 11294 -863
rect 11236 -933 11294 -899
rect 11236 -969 11248 -933
rect 11282 -969 11294 -933
rect 11236 -1003 11294 -969
rect 11236 -1039 11248 -1003
rect 11282 -1039 11294 -1003
rect 11236 -1051 11294 -1039
rect 11494 -863 11552 -851
rect 11494 -899 11506 -863
rect 11540 -899 11552 -863
rect 11494 -933 11552 -899
rect 11494 -969 11506 -933
rect 11540 -969 11552 -933
rect 11494 -1003 11552 -969
rect 11494 -1039 11506 -1003
rect 11540 -1039 11552 -1003
rect 11494 -1051 11552 -1039
rect 11752 -863 11810 -851
rect 11752 -899 11764 -863
rect 11798 -899 11810 -863
rect 11752 -933 11810 -899
rect 11752 -969 11764 -933
rect 11798 -969 11810 -933
rect 11752 -1003 11810 -969
rect 11752 -1039 11764 -1003
rect 11798 -1039 11810 -1003
rect 11752 -1051 11810 -1039
rect 12010 -863 12068 -851
rect 12010 -899 12022 -863
rect 12056 -899 12068 -863
rect 12010 -933 12068 -899
rect 12010 -969 12022 -933
rect 12056 -969 12068 -933
rect 12010 -1003 12068 -969
rect 12010 -1039 12022 -1003
rect 12056 -1039 12068 -1003
rect 12010 -1051 12068 -1039
rect 12268 -863 12326 -851
rect 12268 -899 12280 -863
rect 12314 -899 12326 -863
rect 12268 -933 12326 -899
rect 12268 -969 12280 -933
rect 12314 -969 12326 -933
rect 12268 -1003 12326 -969
rect 12268 -1039 12280 -1003
rect 12314 -1039 12326 -1003
rect 12268 -1051 12326 -1039
rect 12526 -863 12584 -851
rect 12526 -899 12538 -863
rect 12572 -899 12584 -863
rect 12526 -933 12584 -899
rect 12526 -969 12538 -933
rect 12572 -969 12584 -933
rect 12526 -1003 12584 -969
rect 12526 -1039 12538 -1003
rect 12572 -1039 12584 -1003
rect 12526 -1051 12584 -1039
rect 5129 -1282 5187 -1270
rect 5129 -1318 5141 -1282
rect 5175 -1318 5187 -1282
rect 5129 -1352 5187 -1318
rect 5129 -1388 5141 -1352
rect 5175 -1388 5187 -1352
rect 5129 -1422 5187 -1388
rect 5129 -1458 5141 -1422
rect 5175 -1458 5187 -1422
rect 5129 -1470 5187 -1458
rect 5387 -1282 5445 -1270
rect 5387 -1318 5399 -1282
rect 5433 -1318 5445 -1282
rect 5387 -1352 5445 -1318
rect 5387 -1388 5399 -1352
rect 5433 -1388 5445 -1352
rect 5387 -1422 5445 -1388
rect 5387 -1458 5399 -1422
rect 5433 -1458 5445 -1422
rect 5387 -1470 5445 -1458
rect 5645 -1282 5703 -1270
rect 5645 -1318 5657 -1282
rect 5691 -1318 5703 -1282
rect 5645 -1352 5703 -1318
rect 5645 -1388 5657 -1352
rect 5691 -1388 5703 -1352
rect 5645 -1423 5703 -1388
rect 5645 -1459 5657 -1423
rect 5691 -1459 5703 -1423
rect 5645 -1470 5703 -1459
rect 5903 -1282 5961 -1270
rect 5903 -1318 5915 -1282
rect 5949 -1318 5961 -1282
rect 5903 -1352 5961 -1318
rect 5903 -1388 5915 -1352
rect 5949 -1388 5961 -1352
rect 5903 -1422 5961 -1388
rect 5903 -1458 5915 -1422
rect 5949 -1458 5961 -1422
rect 5903 -1470 5961 -1458
rect 6161 -1282 6219 -1270
rect 6161 -1318 6173 -1282
rect 6207 -1318 6219 -1282
rect 6161 -1352 6219 -1318
rect 6161 -1388 6173 -1352
rect 6207 -1388 6219 -1352
rect 6161 -1422 6219 -1388
rect 6161 -1458 6173 -1422
rect 6207 -1458 6219 -1422
rect 6161 -1470 6219 -1458
rect 6419 -1282 6477 -1270
rect 6419 -1318 6431 -1282
rect 6465 -1318 6477 -1282
rect 6419 -1352 6477 -1318
rect 6419 -1388 6431 -1352
rect 6465 -1388 6477 -1352
rect 6419 -1422 6477 -1388
rect 6419 -1458 6431 -1422
rect 6465 -1458 6477 -1422
rect 6419 -1470 6477 -1458
rect 6677 -1282 6735 -1270
rect 6677 -1318 6689 -1282
rect 6723 -1318 6735 -1282
rect 6677 -1352 6735 -1318
rect 6677 -1388 6689 -1352
rect 6723 -1388 6735 -1352
rect 6677 -1422 6735 -1388
rect 6677 -1458 6689 -1422
rect 6723 -1458 6735 -1422
rect 6677 -1470 6735 -1458
rect 6935 -1282 6993 -1270
rect 6935 -1318 6947 -1282
rect 6981 -1318 6993 -1282
rect 6935 -1352 6993 -1318
rect 6935 -1388 6947 -1352
rect 6981 -1388 6993 -1352
rect 6935 -1422 6993 -1388
rect 6935 -1458 6947 -1422
rect 6981 -1458 6993 -1422
rect 6935 -1470 6993 -1458
rect 7193 -1282 7251 -1270
rect 7193 -1318 7205 -1282
rect 7239 -1318 7251 -1282
rect 7193 -1352 7251 -1318
rect 7193 -1388 7205 -1352
rect 7239 -1388 7251 -1352
rect 7193 -1422 7251 -1388
rect 7193 -1458 7205 -1422
rect 7239 -1458 7251 -1422
rect 7193 -1470 7251 -1458
rect 7799 -1282 7857 -1270
rect 7799 -1318 7811 -1282
rect 7845 -1318 7857 -1282
rect 7799 -1352 7857 -1318
rect 7799 -1388 7811 -1352
rect 7845 -1388 7857 -1352
rect 7799 -1422 7857 -1388
rect 7799 -1458 7811 -1422
rect 7845 -1458 7857 -1422
rect 7799 -1470 7857 -1458
rect 8057 -1282 8115 -1270
rect 8057 -1318 8069 -1282
rect 8103 -1318 8115 -1282
rect 8057 -1352 8115 -1318
rect 8057 -1388 8069 -1352
rect 8103 -1388 8115 -1352
rect 8057 -1422 8115 -1388
rect 8057 -1458 8069 -1422
rect 8103 -1458 8115 -1422
rect 8057 -1470 8115 -1458
rect 8315 -1282 8373 -1270
rect 8315 -1318 8327 -1282
rect 8361 -1318 8373 -1282
rect 8315 -1352 8373 -1318
rect 8315 -1388 8327 -1352
rect 8361 -1388 8373 -1352
rect 8315 -1423 8373 -1388
rect 8315 -1459 8327 -1423
rect 8361 -1459 8373 -1423
rect 8315 -1470 8373 -1459
rect 8573 -1282 8631 -1270
rect 8573 -1318 8585 -1282
rect 8619 -1318 8631 -1282
rect 8573 -1352 8631 -1318
rect 8573 -1388 8585 -1352
rect 8619 -1388 8631 -1352
rect 8573 -1422 8631 -1388
rect 8573 -1458 8585 -1422
rect 8619 -1458 8631 -1422
rect 8573 -1470 8631 -1458
rect 8831 -1282 8889 -1270
rect 8831 -1318 8843 -1282
rect 8877 -1318 8889 -1282
rect 8831 -1352 8889 -1318
rect 8831 -1388 8843 -1352
rect 8877 -1388 8889 -1352
rect 8831 -1422 8889 -1388
rect 8831 -1458 8843 -1422
rect 8877 -1458 8889 -1422
rect 8831 -1470 8889 -1458
rect 9089 -1282 9147 -1270
rect 9089 -1318 9101 -1282
rect 9135 -1318 9147 -1282
rect 9089 -1352 9147 -1318
rect 9089 -1388 9101 -1352
rect 9135 -1388 9147 -1352
rect 9089 -1422 9147 -1388
rect 9089 -1458 9101 -1422
rect 9135 -1458 9147 -1422
rect 9089 -1470 9147 -1458
rect 9347 -1282 9405 -1270
rect 9347 -1318 9359 -1282
rect 9393 -1318 9405 -1282
rect 9347 -1352 9405 -1318
rect 9347 -1388 9359 -1352
rect 9393 -1388 9405 -1352
rect 9347 -1422 9405 -1388
rect 9347 -1458 9359 -1422
rect 9393 -1458 9405 -1422
rect 9347 -1470 9405 -1458
rect 9605 -1282 9663 -1270
rect 9605 -1318 9617 -1282
rect 9651 -1318 9663 -1282
rect 9605 -1352 9663 -1318
rect 9605 -1388 9617 -1352
rect 9651 -1388 9663 -1352
rect 9605 -1422 9663 -1388
rect 9605 -1458 9617 -1422
rect 9651 -1458 9663 -1422
rect 9605 -1470 9663 -1458
rect 9863 -1282 9921 -1270
rect 9863 -1318 9875 -1282
rect 9909 -1318 9921 -1282
rect 9863 -1352 9921 -1318
rect 9863 -1388 9875 -1352
rect 9909 -1388 9921 -1352
rect 9863 -1422 9921 -1388
rect 9863 -1458 9875 -1422
rect 9909 -1458 9921 -1422
rect 9863 -1470 9921 -1458
rect 10462 -1281 10520 -1269
rect 10462 -1317 10474 -1281
rect 10508 -1317 10520 -1281
rect 10462 -1351 10520 -1317
rect 10462 -1387 10474 -1351
rect 10508 -1387 10520 -1351
rect 10462 -1421 10520 -1387
rect 10462 -1457 10474 -1421
rect 10508 -1457 10520 -1421
rect 10462 -1469 10520 -1457
rect 10720 -1281 10778 -1269
rect 10720 -1317 10732 -1281
rect 10766 -1317 10778 -1281
rect 10720 -1351 10778 -1317
rect 10720 -1387 10732 -1351
rect 10766 -1387 10778 -1351
rect 10720 -1421 10778 -1387
rect 10720 -1457 10732 -1421
rect 10766 -1457 10778 -1421
rect 10720 -1469 10778 -1457
rect 10978 -1281 11036 -1269
rect 10978 -1317 10990 -1281
rect 11024 -1317 11036 -1281
rect 10978 -1351 11036 -1317
rect 10978 -1387 10990 -1351
rect 11024 -1387 11036 -1351
rect 10978 -1422 11036 -1387
rect 10978 -1458 10990 -1422
rect 11024 -1458 11036 -1422
rect 10978 -1469 11036 -1458
rect 11236 -1281 11294 -1269
rect 11236 -1317 11248 -1281
rect 11282 -1317 11294 -1281
rect 11236 -1351 11294 -1317
rect 11236 -1387 11248 -1351
rect 11282 -1387 11294 -1351
rect 11236 -1421 11294 -1387
rect 11236 -1457 11248 -1421
rect 11282 -1457 11294 -1421
rect 11236 -1469 11294 -1457
rect 11494 -1281 11552 -1269
rect 11494 -1317 11506 -1281
rect 11540 -1317 11552 -1281
rect 11494 -1351 11552 -1317
rect 11494 -1387 11506 -1351
rect 11540 -1387 11552 -1351
rect 11494 -1421 11552 -1387
rect 11494 -1457 11506 -1421
rect 11540 -1457 11552 -1421
rect 11494 -1469 11552 -1457
rect 11752 -1281 11810 -1269
rect 11752 -1317 11764 -1281
rect 11798 -1317 11810 -1281
rect 11752 -1351 11810 -1317
rect 11752 -1387 11764 -1351
rect 11798 -1387 11810 -1351
rect 11752 -1421 11810 -1387
rect 11752 -1457 11764 -1421
rect 11798 -1457 11810 -1421
rect 11752 -1469 11810 -1457
rect 12010 -1281 12068 -1269
rect 12010 -1317 12022 -1281
rect 12056 -1317 12068 -1281
rect 12010 -1351 12068 -1317
rect 12010 -1387 12022 -1351
rect 12056 -1387 12068 -1351
rect 12010 -1421 12068 -1387
rect 12010 -1457 12022 -1421
rect 12056 -1457 12068 -1421
rect 12010 -1469 12068 -1457
rect 12268 -1281 12326 -1269
rect 12268 -1317 12280 -1281
rect 12314 -1317 12326 -1281
rect 12268 -1351 12326 -1317
rect 12268 -1387 12280 -1351
rect 12314 -1387 12326 -1351
rect 12268 -1421 12326 -1387
rect 12268 -1457 12280 -1421
rect 12314 -1457 12326 -1421
rect 12268 -1469 12326 -1457
rect 12526 -1281 12584 -1269
rect 12526 -1317 12538 -1281
rect 12572 -1317 12584 -1281
rect 12526 -1351 12584 -1317
rect 12526 -1387 12538 -1351
rect 12572 -1387 12584 -1351
rect 12526 -1421 12584 -1387
rect 12526 -1457 12538 -1421
rect 12572 -1457 12584 -1421
rect 12526 -1469 12584 -1457
rect 5129 -1700 5187 -1688
rect 5129 -1736 5141 -1700
rect 5175 -1736 5187 -1700
rect 5129 -1770 5187 -1736
rect 5129 -1806 5141 -1770
rect 5175 -1806 5187 -1770
rect 5129 -1840 5187 -1806
rect 5129 -1876 5141 -1840
rect 5175 -1876 5187 -1840
rect 5129 -1888 5187 -1876
rect 5387 -1700 5445 -1688
rect 5387 -1736 5399 -1700
rect 5433 -1736 5445 -1700
rect 5387 -1770 5445 -1736
rect 5387 -1806 5399 -1770
rect 5433 -1806 5445 -1770
rect 5387 -1840 5445 -1806
rect 5387 -1876 5399 -1840
rect 5433 -1876 5445 -1840
rect 5387 -1888 5445 -1876
rect 5645 -1700 5703 -1688
rect 5645 -1736 5657 -1700
rect 5691 -1736 5703 -1700
rect 5645 -1770 5703 -1736
rect 5645 -1806 5657 -1770
rect 5691 -1806 5703 -1770
rect 5645 -1841 5703 -1806
rect 5645 -1877 5657 -1841
rect 5691 -1877 5703 -1841
rect 5645 -1888 5703 -1877
rect 5903 -1700 5961 -1688
rect 5903 -1736 5915 -1700
rect 5949 -1736 5961 -1700
rect 5903 -1770 5961 -1736
rect 5903 -1806 5915 -1770
rect 5949 -1806 5961 -1770
rect 5903 -1840 5961 -1806
rect 5903 -1876 5915 -1840
rect 5949 -1876 5961 -1840
rect 5903 -1888 5961 -1876
rect 6161 -1700 6219 -1688
rect 6161 -1736 6173 -1700
rect 6207 -1736 6219 -1700
rect 6161 -1770 6219 -1736
rect 6161 -1806 6173 -1770
rect 6207 -1806 6219 -1770
rect 6161 -1840 6219 -1806
rect 6161 -1876 6173 -1840
rect 6207 -1876 6219 -1840
rect 6161 -1888 6219 -1876
rect 6419 -1700 6477 -1688
rect 6419 -1736 6431 -1700
rect 6465 -1736 6477 -1700
rect 6419 -1770 6477 -1736
rect 6419 -1806 6431 -1770
rect 6465 -1806 6477 -1770
rect 6419 -1840 6477 -1806
rect 6419 -1876 6431 -1840
rect 6465 -1876 6477 -1840
rect 6419 -1888 6477 -1876
rect 6677 -1700 6735 -1688
rect 6677 -1736 6689 -1700
rect 6723 -1736 6735 -1700
rect 6677 -1770 6735 -1736
rect 6677 -1806 6689 -1770
rect 6723 -1806 6735 -1770
rect 6677 -1840 6735 -1806
rect 6677 -1876 6689 -1840
rect 6723 -1876 6735 -1840
rect 6677 -1888 6735 -1876
rect 6935 -1700 6993 -1688
rect 6935 -1736 6947 -1700
rect 6981 -1736 6993 -1700
rect 6935 -1770 6993 -1736
rect 6935 -1806 6947 -1770
rect 6981 -1806 6993 -1770
rect 6935 -1840 6993 -1806
rect 6935 -1876 6947 -1840
rect 6981 -1876 6993 -1840
rect 6935 -1888 6993 -1876
rect 7193 -1700 7251 -1688
rect 7193 -1736 7205 -1700
rect 7239 -1736 7251 -1700
rect 7193 -1770 7251 -1736
rect 7193 -1806 7205 -1770
rect 7239 -1806 7251 -1770
rect 7193 -1840 7251 -1806
rect 7193 -1876 7205 -1840
rect 7239 -1876 7251 -1840
rect 7193 -1888 7251 -1876
rect 7799 -1700 7857 -1688
rect 7799 -1736 7811 -1700
rect 7845 -1736 7857 -1700
rect 7799 -1770 7857 -1736
rect 7799 -1806 7811 -1770
rect 7845 -1806 7857 -1770
rect 7799 -1840 7857 -1806
rect 7799 -1876 7811 -1840
rect 7845 -1876 7857 -1840
rect 7799 -1888 7857 -1876
rect 8057 -1700 8115 -1688
rect 8057 -1736 8069 -1700
rect 8103 -1736 8115 -1700
rect 8057 -1770 8115 -1736
rect 8057 -1806 8069 -1770
rect 8103 -1806 8115 -1770
rect 8057 -1840 8115 -1806
rect 8057 -1876 8069 -1840
rect 8103 -1876 8115 -1840
rect 8057 -1888 8115 -1876
rect 8315 -1700 8373 -1688
rect 8315 -1736 8327 -1700
rect 8361 -1736 8373 -1700
rect 8315 -1770 8373 -1736
rect 8315 -1806 8327 -1770
rect 8361 -1806 8373 -1770
rect 8315 -1841 8373 -1806
rect 8315 -1877 8327 -1841
rect 8361 -1877 8373 -1841
rect 8315 -1888 8373 -1877
rect 8573 -1700 8631 -1688
rect 8573 -1736 8585 -1700
rect 8619 -1736 8631 -1700
rect 8573 -1770 8631 -1736
rect 8573 -1806 8585 -1770
rect 8619 -1806 8631 -1770
rect 8573 -1840 8631 -1806
rect 8573 -1876 8585 -1840
rect 8619 -1876 8631 -1840
rect 8573 -1888 8631 -1876
rect 8831 -1700 8889 -1688
rect 8831 -1736 8843 -1700
rect 8877 -1736 8889 -1700
rect 8831 -1770 8889 -1736
rect 8831 -1806 8843 -1770
rect 8877 -1806 8889 -1770
rect 8831 -1840 8889 -1806
rect 8831 -1876 8843 -1840
rect 8877 -1876 8889 -1840
rect 8831 -1888 8889 -1876
rect 9089 -1700 9147 -1688
rect 9089 -1736 9101 -1700
rect 9135 -1736 9147 -1700
rect 9089 -1770 9147 -1736
rect 9089 -1806 9101 -1770
rect 9135 -1806 9147 -1770
rect 9089 -1840 9147 -1806
rect 9089 -1876 9101 -1840
rect 9135 -1876 9147 -1840
rect 9089 -1888 9147 -1876
rect 9347 -1700 9405 -1688
rect 9347 -1736 9359 -1700
rect 9393 -1736 9405 -1700
rect 9347 -1770 9405 -1736
rect 9347 -1806 9359 -1770
rect 9393 -1806 9405 -1770
rect 9347 -1840 9405 -1806
rect 9347 -1876 9359 -1840
rect 9393 -1876 9405 -1840
rect 9347 -1888 9405 -1876
rect 9605 -1700 9663 -1688
rect 9605 -1736 9617 -1700
rect 9651 -1736 9663 -1700
rect 9605 -1770 9663 -1736
rect 9605 -1806 9617 -1770
rect 9651 -1806 9663 -1770
rect 9605 -1840 9663 -1806
rect 9605 -1876 9617 -1840
rect 9651 -1876 9663 -1840
rect 9605 -1888 9663 -1876
rect 9863 -1700 9921 -1688
rect 9863 -1736 9875 -1700
rect 9909 -1736 9921 -1700
rect 9863 -1770 9921 -1736
rect 9863 -1806 9875 -1770
rect 9909 -1806 9921 -1770
rect 9863 -1840 9921 -1806
rect 9863 -1876 9875 -1840
rect 9909 -1876 9921 -1840
rect 9863 -1888 9921 -1876
rect 10462 -1699 10520 -1687
rect 10462 -1735 10474 -1699
rect 10508 -1735 10520 -1699
rect 10462 -1769 10520 -1735
rect 10462 -1805 10474 -1769
rect 10508 -1805 10520 -1769
rect 10462 -1839 10520 -1805
rect 10462 -1875 10474 -1839
rect 10508 -1875 10520 -1839
rect 10462 -1887 10520 -1875
rect 10720 -1699 10778 -1687
rect 10720 -1735 10732 -1699
rect 10766 -1735 10778 -1699
rect 10720 -1769 10778 -1735
rect 10720 -1805 10732 -1769
rect 10766 -1805 10778 -1769
rect 10720 -1839 10778 -1805
rect 10720 -1875 10732 -1839
rect 10766 -1875 10778 -1839
rect 10720 -1887 10778 -1875
rect 10978 -1699 11036 -1687
rect 10978 -1735 10990 -1699
rect 11024 -1735 11036 -1699
rect 10978 -1769 11036 -1735
rect 10978 -1805 10990 -1769
rect 11024 -1805 11036 -1769
rect 10978 -1840 11036 -1805
rect 10978 -1876 10990 -1840
rect 11024 -1876 11036 -1840
rect 10978 -1887 11036 -1876
rect 11236 -1699 11294 -1687
rect 11236 -1735 11248 -1699
rect 11282 -1735 11294 -1699
rect 11236 -1769 11294 -1735
rect 11236 -1805 11248 -1769
rect 11282 -1805 11294 -1769
rect 11236 -1839 11294 -1805
rect 11236 -1875 11248 -1839
rect 11282 -1875 11294 -1839
rect 11236 -1887 11294 -1875
rect 11494 -1699 11552 -1687
rect 11494 -1735 11506 -1699
rect 11540 -1735 11552 -1699
rect 11494 -1769 11552 -1735
rect 11494 -1805 11506 -1769
rect 11540 -1805 11552 -1769
rect 11494 -1839 11552 -1805
rect 11494 -1875 11506 -1839
rect 11540 -1875 11552 -1839
rect 11494 -1887 11552 -1875
rect 11752 -1699 11810 -1687
rect 11752 -1735 11764 -1699
rect 11798 -1735 11810 -1699
rect 11752 -1769 11810 -1735
rect 11752 -1805 11764 -1769
rect 11798 -1805 11810 -1769
rect 11752 -1839 11810 -1805
rect 11752 -1875 11764 -1839
rect 11798 -1875 11810 -1839
rect 11752 -1887 11810 -1875
rect 12010 -1699 12068 -1687
rect 12010 -1735 12022 -1699
rect 12056 -1735 12068 -1699
rect 12010 -1769 12068 -1735
rect 12010 -1805 12022 -1769
rect 12056 -1805 12068 -1769
rect 12010 -1839 12068 -1805
rect 12010 -1875 12022 -1839
rect 12056 -1875 12068 -1839
rect 12010 -1887 12068 -1875
rect 12268 -1699 12326 -1687
rect 12268 -1735 12280 -1699
rect 12314 -1735 12326 -1699
rect 12268 -1769 12326 -1735
rect 12268 -1805 12280 -1769
rect 12314 -1805 12326 -1769
rect 12268 -1839 12326 -1805
rect 12268 -1875 12280 -1839
rect 12314 -1875 12326 -1839
rect 12268 -1887 12326 -1875
rect 12526 -1699 12584 -1687
rect 12526 -1735 12538 -1699
rect 12572 -1735 12584 -1699
rect 12526 -1769 12584 -1735
rect 12526 -1805 12538 -1769
rect 12572 -1805 12584 -1769
rect 12526 -1839 12584 -1805
rect 12526 -1875 12538 -1839
rect 12572 -1875 12584 -1839
rect 12526 -1887 12584 -1875
rect 5009 -2354 5067 -2340
rect 5009 -2388 5021 -2354
rect 5055 -2388 5067 -2354
rect 5009 -2422 5067 -2388
rect 5009 -2458 5021 -2422
rect 5055 -2458 5067 -2422
rect 5009 -2492 5067 -2458
rect 5009 -2526 5021 -2492
rect 5055 -2526 5067 -2492
rect 5009 -2540 5067 -2526
rect 5267 -2354 5325 -2340
rect 5267 -2388 5279 -2354
rect 5313 -2388 5325 -2354
rect 5267 -2422 5325 -2388
rect 5267 -2458 5279 -2422
rect 5313 -2458 5325 -2422
rect 5267 -2492 5325 -2458
rect 5267 -2526 5279 -2492
rect 5313 -2526 5325 -2492
rect 5267 -2540 5325 -2526
rect 5549 -2354 5607 -2340
rect 5549 -2388 5561 -2354
rect 5595 -2388 5607 -2354
rect 5549 -2422 5607 -2388
rect 5549 -2458 5561 -2422
rect 5595 -2458 5607 -2422
rect 5549 -2492 5607 -2458
rect 5549 -2526 5561 -2492
rect 5595 -2526 5607 -2492
rect 5549 -2540 5607 -2526
rect 5807 -2354 5865 -2340
rect 5807 -2388 5819 -2354
rect 5853 -2388 5865 -2354
rect 5807 -2422 5865 -2388
rect 5807 -2458 5819 -2422
rect 5853 -2458 5865 -2422
rect 5807 -2492 5865 -2458
rect 5807 -2526 5819 -2492
rect 5853 -2526 5865 -2492
rect 5807 -2540 5865 -2526
rect 6029 -2354 6087 -2340
rect 6029 -2388 6041 -2354
rect 6075 -2388 6087 -2354
rect 6029 -2422 6087 -2388
rect 6029 -2458 6041 -2422
rect 6075 -2458 6087 -2422
rect 6029 -2492 6087 -2458
rect 6029 -2526 6041 -2492
rect 6075 -2526 6087 -2492
rect 6029 -2540 6087 -2526
rect 6287 -2354 6345 -2340
rect 6287 -2388 6299 -2354
rect 6333 -2388 6345 -2354
rect 6287 -2422 6345 -2388
rect 6287 -2458 6299 -2422
rect 6333 -2458 6345 -2422
rect 6287 -2492 6345 -2458
rect 6287 -2526 6299 -2492
rect 6333 -2526 6345 -2492
rect 6287 -2540 6345 -2526
rect 6532 -2352 6590 -2338
rect 6532 -2386 6544 -2352
rect 6578 -2386 6590 -2352
rect 6532 -2420 6590 -2386
rect 6532 -2456 6544 -2420
rect 6578 -2456 6590 -2420
rect 6532 -2490 6590 -2456
rect 6532 -2524 6544 -2490
rect 6578 -2524 6590 -2490
rect 6532 -2538 6590 -2524
rect 6790 -2352 6848 -2338
rect 6790 -2386 6802 -2352
rect 6836 -2386 6848 -2352
rect 6790 -2420 6848 -2386
rect 6790 -2456 6802 -2420
rect 6836 -2456 6848 -2420
rect 6790 -2490 6848 -2456
rect 6790 -2524 6802 -2490
rect 6836 -2524 6848 -2490
rect 6790 -2538 6848 -2524
rect 7042 -2342 7100 -2328
rect 7042 -2376 7054 -2342
rect 7088 -2376 7100 -2342
rect 7042 -2410 7100 -2376
rect 7042 -2446 7054 -2410
rect 7088 -2446 7100 -2410
rect 7042 -2480 7100 -2446
rect 7042 -2514 7054 -2480
rect 7088 -2514 7100 -2480
rect 7042 -2528 7100 -2514
rect 7300 -2342 7358 -2328
rect 7300 -2376 7312 -2342
rect 7346 -2376 7358 -2342
rect 7300 -2410 7358 -2376
rect 7300 -2446 7312 -2410
rect 7346 -2446 7358 -2410
rect 7300 -2480 7358 -2446
rect 7300 -2514 7312 -2480
rect 7346 -2514 7358 -2480
rect 7300 -2528 7358 -2514
rect 7679 -2354 7737 -2340
rect 7679 -2388 7691 -2354
rect 7725 -2388 7737 -2354
rect 7679 -2422 7737 -2388
rect 7679 -2458 7691 -2422
rect 7725 -2458 7737 -2422
rect 7679 -2492 7737 -2458
rect 7679 -2526 7691 -2492
rect 7725 -2526 7737 -2492
rect 7679 -2540 7737 -2526
rect 7937 -2354 7995 -2340
rect 7937 -2388 7949 -2354
rect 7983 -2388 7995 -2354
rect 7937 -2422 7995 -2388
rect 7937 -2458 7949 -2422
rect 7983 -2458 7995 -2422
rect 7937 -2492 7995 -2458
rect 7937 -2526 7949 -2492
rect 7983 -2526 7995 -2492
rect 7937 -2540 7995 -2526
rect 8219 -2354 8277 -2340
rect 8219 -2388 8231 -2354
rect 8265 -2388 8277 -2354
rect 8219 -2422 8277 -2388
rect 8219 -2458 8231 -2422
rect 8265 -2458 8277 -2422
rect 8219 -2492 8277 -2458
rect 8219 -2526 8231 -2492
rect 8265 -2526 8277 -2492
rect 8219 -2540 8277 -2526
rect 8477 -2354 8535 -2340
rect 8477 -2388 8489 -2354
rect 8523 -2388 8535 -2354
rect 8477 -2422 8535 -2388
rect 8477 -2458 8489 -2422
rect 8523 -2458 8535 -2422
rect 8477 -2492 8535 -2458
rect 8477 -2526 8489 -2492
rect 8523 -2526 8535 -2492
rect 8477 -2540 8535 -2526
rect 8699 -2354 8757 -2340
rect 8699 -2388 8711 -2354
rect 8745 -2388 8757 -2354
rect 8699 -2422 8757 -2388
rect 8699 -2458 8711 -2422
rect 8745 -2458 8757 -2422
rect 8699 -2492 8757 -2458
rect 8699 -2526 8711 -2492
rect 8745 -2526 8757 -2492
rect 8699 -2540 8757 -2526
rect 8957 -2354 9015 -2340
rect 8957 -2388 8969 -2354
rect 9003 -2388 9015 -2354
rect 8957 -2422 9015 -2388
rect 8957 -2458 8969 -2422
rect 9003 -2458 9015 -2422
rect 8957 -2492 9015 -2458
rect 8957 -2526 8969 -2492
rect 9003 -2526 9015 -2492
rect 8957 -2540 9015 -2526
rect 9202 -2352 9260 -2338
rect 9202 -2386 9214 -2352
rect 9248 -2386 9260 -2352
rect 9202 -2420 9260 -2386
rect 9202 -2456 9214 -2420
rect 9248 -2456 9260 -2420
rect 9202 -2490 9260 -2456
rect 9202 -2524 9214 -2490
rect 9248 -2524 9260 -2490
rect 9202 -2538 9260 -2524
rect 9460 -2352 9518 -2338
rect 9460 -2386 9472 -2352
rect 9506 -2386 9518 -2352
rect 9460 -2420 9518 -2386
rect 9460 -2456 9472 -2420
rect 9506 -2456 9518 -2420
rect 9460 -2490 9518 -2456
rect 9460 -2524 9472 -2490
rect 9506 -2524 9518 -2490
rect 9460 -2538 9518 -2524
rect 9712 -2342 9770 -2328
rect 9712 -2376 9724 -2342
rect 9758 -2376 9770 -2342
rect 9712 -2410 9770 -2376
rect 9712 -2446 9724 -2410
rect 9758 -2446 9770 -2410
rect 9712 -2480 9770 -2446
rect 9712 -2514 9724 -2480
rect 9758 -2514 9770 -2480
rect 9712 -2528 9770 -2514
rect 9970 -2342 10028 -2328
rect 9970 -2376 9982 -2342
rect 10016 -2376 10028 -2342
rect 9970 -2410 10028 -2376
rect 9970 -2446 9982 -2410
rect 10016 -2446 10028 -2410
rect 9970 -2480 10028 -2446
rect 9970 -2514 9982 -2480
rect 10016 -2514 10028 -2480
rect 9970 -2528 10028 -2514
rect 10342 -2353 10400 -2339
rect 10342 -2387 10354 -2353
rect 10388 -2387 10400 -2353
rect 10342 -2421 10400 -2387
rect 10342 -2457 10354 -2421
rect 10388 -2457 10400 -2421
rect 10342 -2491 10400 -2457
rect 10342 -2525 10354 -2491
rect 10388 -2525 10400 -2491
rect 10342 -2539 10400 -2525
rect 10600 -2353 10658 -2339
rect 10600 -2387 10612 -2353
rect 10646 -2387 10658 -2353
rect 10600 -2421 10658 -2387
rect 10600 -2457 10612 -2421
rect 10646 -2457 10658 -2421
rect 10600 -2491 10658 -2457
rect 10600 -2525 10612 -2491
rect 10646 -2525 10658 -2491
rect 10600 -2539 10658 -2525
rect 10882 -2353 10940 -2339
rect 10882 -2387 10894 -2353
rect 10928 -2387 10940 -2353
rect 10882 -2421 10940 -2387
rect 10882 -2457 10894 -2421
rect 10928 -2457 10940 -2421
rect 10882 -2491 10940 -2457
rect 10882 -2525 10894 -2491
rect 10928 -2525 10940 -2491
rect 10882 -2539 10940 -2525
rect 11140 -2353 11198 -2339
rect 11140 -2387 11152 -2353
rect 11186 -2387 11198 -2353
rect 11140 -2421 11198 -2387
rect 11140 -2457 11152 -2421
rect 11186 -2457 11198 -2421
rect 11140 -2491 11198 -2457
rect 11140 -2525 11152 -2491
rect 11186 -2525 11198 -2491
rect 11140 -2539 11198 -2525
rect 11362 -2353 11420 -2339
rect 11362 -2387 11374 -2353
rect 11408 -2387 11420 -2353
rect 11362 -2421 11420 -2387
rect 11362 -2457 11374 -2421
rect 11408 -2457 11420 -2421
rect 11362 -2491 11420 -2457
rect 11362 -2525 11374 -2491
rect 11408 -2525 11420 -2491
rect 11362 -2539 11420 -2525
rect 11620 -2353 11678 -2339
rect 11620 -2387 11632 -2353
rect 11666 -2387 11678 -2353
rect 11620 -2421 11678 -2387
rect 11620 -2457 11632 -2421
rect 11666 -2457 11678 -2421
rect 11620 -2491 11678 -2457
rect 11620 -2525 11632 -2491
rect 11666 -2525 11678 -2491
rect 11620 -2539 11678 -2525
rect 11865 -2351 11923 -2337
rect 11865 -2385 11877 -2351
rect 11911 -2385 11923 -2351
rect 11865 -2419 11923 -2385
rect 11865 -2455 11877 -2419
rect 11911 -2455 11923 -2419
rect 11865 -2489 11923 -2455
rect 11865 -2523 11877 -2489
rect 11911 -2523 11923 -2489
rect 11865 -2537 11923 -2523
rect 12123 -2351 12181 -2337
rect 12123 -2385 12135 -2351
rect 12169 -2385 12181 -2351
rect 12123 -2419 12181 -2385
rect 12123 -2455 12135 -2419
rect 12169 -2455 12181 -2419
rect 12123 -2489 12181 -2455
rect 12123 -2523 12135 -2489
rect 12169 -2523 12181 -2489
rect 12123 -2537 12181 -2523
rect 12375 -2341 12433 -2327
rect 12375 -2375 12387 -2341
rect 12421 -2375 12433 -2341
rect 12375 -2409 12433 -2375
rect 12375 -2445 12387 -2409
rect 12421 -2445 12433 -2409
rect 12375 -2479 12433 -2445
rect 12375 -2513 12387 -2479
rect 12421 -2513 12433 -2479
rect 12375 -2527 12433 -2513
rect 12633 -2341 12691 -2327
rect 12633 -2375 12645 -2341
rect 12679 -2375 12691 -2341
rect 12633 -2409 12691 -2375
rect 12633 -2445 12645 -2409
rect 12679 -2445 12691 -2409
rect 12633 -2479 12691 -2445
rect 12633 -2513 12645 -2479
rect 12679 -2513 12691 -2479
rect 12633 -2527 12691 -2513
rect 12674 -4248 12732 -4236
rect 12674 -4308 12686 -4248
rect 12720 -4308 12732 -4248
rect 12674 -4320 12732 -4308
rect 12762 -4248 12820 -4236
rect 12762 -4308 12774 -4248
rect 12808 -4308 12820 -4248
rect 12762 -4320 12820 -4308
rect 13064 -4248 13122 -4236
rect 13064 -4308 13076 -4248
rect 13110 -4308 13122 -4248
rect 13064 -4320 13122 -4308
rect 13152 -4248 13210 -4236
rect 13152 -4308 13164 -4248
rect 13198 -4308 13210 -4248
rect 13152 -4320 13210 -4308
rect 5129 -5096 5187 -5084
rect 5129 -5132 5141 -5096
rect 5175 -5132 5187 -5096
rect 5129 -5166 5187 -5132
rect 5129 -5202 5141 -5166
rect 5175 -5202 5187 -5166
rect 5129 -5236 5187 -5202
rect 5129 -5272 5141 -5236
rect 5175 -5272 5187 -5236
rect 5129 -5284 5187 -5272
rect 5387 -5096 5445 -5084
rect 5387 -5132 5399 -5096
rect 5433 -5132 5445 -5096
rect 5387 -5166 5445 -5132
rect 5387 -5202 5399 -5166
rect 5433 -5202 5445 -5166
rect 5387 -5236 5445 -5202
rect 5387 -5272 5399 -5236
rect 5433 -5272 5445 -5236
rect 5387 -5284 5445 -5272
rect 5645 -5096 5703 -5084
rect 5645 -5132 5657 -5096
rect 5691 -5132 5703 -5096
rect 5645 -5166 5703 -5132
rect 5645 -5202 5657 -5166
rect 5691 -5202 5703 -5166
rect 5645 -5237 5703 -5202
rect 5645 -5273 5657 -5237
rect 5691 -5273 5703 -5237
rect 5645 -5284 5703 -5273
rect 5903 -5096 5961 -5084
rect 5903 -5132 5915 -5096
rect 5949 -5132 5961 -5096
rect 5903 -5166 5961 -5132
rect 5903 -5202 5915 -5166
rect 5949 -5202 5961 -5166
rect 5903 -5236 5961 -5202
rect 5903 -5272 5915 -5236
rect 5949 -5272 5961 -5236
rect 5903 -5284 5961 -5272
rect 6161 -5096 6219 -5084
rect 6161 -5132 6173 -5096
rect 6207 -5132 6219 -5096
rect 6161 -5166 6219 -5132
rect 6161 -5202 6173 -5166
rect 6207 -5202 6219 -5166
rect 6161 -5236 6219 -5202
rect 6161 -5272 6173 -5236
rect 6207 -5272 6219 -5236
rect 6161 -5284 6219 -5272
rect 6419 -5096 6477 -5084
rect 6419 -5132 6431 -5096
rect 6465 -5132 6477 -5096
rect 6419 -5166 6477 -5132
rect 6419 -5202 6431 -5166
rect 6465 -5202 6477 -5166
rect 6419 -5236 6477 -5202
rect 6419 -5272 6431 -5236
rect 6465 -5272 6477 -5236
rect 6419 -5284 6477 -5272
rect 6677 -5096 6735 -5084
rect 6677 -5132 6689 -5096
rect 6723 -5132 6735 -5096
rect 6677 -5166 6735 -5132
rect 6677 -5202 6689 -5166
rect 6723 -5202 6735 -5166
rect 6677 -5236 6735 -5202
rect 6677 -5272 6689 -5236
rect 6723 -5272 6735 -5236
rect 6677 -5284 6735 -5272
rect 6935 -5096 6993 -5084
rect 6935 -5132 6947 -5096
rect 6981 -5132 6993 -5096
rect 6935 -5166 6993 -5132
rect 6935 -5202 6947 -5166
rect 6981 -5202 6993 -5166
rect 6935 -5236 6993 -5202
rect 6935 -5272 6947 -5236
rect 6981 -5272 6993 -5236
rect 6935 -5284 6993 -5272
rect 7193 -5096 7251 -5084
rect 7193 -5132 7205 -5096
rect 7239 -5132 7251 -5096
rect 7193 -5166 7251 -5132
rect 7193 -5202 7205 -5166
rect 7239 -5202 7251 -5166
rect 7193 -5236 7251 -5202
rect 7193 -5272 7205 -5236
rect 7239 -5272 7251 -5236
rect 7193 -5284 7251 -5272
rect 7799 -5096 7857 -5084
rect 7799 -5132 7811 -5096
rect 7845 -5132 7857 -5096
rect 7799 -5166 7857 -5132
rect 7799 -5202 7811 -5166
rect 7845 -5202 7857 -5166
rect 7799 -5236 7857 -5202
rect 7799 -5272 7811 -5236
rect 7845 -5272 7857 -5236
rect 7799 -5284 7857 -5272
rect 8057 -5096 8115 -5084
rect 8057 -5132 8069 -5096
rect 8103 -5132 8115 -5096
rect 8057 -5166 8115 -5132
rect 8057 -5202 8069 -5166
rect 8103 -5202 8115 -5166
rect 8057 -5236 8115 -5202
rect 8057 -5272 8069 -5236
rect 8103 -5272 8115 -5236
rect 8057 -5284 8115 -5272
rect 8315 -5096 8373 -5084
rect 8315 -5132 8327 -5096
rect 8361 -5132 8373 -5096
rect 8315 -5166 8373 -5132
rect 8315 -5202 8327 -5166
rect 8361 -5202 8373 -5166
rect 8315 -5237 8373 -5202
rect 8315 -5273 8327 -5237
rect 8361 -5273 8373 -5237
rect 8315 -5284 8373 -5273
rect 8573 -5096 8631 -5084
rect 8573 -5132 8585 -5096
rect 8619 -5132 8631 -5096
rect 8573 -5166 8631 -5132
rect 8573 -5202 8585 -5166
rect 8619 -5202 8631 -5166
rect 8573 -5236 8631 -5202
rect 8573 -5272 8585 -5236
rect 8619 -5272 8631 -5236
rect 8573 -5284 8631 -5272
rect 8831 -5096 8889 -5084
rect 8831 -5132 8843 -5096
rect 8877 -5132 8889 -5096
rect 8831 -5166 8889 -5132
rect 8831 -5202 8843 -5166
rect 8877 -5202 8889 -5166
rect 8831 -5236 8889 -5202
rect 8831 -5272 8843 -5236
rect 8877 -5272 8889 -5236
rect 8831 -5284 8889 -5272
rect 9089 -5096 9147 -5084
rect 9089 -5132 9101 -5096
rect 9135 -5132 9147 -5096
rect 9089 -5166 9147 -5132
rect 9089 -5202 9101 -5166
rect 9135 -5202 9147 -5166
rect 9089 -5236 9147 -5202
rect 9089 -5272 9101 -5236
rect 9135 -5272 9147 -5236
rect 9089 -5284 9147 -5272
rect 9347 -5096 9405 -5084
rect 9347 -5132 9359 -5096
rect 9393 -5132 9405 -5096
rect 9347 -5166 9405 -5132
rect 9347 -5202 9359 -5166
rect 9393 -5202 9405 -5166
rect 9347 -5236 9405 -5202
rect 9347 -5272 9359 -5236
rect 9393 -5272 9405 -5236
rect 9347 -5284 9405 -5272
rect 9605 -5096 9663 -5084
rect 9605 -5132 9617 -5096
rect 9651 -5132 9663 -5096
rect 9605 -5166 9663 -5132
rect 9605 -5202 9617 -5166
rect 9651 -5202 9663 -5166
rect 9605 -5236 9663 -5202
rect 9605 -5272 9617 -5236
rect 9651 -5272 9663 -5236
rect 9605 -5284 9663 -5272
rect 9863 -5096 9921 -5084
rect 9863 -5132 9875 -5096
rect 9909 -5132 9921 -5096
rect 9863 -5166 9921 -5132
rect 9863 -5202 9875 -5166
rect 9909 -5202 9921 -5166
rect 9863 -5236 9921 -5202
rect 9863 -5272 9875 -5236
rect 9909 -5272 9921 -5236
rect 9863 -5284 9921 -5272
rect 10462 -5095 10520 -5083
rect 10462 -5131 10474 -5095
rect 10508 -5131 10520 -5095
rect 10462 -5165 10520 -5131
rect 10462 -5201 10474 -5165
rect 10508 -5201 10520 -5165
rect 10462 -5235 10520 -5201
rect 10462 -5271 10474 -5235
rect 10508 -5271 10520 -5235
rect 10462 -5283 10520 -5271
rect 10720 -5095 10778 -5083
rect 10720 -5131 10732 -5095
rect 10766 -5131 10778 -5095
rect 10720 -5165 10778 -5131
rect 10720 -5201 10732 -5165
rect 10766 -5201 10778 -5165
rect 10720 -5235 10778 -5201
rect 10720 -5271 10732 -5235
rect 10766 -5271 10778 -5235
rect 10720 -5283 10778 -5271
rect 10978 -5095 11036 -5083
rect 10978 -5131 10990 -5095
rect 11024 -5131 11036 -5095
rect 10978 -5165 11036 -5131
rect 10978 -5201 10990 -5165
rect 11024 -5201 11036 -5165
rect 10978 -5236 11036 -5201
rect 10978 -5272 10990 -5236
rect 11024 -5272 11036 -5236
rect 10978 -5283 11036 -5272
rect 11236 -5095 11294 -5083
rect 11236 -5131 11248 -5095
rect 11282 -5131 11294 -5095
rect 11236 -5165 11294 -5131
rect 11236 -5201 11248 -5165
rect 11282 -5201 11294 -5165
rect 11236 -5235 11294 -5201
rect 11236 -5271 11248 -5235
rect 11282 -5271 11294 -5235
rect 11236 -5283 11294 -5271
rect 11494 -5095 11552 -5083
rect 11494 -5131 11506 -5095
rect 11540 -5131 11552 -5095
rect 11494 -5165 11552 -5131
rect 11494 -5201 11506 -5165
rect 11540 -5201 11552 -5165
rect 11494 -5235 11552 -5201
rect 11494 -5271 11506 -5235
rect 11540 -5271 11552 -5235
rect 11494 -5283 11552 -5271
rect 11752 -5095 11810 -5083
rect 11752 -5131 11764 -5095
rect 11798 -5131 11810 -5095
rect 11752 -5165 11810 -5131
rect 11752 -5201 11764 -5165
rect 11798 -5201 11810 -5165
rect 11752 -5235 11810 -5201
rect 11752 -5271 11764 -5235
rect 11798 -5271 11810 -5235
rect 11752 -5283 11810 -5271
rect 12010 -5095 12068 -5083
rect 12010 -5131 12022 -5095
rect 12056 -5131 12068 -5095
rect 12010 -5165 12068 -5131
rect 12010 -5201 12022 -5165
rect 12056 -5201 12068 -5165
rect 12010 -5235 12068 -5201
rect 12010 -5271 12022 -5235
rect 12056 -5271 12068 -5235
rect 12010 -5283 12068 -5271
rect 12268 -5095 12326 -5083
rect 12268 -5131 12280 -5095
rect 12314 -5131 12326 -5095
rect 12268 -5165 12326 -5131
rect 12268 -5201 12280 -5165
rect 12314 -5201 12326 -5165
rect 12268 -5235 12326 -5201
rect 12268 -5271 12280 -5235
rect 12314 -5271 12326 -5235
rect 12268 -5283 12326 -5271
rect 12526 -5095 12584 -5083
rect 12526 -5131 12538 -5095
rect 12572 -5131 12584 -5095
rect 12526 -5165 12584 -5131
rect 12526 -5201 12538 -5165
rect 12572 -5201 12584 -5165
rect 12526 -5235 12584 -5201
rect 12526 -5271 12538 -5235
rect 12572 -5271 12584 -5235
rect 12526 -5283 12584 -5271
rect 5129 -5514 5187 -5502
rect 5129 -5550 5141 -5514
rect 5175 -5550 5187 -5514
rect 5129 -5584 5187 -5550
rect 5129 -5620 5141 -5584
rect 5175 -5620 5187 -5584
rect 5129 -5654 5187 -5620
rect 5129 -5690 5141 -5654
rect 5175 -5690 5187 -5654
rect 5129 -5702 5187 -5690
rect 5387 -5514 5445 -5502
rect 5387 -5550 5399 -5514
rect 5433 -5550 5445 -5514
rect 5387 -5584 5445 -5550
rect 5387 -5620 5399 -5584
rect 5433 -5620 5445 -5584
rect 5387 -5654 5445 -5620
rect 5387 -5690 5399 -5654
rect 5433 -5690 5445 -5654
rect 5387 -5702 5445 -5690
rect 5645 -5514 5703 -5502
rect 5645 -5550 5657 -5514
rect 5691 -5550 5703 -5514
rect 5645 -5584 5703 -5550
rect 5645 -5620 5657 -5584
rect 5691 -5620 5703 -5584
rect 5645 -5655 5703 -5620
rect 5645 -5691 5657 -5655
rect 5691 -5691 5703 -5655
rect 5645 -5702 5703 -5691
rect 5903 -5514 5961 -5502
rect 5903 -5550 5915 -5514
rect 5949 -5550 5961 -5514
rect 5903 -5584 5961 -5550
rect 5903 -5620 5915 -5584
rect 5949 -5620 5961 -5584
rect 5903 -5654 5961 -5620
rect 5903 -5690 5915 -5654
rect 5949 -5690 5961 -5654
rect 5903 -5702 5961 -5690
rect 6161 -5514 6219 -5502
rect 6161 -5550 6173 -5514
rect 6207 -5550 6219 -5514
rect 6161 -5584 6219 -5550
rect 6161 -5620 6173 -5584
rect 6207 -5620 6219 -5584
rect 6161 -5654 6219 -5620
rect 6161 -5690 6173 -5654
rect 6207 -5690 6219 -5654
rect 6161 -5702 6219 -5690
rect 6419 -5514 6477 -5502
rect 6419 -5550 6431 -5514
rect 6465 -5550 6477 -5514
rect 6419 -5584 6477 -5550
rect 6419 -5620 6431 -5584
rect 6465 -5620 6477 -5584
rect 6419 -5654 6477 -5620
rect 6419 -5690 6431 -5654
rect 6465 -5690 6477 -5654
rect 6419 -5702 6477 -5690
rect 6677 -5514 6735 -5502
rect 6677 -5550 6689 -5514
rect 6723 -5550 6735 -5514
rect 6677 -5584 6735 -5550
rect 6677 -5620 6689 -5584
rect 6723 -5620 6735 -5584
rect 6677 -5654 6735 -5620
rect 6677 -5690 6689 -5654
rect 6723 -5690 6735 -5654
rect 6677 -5702 6735 -5690
rect 6935 -5514 6993 -5502
rect 6935 -5550 6947 -5514
rect 6981 -5550 6993 -5514
rect 6935 -5584 6993 -5550
rect 6935 -5620 6947 -5584
rect 6981 -5620 6993 -5584
rect 6935 -5654 6993 -5620
rect 6935 -5690 6947 -5654
rect 6981 -5690 6993 -5654
rect 6935 -5702 6993 -5690
rect 7193 -5514 7251 -5502
rect 7193 -5550 7205 -5514
rect 7239 -5550 7251 -5514
rect 7193 -5584 7251 -5550
rect 7193 -5620 7205 -5584
rect 7239 -5620 7251 -5584
rect 7193 -5654 7251 -5620
rect 7193 -5690 7205 -5654
rect 7239 -5690 7251 -5654
rect 7193 -5702 7251 -5690
rect 7799 -5514 7857 -5502
rect 7799 -5550 7811 -5514
rect 7845 -5550 7857 -5514
rect 7799 -5584 7857 -5550
rect 7799 -5620 7811 -5584
rect 7845 -5620 7857 -5584
rect 7799 -5654 7857 -5620
rect 7799 -5690 7811 -5654
rect 7845 -5690 7857 -5654
rect 7799 -5702 7857 -5690
rect 8057 -5514 8115 -5502
rect 8057 -5550 8069 -5514
rect 8103 -5550 8115 -5514
rect 8057 -5584 8115 -5550
rect 8057 -5620 8069 -5584
rect 8103 -5620 8115 -5584
rect 8057 -5654 8115 -5620
rect 8057 -5690 8069 -5654
rect 8103 -5690 8115 -5654
rect 8057 -5702 8115 -5690
rect 8315 -5514 8373 -5502
rect 8315 -5550 8327 -5514
rect 8361 -5550 8373 -5514
rect 8315 -5584 8373 -5550
rect 8315 -5620 8327 -5584
rect 8361 -5620 8373 -5584
rect 8315 -5655 8373 -5620
rect 8315 -5691 8327 -5655
rect 8361 -5691 8373 -5655
rect 8315 -5702 8373 -5691
rect 8573 -5514 8631 -5502
rect 8573 -5550 8585 -5514
rect 8619 -5550 8631 -5514
rect 8573 -5584 8631 -5550
rect 8573 -5620 8585 -5584
rect 8619 -5620 8631 -5584
rect 8573 -5654 8631 -5620
rect 8573 -5690 8585 -5654
rect 8619 -5690 8631 -5654
rect 8573 -5702 8631 -5690
rect 8831 -5514 8889 -5502
rect 8831 -5550 8843 -5514
rect 8877 -5550 8889 -5514
rect 8831 -5584 8889 -5550
rect 8831 -5620 8843 -5584
rect 8877 -5620 8889 -5584
rect 8831 -5654 8889 -5620
rect 8831 -5690 8843 -5654
rect 8877 -5690 8889 -5654
rect 8831 -5702 8889 -5690
rect 9089 -5514 9147 -5502
rect 9089 -5550 9101 -5514
rect 9135 -5550 9147 -5514
rect 9089 -5584 9147 -5550
rect 9089 -5620 9101 -5584
rect 9135 -5620 9147 -5584
rect 9089 -5654 9147 -5620
rect 9089 -5690 9101 -5654
rect 9135 -5690 9147 -5654
rect 9089 -5702 9147 -5690
rect 9347 -5514 9405 -5502
rect 9347 -5550 9359 -5514
rect 9393 -5550 9405 -5514
rect 9347 -5584 9405 -5550
rect 9347 -5620 9359 -5584
rect 9393 -5620 9405 -5584
rect 9347 -5654 9405 -5620
rect 9347 -5690 9359 -5654
rect 9393 -5690 9405 -5654
rect 9347 -5702 9405 -5690
rect 9605 -5514 9663 -5502
rect 9605 -5550 9617 -5514
rect 9651 -5550 9663 -5514
rect 9605 -5584 9663 -5550
rect 9605 -5620 9617 -5584
rect 9651 -5620 9663 -5584
rect 9605 -5654 9663 -5620
rect 9605 -5690 9617 -5654
rect 9651 -5690 9663 -5654
rect 9605 -5702 9663 -5690
rect 9863 -5514 9921 -5502
rect 9863 -5550 9875 -5514
rect 9909 -5550 9921 -5514
rect 9863 -5584 9921 -5550
rect 9863 -5620 9875 -5584
rect 9909 -5620 9921 -5584
rect 9863 -5654 9921 -5620
rect 9863 -5690 9875 -5654
rect 9909 -5690 9921 -5654
rect 9863 -5702 9921 -5690
rect 10462 -5513 10520 -5501
rect 10462 -5549 10474 -5513
rect 10508 -5549 10520 -5513
rect 10462 -5583 10520 -5549
rect 10462 -5619 10474 -5583
rect 10508 -5619 10520 -5583
rect 10462 -5653 10520 -5619
rect 10462 -5689 10474 -5653
rect 10508 -5689 10520 -5653
rect 10462 -5701 10520 -5689
rect 10720 -5513 10778 -5501
rect 10720 -5549 10732 -5513
rect 10766 -5549 10778 -5513
rect 10720 -5583 10778 -5549
rect 10720 -5619 10732 -5583
rect 10766 -5619 10778 -5583
rect 10720 -5653 10778 -5619
rect 10720 -5689 10732 -5653
rect 10766 -5689 10778 -5653
rect 10720 -5701 10778 -5689
rect 10978 -5513 11036 -5501
rect 10978 -5549 10990 -5513
rect 11024 -5549 11036 -5513
rect 10978 -5583 11036 -5549
rect 10978 -5619 10990 -5583
rect 11024 -5619 11036 -5583
rect 10978 -5654 11036 -5619
rect 10978 -5690 10990 -5654
rect 11024 -5690 11036 -5654
rect 10978 -5701 11036 -5690
rect 11236 -5513 11294 -5501
rect 11236 -5549 11248 -5513
rect 11282 -5549 11294 -5513
rect 11236 -5583 11294 -5549
rect 11236 -5619 11248 -5583
rect 11282 -5619 11294 -5583
rect 11236 -5653 11294 -5619
rect 11236 -5689 11248 -5653
rect 11282 -5689 11294 -5653
rect 11236 -5701 11294 -5689
rect 11494 -5513 11552 -5501
rect 11494 -5549 11506 -5513
rect 11540 -5549 11552 -5513
rect 11494 -5583 11552 -5549
rect 11494 -5619 11506 -5583
rect 11540 -5619 11552 -5583
rect 11494 -5653 11552 -5619
rect 11494 -5689 11506 -5653
rect 11540 -5689 11552 -5653
rect 11494 -5701 11552 -5689
rect 11752 -5513 11810 -5501
rect 11752 -5549 11764 -5513
rect 11798 -5549 11810 -5513
rect 11752 -5583 11810 -5549
rect 11752 -5619 11764 -5583
rect 11798 -5619 11810 -5583
rect 11752 -5653 11810 -5619
rect 11752 -5689 11764 -5653
rect 11798 -5689 11810 -5653
rect 11752 -5701 11810 -5689
rect 12010 -5513 12068 -5501
rect 12010 -5549 12022 -5513
rect 12056 -5549 12068 -5513
rect 12010 -5583 12068 -5549
rect 12010 -5619 12022 -5583
rect 12056 -5619 12068 -5583
rect 12010 -5653 12068 -5619
rect 12010 -5689 12022 -5653
rect 12056 -5689 12068 -5653
rect 12010 -5701 12068 -5689
rect 12268 -5513 12326 -5501
rect 12268 -5549 12280 -5513
rect 12314 -5549 12326 -5513
rect 12268 -5583 12326 -5549
rect 12268 -5619 12280 -5583
rect 12314 -5619 12326 -5583
rect 12268 -5653 12326 -5619
rect 12268 -5689 12280 -5653
rect 12314 -5689 12326 -5653
rect 12268 -5701 12326 -5689
rect 12526 -5513 12584 -5501
rect 12526 -5549 12538 -5513
rect 12572 -5549 12584 -5513
rect 12526 -5583 12584 -5549
rect 12526 -5619 12538 -5583
rect 12572 -5619 12584 -5583
rect 12526 -5653 12584 -5619
rect 12526 -5689 12538 -5653
rect 12572 -5689 12584 -5653
rect 12526 -5701 12584 -5689
rect 5129 -5932 5187 -5920
rect 5129 -5968 5141 -5932
rect 5175 -5968 5187 -5932
rect 5129 -6002 5187 -5968
rect 5129 -6038 5141 -6002
rect 5175 -6038 5187 -6002
rect 5129 -6072 5187 -6038
rect 5129 -6108 5141 -6072
rect 5175 -6108 5187 -6072
rect 5129 -6120 5187 -6108
rect 5387 -5932 5445 -5920
rect 5387 -5968 5399 -5932
rect 5433 -5968 5445 -5932
rect 5387 -6002 5445 -5968
rect 5387 -6038 5399 -6002
rect 5433 -6038 5445 -6002
rect 5387 -6072 5445 -6038
rect 5387 -6108 5399 -6072
rect 5433 -6108 5445 -6072
rect 5387 -6120 5445 -6108
rect 5645 -5932 5703 -5920
rect 5645 -5968 5657 -5932
rect 5691 -5968 5703 -5932
rect 5645 -6002 5703 -5968
rect 5645 -6038 5657 -6002
rect 5691 -6038 5703 -6002
rect 5645 -6073 5703 -6038
rect 5645 -6109 5657 -6073
rect 5691 -6109 5703 -6073
rect 5645 -6120 5703 -6109
rect 5903 -5932 5961 -5920
rect 5903 -5968 5915 -5932
rect 5949 -5968 5961 -5932
rect 5903 -6002 5961 -5968
rect 5903 -6038 5915 -6002
rect 5949 -6038 5961 -6002
rect 5903 -6072 5961 -6038
rect 5903 -6108 5915 -6072
rect 5949 -6108 5961 -6072
rect 5903 -6120 5961 -6108
rect 6161 -5932 6219 -5920
rect 6161 -5968 6173 -5932
rect 6207 -5968 6219 -5932
rect 6161 -6002 6219 -5968
rect 6161 -6038 6173 -6002
rect 6207 -6038 6219 -6002
rect 6161 -6072 6219 -6038
rect 6161 -6108 6173 -6072
rect 6207 -6108 6219 -6072
rect 6161 -6120 6219 -6108
rect 6419 -5932 6477 -5920
rect 6419 -5968 6431 -5932
rect 6465 -5968 6477 -5932
rect 6419 -6002 6477 -5968
rect 6419 -6038 6431 -6002
rect 6465 -6038 6477 -6002
rect 6419 -6072 6477 -6038
rect 6419 -6108 6431 -6072
rect 6465 -6108 6477 -6072
rect 6419 -6120 6477 -6108
rect 6677 -5932 6735 -5920
rect 6677 -5968 6689 -5932
rect 6723 -5968 6735 -5932
rect 6677 -6002 6735 -5968
rect 6677 -6038 6689 -6002
rect 6723 -6038 6735 -6002
rect 6677 -6072 6735 -6038
rect 6677 -6108 6689 -6072
rect 6723 -6108 6735 -6072
rect 6677 -6120 6735 -6108
rect 6935 -5932 6993 -5920
rect 6935 -5968 6947 -5932
rect 6981 -5968 6993 -5932
rect 6935 -6002 6993 -5968
rect 6935 -6038 6947 -6002
rect 6981 -6038 6993 -6002
rect 6935 -6072 6993 -6038
rect 6935 -6108 6947 -6072
rect 6981 -6108 6993 -6072
rect 6935 -6120 6993 -6108
rect 7193 -5932 7251 -5920
rect 7193 -5968 7205 -5932
rect 7239 -5968 7251 -5932
rect 7193 -6002 7251 -5968
rect 7193 -6038 7205 -6002
rect 7239 -6038 7251 -6002
rect 7193 -6072 7251 -6038
rect 7193 -6108 7205 -6072
rect 7239 -6108 7251 -6072
rect 7193 -6120 7251 -6108
rect 7799 -5932 7857 -5920
rect 7799 -5968 7811 -5932
rect 7845 -5968 7857 -5932
rect 7799 -6002 7857 -5968
rect 7799 -6038 7811 -6002
rect 7845 -6038 7857 -6002
rect 7799 -6072 7857 -6038
rect 7799 -6108 7811 -6072
rect 7845 -6108 7857 -6072
rect 7799 -6120 7857 -6108
rect 8057 -5932 8115 -5920
rect 8057 -5968 8069 -5932
rect 8103 -5968 8115 -5932
rect 8057 -6002 8115 -5968
rect 8057 -6038 8069 -6002
rect 8103 -6038 8115 -6002
rect 8057 -6072 8115 -6038
rect 8057 -6108 8069 -6072
rect 8103 -6108 8115 -6072
rect 8057 -6120 8115 -6108
rect 8315 -5932 8373 -5920
rect 8315 -5968 8327 -5932
rect 8361 -5968 8373 -5932
rect 8315 -6002 8373 -5968
rect 8315 -6038 8327 -6002
rect 8361 -6038 8373 -6002
rect 8315 -6073 8373 -6038
rect 8315 -6109 8327 -6073
rect 8361 -6109 8373 -6073
rect 8315 -6120 8373 -6109
rect 8573 -5932 8631 -5920
rect 8573 -5968 8585 -5932
rect 8619 -5968 8631 -5932
rect 8573 -6002 8631 -5968
rect 8573 -6038 8585 -6002
rect 8619 -6038 8631 -6002
rect 8573 -6072 8631 -6038
rect 8573 -6108 8585 -6072
rect 8619 -6108 8631 -6072
rect 8573 -6120 8631 -6108
rect 8831 -5932 8889 -5920
rect 8831 -5968 8843 -5932
rect 8877 -5968 8889 -5932
rect 8831 -6002 8889 -5968
rect 8831 -6038 8843 -6002
rect 8877 -6038 8889 -6002
rect 8831 -6072 8889 -6038
rect 8831 -6108 8843 -6072
rect 8877 -6108 8889 -6072
rect 8831 -6120 8889 -6108
rect 9089 -5932 9147 -5920
rect 9089 -5968 9101 -5932
rect 9135 -5968 9147 -5932
rect 9089 -6002 9147 -5968
rect 9089 -6038 9101 -6002
rect 9135 -6038 9147 -6002
rect 9089 -6072 9147 -6038
rect 9089 -6108 9101 -6072
rect 9135 -6108 9147 -6072
rect 9089 -6120 9147 -6108
rect 9347 -5932 9405 -5920
rect 9347 -5968 9359 -5932
rect 9393 -5968 9405 -5932
rect 9347 -6002 9405 -5968
rect 9347 -6038 9359 -6002
rect 9393 -6038 9405 -6002
rect 9347 -6072 9405 -6038
rect 9347 -6108 9359 -6072
rect 9393 -6108 9405 -6072
rect 9347 -6120 9405 -6108
rect 9605 -5932 9663 -5920
rect 9605 -5968 9617 -5932
rect 9651 -5968 9663 -5932
rect 9605 -6002 9663 -5968
rect 9605 -6038 9617 -6002
rect 9651 -6038 9663 -6002
rect 9605 -6072 9663 -6038
rect 9605 -6108 9617 -6072
rect 9651 -6108 9663 -6072
rect 9605 -6120 9663 -6108
rect 9863 -5932 9921 -5920
rect 9863 -5968 9875 -5932
rect 9909 -5968 9921 -5932
rect 9863 -6002 9921 -5968
rect 9863 -6038 9875 -6002
rect 9909 -6038 9921 -6002
rect 9863 -6072 9921 -6038
rect 9863 -6108 9875 -6072
rect 9909 -6108 9921 -6072
rect 9863 -6120 9921 -6108
rect 10462 -5931 10520 -5919
rect 10462 -5967 10474 -5931
rect 10508 -5967 10520 -5931
rect 10462 -6001 10520 -5967
rect 10462 -6037 10474 -6001
rect 10508 -6037 10520 -6001
rect 10462 -6071 10520 -6037
rect 10462 -6107 10474 -6071
rect 10508 -6107 10520 -6071
rect 10462 -6119 10520 -6107
rect 10720 -5931 10778 -5919
rect 10720 -5967 10732 -5931
rect 10766 -5967 10778 -5931
rect 10720 -6001 10778 -5967
rect 10720 -6037 10732 -6001
rect 10766 -6037 10778 -6001
rect 10720 -6071 10778 -6037
rect 10720 -6107 10732 -6071
rect 10766 -6107 10778 -6071
rect 10720 -6119 10778 -6107
rect 10978 -5931 11036 -5919
rect 10978 -5967 10990 -5931
rect 11024 -5967 11036 -5931
rect 10978 -6001 11036 -5967
rect 10978 -6037 10990 -6001
rect 11024 -6037 11036 -6001
rect 10978 -6072 11036 -6037
rect 10978 -6108 10990 -6072
rect 11024 -6108 11036 -6072
rect 10978 -6119 11036 -6108
rect 11236 -5931 11294 -5919
rect 11236 -5967 11248 -5931
rect 11282 -5967 11294 -5931
rect 11236 -6001 11294 -5967
rect 11236 -6037 11248 -6001
rect 11282 -6037 11294 -6001
rect 11236 -6071 11294 -6037
rect 11236 -6107 11248 -6071
rect 11282 -6107 11294 -6071
rect 11236 -6119 11294 -6107
rect 11494 -5931 11552 -5919
rect 11494 -5967 11506 -5931
rect 11540 -5967 11552 -5931
rect 11494 -6001 11552 -5967
rect 11494 -6037 11506 -6001
rect 11540 -6037 11552 -6001
rect 11494 -6071 11552 -6037
rect 11494 -6107 11506 -6071
rect 11540 -6107 11552 -6071
rect 11494 -6119 11552 -6107
rect 11752 -5931 11810 -5919
rect 11752 -5967 11764 -5931
rect 11798 -5967 11810 -5931
rect 11752 -6001 11810 -5967
rect 11752 -6037 11764 -6001
rect 11798 -6037 11810 -6001
rect 11752 -6071 11810 -6037
rect 11752 -6107 11764 -6071
rect 11798 -6107 11810 -6071
rect 11752 -6119 11810 -6107
rect 12010 -5931 12068 -5919
rect 12010 -5967 12022 -5931
rect 12056 -5967 12068 -5931
rect 12010 -6001 12068 -5967
rect 12010 -6037 12022 -6001
rect 12056 -6037 12068 -6001
rect 12010 -6071 12068 -6037
rect 12010 -6107 12022 -6071
rect 12056 -6107 12068 -6071
rect 12010 -6119 12068 -6107
rect 12268 -5931 12326 -5919
rect 12268 -5967 12280 -5931
rect 12314 -5967 12326 -5931
rect 12268 -6001 12326 -5967
rect 12268 -6037 12280 -6001
rect 12314 -6037 12326 -6001
rect 12268 -6071 12326 -6037
rect 12268 -6107 12280 -6071
rect 12314 -6107 12326 -6071
rect 12268 -6119 12326 -6107
rect 12526 -5931 12584 -5919
rect 12526 -5967 12538 -5931
rect 12572 -5967 12584 -5931
rect 12526 -6001 12584 -5967
rect 12526 -6037 12538 -6001
rect 12572 -6037 12584 -6001
rect 12526 -6071 12584 -6037
rect 12526 -6107 12538 -6071
rect 12572 -6107 12584 -6071
rect 12526 -6119 12584 -6107
rect 5129 -6350 5187 -6338
rect 5129 -6386 5141 -6350
rect 5175 -6386 5187 -6350
rect 5129 -6420 5187 -6386
rect 5129 -6456 5141 -6420
rect 5175 -6456 5187 -6420
rect 5129 -6490 5187 -6456
rect 5129 -6526 5141 -6490
rect 5175 -6526 5187 -6490
rect 5129 -6538 5187 -6526
rect 5387 -6350 5445 -6338
rect 5387 -6386 5399 -6350
rect 5433 -6386 5445 -6350
rect 5387 -6420 5445 -6386
rect 5387 -6456 5399 -6420
rect 5433 -6456 5445 -6420
rect 5387 -6490 5445 -6456
rect 5387 -6526 5399 -6490
rect 5433 -6526 5445 -6490
rect 5387 -6538 5445 -6526
rect 5645 -6350 5703 -6338
rect 5645 -6386 5657 -6350
rect 5691 -6386 5703 -6350
rect 5645 -6420 5703 -6386
rect 5645 -6456 5657 -6420
rect 5691 -6456 5703 -6420
rect 5645 -6491 5703 -6456
rect 5645 -6527 5657 -6491
rect 5691 -6527 5703 -6491
rect 5645 -6538 5703 -6527
rect 5903 -6350 5961 -6338
rect 5903 -6386 5915 -6350
rect 5949 -6386 5961 -6350
rect 5903 -6420 5961 -6386
rect 5903 -6456 5915 -6420
rect 5949 -6456 5961 -6420
rect 5903 -6490 5961 -6456
rect 5903 -6526 5915 -6490
rect 5949 -6526 5961 -6490
rect 5903 -6538 5961 -6526
rect 6161 -6350 6219 -6338
rect 6161 -6386 6173 -6350
rect 6207 -6386 6219 -6350
rect 6161 -6420 6219 -6386
rect 6161 -6456 6173 -6420
rect 6207 -6456 6219 -6420
rect 6161 -6490 6219 -6456
rect 6161 -6526 6173 -6490
rect 6207 -6526 6219 -6490
rect 6161 -6538 6219 -6526
rect 6419 -6350 6477 -6338
rect 6419 -6386 6431 -6350
rect 6465 -6386 6477 -6350
rect 6419 -6420 6477 -6386
rect 6419 -6456 6431 -6420
rect 6465 -6456 6477 -6420
rect 6419 -6490 6477 -6456
rect 6419 -6526 6431 -6490
rect 6465 -6526 6477 -6490
rect 6419 -6538 6477 -6526
rect 6677 -6350 6735 -6338
rect 6677 -6386 6689 -6350
rect 6723 -6386 6735 -6350
rect 6677 -6420 6735 -6386
rect 6677 -6456 6689 -6420
rect 6723 -6456 6735 -6420
rect 6677 -6490 6735 -6456
rect 6677 -6526 6689 -6490
rect 6723 -6526 6735 -6490
rect 6677 -6538 6735 -6526
rect 6935 -6350 6993 -6338
rect 6935 -6386 6947 -6350
rect 6981 -6386 6993 -6350
rect 6935 -6420 6993 -6386
rect 6935 -6456 6947 -6420
rect 6981 -6456 6993 -6420
rect 6935 -6490 6993 -6456
rect 6935 -6526 6947 -6490
rect 6981 -6526 6993 -6490
rect 6935 -6538 6993 -6526
rect 7193 -6350 7251 -6338
rect 7193 -6386 7205 -6350
rect 7239 -6386 7251 -6350
rect 7193 -6420 7251 -6386
rect 7193 -6456 7205 -6420
rect 7239 -6456 7251 -6420
rect 7193 -6490 7251 -6456
rect 7193 -6526 7205 -6490
rect 7239 -6526 7251 -6490
rect 7193 -6538 7251 -6526
rect 7799 -6350 7857 -6338
rect 7799 -6386 7811 -6350
rect 7845 -6386 7857 -6350
rect 7799 -6420 7857 -6386
rect 7799 -6456 7811 -6420
rect 7845 -6456 7857 -6420
rect 7799 -6490 7857 -6456
rect 7799 -6526 7811 -6490
rect 7845 -6526 7857 -6490
rect 7799 -6538 7857 -6526
rect 8057 -6350 8115 -6338
rect 8057 -6386 8069 -6350
rect 8103 -6386 8115 -6350
rect 8057 -6420 8115 -6386
rect 8057 -6456 8069 -6420
rect 8103 -6456 8115 -6420
rect 8057 -6490 8115 -6456
rect 8057 -6526 8069 -6490
rect 8103 -6526 8115 -6490
rect 8057 -6538 8115 -6526
rect 8315 -6350 8373 -6338
rect 8315 -6386 8327 -6350
rect 8361 -6386 8373 -6350
rect 8315 -6420 8373 -6386
rect 8315 -6456 8327 -6420
rect 8361 -6456 8373 -6420
rect 8315 -6491 8373 -6456
rect 8315 -6527 8327 -6491
rect 8361 -6527 8373 -6491
rect 8315 -6538 8373 -6527
rect 8573 -6350 8631 -6338
rect 8573 -6386 8585 -6350
rect 8619 -6386 8631 -6350
rect 8573 -6420 8631 -6386
rect 8573 -6456 8585 -6420
rect 8619 -6456 8631 -6420
rect 8573 -6490 8631 -6456
rect 8573 -6526 8585 -6490
rect 8619 -6526 8631 -6490
rect 8573 -6538 8631 -6526
rect 8831 -6350 8889 -6338
rect 8831 -6386 8843 -6350
rect 8877 -6386 8889 -6350
rect 8831 -6420 8889 -6386
rect 8831 -6456 8843 -6420
rect 8877 -6456 8889 -6420
rect 8831 -6490 8889 -6456
rect 8831 -6526 8843 -6490
rect 8877 -6526 8889 -6490
rect 8831 -6538 8889 -6526
rect 9089 -6350 9147 -6338
rect 9089 -6386 9101 -6350
rect 9135 -6386 9147 -6350
rect 9089 -6420 9147 -6386
rect 9089 -6456 9101 -6420
rect 9135 -6456 9147 -6420
rect 9089 -6490 9147 -6456
rect 9089 -6526 9101 -6490
rect 9135 -6526 9147 -6490
rect 9089 -6538 9147 -6526
rect 9347 -6350 9405 -6338
rect 9347 -6386 9359 -6350
rect 9393 -6386 9405 -6350
rect 9347 -6420 9405 -6386
rect 9347 -6456 9359 -6420
rect 9393 -6456 9405 -6420
rect 9347 -6490 9405 -6456
rect 9347 -6526 9359 -6490
rect 9393 -6526 9405 -6490
rect 9347 -6538 9405 -6526
rect 9605 -6350 9663 -6338
rect 9605 -6386 9617 -6350
rect 9651 -6386 9663 -6350
rect 9605 -6420 9663 -6386
rect 9605 -6456 9617 -6420
rect 9651 -6456 9663 -6420
rect 9605 -6490 9663 -6456
rect 9605 -6526 9617 -6490
rect 9651 -6526 9663 -6490
rect 9605 -6538 9663 -6526
rect 9863 -6350 9921 -6338
rect 9863 -6386 9875 -6350
rect 9909 -6386 9921 -6350
rect 9863 -6420 9921 -6386
rect 9863 -6456 9875 -6420
rect 9909 -6456 9921 -6420
rect 9863 -6490 9921 -6456
rect 9863 -6526 9875 -6490
rect 9909 -6526 9921 -6490
rect 9863 -6538 9921 -6526
rect 10462 -6349 10520 -6337
rect 10462 -6385 10474 -6349
rect 10508 -6385 10520 -6349
rect 10462 -6419 10520 -6385
rect 10462 -6455 10474 -6419
rect 10508 -6455 10520 -6419
rect 10462 -6489 10520 -6455
rect 10462 -6525 10474 -6489
rect 10508 -6525 10520 -6489
rect 10462 -6537 10520 -6525
rect 10720 -6349 10778 -6337
rect 10720 -6385 10732 -6349
rect 10766 -6385 10778 -6349
rect 10720 -6419 10778 -6385
rect 10720 -6455 10732 -6419
rect 10766 -6455 10778 -6419
rect 10720 -6489 10778 -6455
rect 10720 -6525 10732 -6489
rect 10766 -6525 10778 -6489
rect 10720 -6537 10778 -6525
rect 10978 -6349 11036 -6337
rect 10978 -6385 10990 -6349
rect 11024 -6385 11036 -6349
rect 10978 -6419 11036 -6385
rect 10978 -6455 10990 -6419
rect 11024 -6455 11036 -6419
rect 10978 -6490 11036 -6455
rect 10978 -6526 10990 -6490
rect 11024 -6526 11036 -6490
rect 10978 -6537 11036 -6526
rect 11236 -6349 11294 -6337
rect 11236 -6385 11248 -6349
rect 11282 -6385 11294 -6349
rect 11236 -6419 11294 -6385
rect 11236 -6455 11248 -6419
rect 11282 -6455 11294 -6419
rect 11236 -6489 11294 -6455
rect 11236 -6525 11248 -6489
rect 11282 -6525 11294 -6489
rect 11236 -6537 11294 -6525
rect 11494 -6349 11552 -6337
rect 11494 -6385 11506 -6349
rect 11540 -6385 11552 -6349
rect 11494 -6419 11552 -6385
rect 11494 -6455 11506 -6419
rect 11540 -6455 11552 -6419
rect 11494 -6489 11552 -6455
rect 11494 -6525 11506 -6489
rect 11540 -6525 11552 -6489
rect 11494 -6537 11552 -6525
rect 11752 -6349 11810 -6337
rect 11752 -6385 11764 -6349
rect 11798 -6385 11810 -6349
rect 11752 -6419 11810 -6385
rect 11752 -6455 11764 -6419
rect 11798 -6455 11810 -6419
rect 11752 -6489 11810 -6455
rect 11752 -6525 11764 -6489
rect 11798 -6525 11810 -6489
rect 11752 -6537 11810 -6525
rect 12010 -6349 12068 -6337
rect 12010 -6385 12022 -6349
rect 12056 -6385 12068 -6349
rect 12010 -6419 12068 -6385
rect 12010 -6455 12022 -6419
rect 12056 -6455 12068 -6419
rect 12010 -6489 12068 -6455
rect 12010 -6525 12022 -6489
rect 12056 -6525 12068 -6489
rect 12010 -6537 12068 -6525
rect 12268 -6349 12326 -6337
rect 12268 -6385 12280 -6349
rect 12314 -6385 12326 -6349
rect 12268 -6419 12326 -6385
rect 12268 -6455 12280 -6419
rect 12314 -6455 12326 -6419
rect 12268 -6489 12326 -6455
rect 12268 -6525 12280 -6489
rect 12314 -6525 12326 -6489
rect 12268 -6537 12326 -6525
rect 12526 -6349 12584 -6337
rect 12526 -6385 12538 -6349
rect 12572 -6385 12584 -6349
rect 12526 -6419 12584 -6385
rect 12526 -6455 12538 -6419
rect 12572 -6455 12584 -6419
rect 12526 -6489 12584 -6455
rect 12526 -6525 12538 -6489
rect 12572 -6525 12584 -6489
rect 12526 -6537 12584 -6525
rect 5129 -6768 5187 -6756
rect 5129 -6804 5141 -6768
rect 5175 -6804 5187 -6768
rect 5129 -6838 5187 -6804
rect 5129 -6874 5141 -6838
rect 5175 -6874 5187 -6838
rect 5129 -6908 5187 -6874
rect 5129 -6944 5141 -6908
rect 5175 -6944 5187 -6908
rect 5129 -6956 5187 -6944
rect 5387 -6768 5445 -6756
rect 5387 -6804 5399 -6768
rect 5433 -6804 5445 -6768
rect 5387 -6838 5445 -6804
rect 5387 -6874 5399 -6838
rect 5433 -6874 5445 -6838
rect 5387 -6908 5445 -6874
rect 5387 -6944 5399 -6908
rect 5433 -6944 5445 -6908
rect 5387 -6956 5445 -6944
rect 5645 -6768 5703 -6756
rect 5645 -6804 5657 -6768
rect 5691 -6804 5703 -6768
rect 5645 -6838 5703 -6804
rect 5645 -6874 5657 -6838
rect 5691 -6874 5703 -6838
rect 5645 -6909 5703 -6874
rect 5645 -6945 5657 -6909
rect 5691 -6945 5703 -6909
rect 5645 -6956 5703 -6945
rect 5903 -6768 5961 -6756
rect 5903 -6804 5915 -6768
rect 5949 -6804 5961 -6768
rect 5903 -6838 5961 -6804
rect 5903 -6874 5915 -6838
rect 5949 -6874 5961 -6838
rect 5903 -6908 5961 -6874
rect 5903 -6944 5915 -6908
rect 5949 -6944 5961 -6908
rect 5903 -6956 5961 -6944
rect 6161 -6768 6219 -6756
rect 6161 -6804 6173 -6768
rect 6207 -6804 6219 -6768
rect 6161 -6838 6219 -6804
rect 6161 -6874 6173 -6838
rect 6207 -6874 6219 -6838
rect 6161 -6908 6219 -6874
rect 6161 -6944 6173 -6908
rect 6207 -6944 6219 -6908
rect 6161 -6956 6219 -6944
rect 6419 -6768 6477 -6756
rect 6419 -6804 6431 -6768
rect 6465 -6804 6477 -6768
rect 6419 -6838 6477 -6804
rect 6419 -6874 6431 -6838
rect 6465 -6874 6477 -6838
rect 6419 -6908 6477 -6874
rect 6419 -6944 6431 -6908
rect 6465 -6944 6477 -6908
rect 6419 -6956 6477 -6944
rect 6677 -6768 6735 -6756
rect 6677 -6804 6689 -6768
rect 6723 -6804 6735 -6768
rect 6677 -6838 6735 -6804
rect 6677 -6874 6689 -6838
rect 6723 -6874 6735 -6838
rect 6677 -6908 6735 -6874
rect 6677 -6944 6689 -6908
rect 6723 -6944 6735 -6908
rect 6677 -6956 6735 -6944
rect 6935 -6768 6993 -6756
rect 6935 -6804 6947 -6768
rect 6981 -6804 6993 -6768
rect 6935 -6838 6993 -6804
rect 6935 -6874 6947 -6838
rect 6981 -6874 6993 -6838
rect 6935 -6908 6993 -6874
rect 6935 -6944 6947 -6908
rect 6981 -6944 6993 -6908
rect 6935 -6956 6993 -6944
rect 7193 -6768 7251 -6756
rect 7193 -6804 7205 -6768
rect 7239 -6804 7251 -6768
rect 7193 -6838 7251 -6804
rect 7193 -6874 7205 -6838
rect 7239 -6874 7251 -6838
rect 7193 -6908 7251 -6874
rect 7193 -6944 7205 -6908
rect 7239 -6944 7251 -6908
rect 7193 -6956 7251 -6944
rect 7799 -6768 7857 -6756
rect 7799 -6804 7811 -6768
rect 7845 -6804 7857 -6768
rect 7799 -6838 7857 -6804
rect 7799 -6874 7811 -6838
rect 7845 -6874 7857 -6838
rect 7799 -6908 7857 -6874
rect 7799 -6944 7811 -6908
rect 7845 -6944 7857 -6908
rect 7799 -6956 7857 -6944
rect 8057 -6768 8115 -6756
rect 8057 -6804 8069 -6768
rect 8103 -6804 8115 -6768
rect 8057 -6838 8115 -6804
rect 8057 -6874 8069 -6838
rect 8103 -6874 8115 -6838
rect 8057 -6908 8115 -6874
rect 8057 -6944 8069 -6908
rect 8103 -6944 8115 -6908
rect 8057 -6956 8115 -6944
rect 8315 -6768 8373 -6756
rect 8315 -6804 8327 -6768
rect 8361 -6804 8373 -6768
rect 8315 -6838 8373 -6804
rect 8315 -6874 8327 -6838
rect 8361 -6874 8373 -6838
rect 8315 -6909 8373 -6874
rect 8315 -6945 8327 -6909
rect 8361 -6945 8373 -6909
rect 8315 -6956 8373 -6945
rect 8573 -6768 8631 -6756
rect 8573 -6804 8585 -6768
rect 8619 -6804 8631 -6768
rect 8573 -6838 8631 -6804
rect 8573 -6874 8585 -6838
rect 8619 -6874 8631 -6838
rect 8573 -6908 8631 -6874
rect 8573 -6944 8585 -6908
rect 8619 -6944 8631 -6908
rect 8573 -6956 8631 -6944
rect 8831 -6768 8889 -6756
rect 8831 -6804 8843 -6768
rect 8877 -6804 8889 -6768
rect 8831 -6838 8889 -6804
rect 8831 -6874 8843 -6838
rect 8877 -6874 8889 -6838
rect 8831 -6908 8889 -6874
rect 8831 -6944 8843 -6908
rect 8877 -6944 8889 -6908
rect 8831 -6956 8889 -6944
rect 9089 -6768 9147 -6756
rect 9089 -6804 9101 -6768
rect 9135 -6804 9147 -6768
rect 9089 -6838 9147 -6804
rect 9089 -6874 9101 -6838
rect 9135 -6874 9147 -6838
rect 9089 -6908 9147 -6874
rect 9089 -6944 9101 -6908
rect 9135 -6944 9147 -6908
rect 9089 -6956 9147 -6944
rect 9347 -6768 9405 -6756
rect 9347 -6804 9359 -6768
rect 9393 -6804 9405 -6768
rect 9347 -6838 9405 -6804
rect 9347 -6874 9359 -6838
rect 9393 -6874 9405 -6838
rect 9347 -6908 9405 -6874
rect 9347 -6944 9359 -6908
rect 9393 -6944 9405 -6908
rect 9347 -6956 9405 -6944
rect 9605 -6768 9663 -6756
rect 9605 -6804 9617 -6768
rect 9651 -6804 9663 -6768
rect 9605 -6838 9663 -6804
rect 9605 -6874 9617 -6838
rect 9651 -6874 9663 -6838
rect 9605 -6908 9663 -6874
rect 9605 -6944 9617 -6908
rect 9651 -6944 9663 -6908
rect 9605 -6956 9663 -6944
rect 9863 -6768 9921 -6756
rect 9863 -6804 9875 -6768
rect 9909 -6804 9921 -6768
rect 9863 -6838 9921 -6804
rect 9863 -6874 9875 -6838
rect 9909 -6874 9921 -6838
rect 9863 -6908 9921 -6874
rect 9863 -6944 9875 -6908
rect 9909 -6944 9921 -6908
rect 9863 -6956 9921 -6944
rect 10462 -6767 10520 -6755
rect 10462 -6803 10474 -6767
rect 10508 -6803 10520 -6767
rect 10462 -6837 10520 -6803
rect 10462 -6873 10474 -6837
rect 10508 -6873 10520 -6837
rect 10462 -6907 10520 -6873
rect 10462 -6943 10474 -6907
rect 10508 -6943 10520 -6907
rect 10462 -6955 10520 -6943
rect 10720 -6767 10778 -6755
rect 10720 -6803 10732 -6767
rect 10766 -6803 10778 -6767
rect 10720 -6837 10778 -6803
rect 10720 -6873 10732 -6837
rect 10766 -6873 10778 -6837
rect 10720 -6907 10778 -6873
rect 10720 -6943 10732 -6907
rect 10766 -6943 10778 -6907
rect 10720 -6955 10778 -6943
rect 10978 -6767 11036 -6755
rect 10978 -6803 10990 -6767
rect 11024 -6803 11036 -6767
rect 10978 -6837 11036 -6803
rect 10978 -6873 10990 -6837
rect 11024 -6873 11036 -6837
rect 10978 -6908 11036 -6873
rect 10978 -6944 10990 -6908
rect 11024 -6944 11036 -6908
rect 10978 -6955 11036 -6944
rect 11236 -6767 11294 -6755
rect 11236 -6803 11248 -6767
rect 11282 -6803 11294 -6767
rect 11236 -6837 11294 -6803
rect 11236 -6873 11248 -6837
rect 11282 -6873 11294 -6837
rect 11236 -6907 11294 -6873
rect 11236 -6943 11248 -6907
rect 11282 -6943 11294 -6907
rect 11236 -6955 11294 -6943
rect 11494 -6767 11552 -6755
rect 11494 -6803 11506 -6767
rect 11540 -6803 11552 -6767
rect 11494 -6837 11552 -6803
rect 11494 -6873 11506 -6837
rect 11540 -6873 11552 -6837
rect 11494 -6907 11552 -6873
rect 11494 -6943 11506 -6907
rect 11540 -6943 11552 -6907
rect 11494 -6955 11552 -6943
rect 11752 -6767 11810 -6755
rect 11752 -6803 11764 -6767
rect 11798 -6803 11810 -6767
rect 11752 -6837 11810 -6803
rect 11752 -6873 11764 -6837
rect 11798 -6873 11810 -6837
rect 11752 -6907 11810 -6873
rect 11752 -6943 11764 -6907
rect 11798 -6943 11810 -6907
rect 11752 -6955 11810 -6943
rect 12010 -6767 12068 -6755
rect 12010 -6803 12022 -6767
rect 12056 -6803 12068 -6767
rect 12010 -6837 12068 -6803
rect 12010 -6873 12022 -6837
rect 12056 -6873 12068 -6837
rect 12010 -6907 12068 -6873
rect 12010 -6943 12022 -6907
rect 12056 -6943 12068 -6907
rect 12010 -6955 12068 -6943
rect 12268 -6767 12326 -6755
rect 12268 -6803 12280 -6767
rect 12314 -6803 12326 -6767
rect 12268 -6837 12326 -6803
rect 12268 -6873 12280 -6837
rect 12314 -6873 12326 -6837
rect 12268 -6907 12326 -6873
rect 12268 -6943 12280 -6907
rect 12314 -6943 12326 -6907
rect 12268 -6955 12326 -6943
rect 12526 -6767 12584 -6755
rect 12526 -6803 12538 -6767
rect 12572 -6803 12584 -6767
rect 12526 -6837 12584 -6803
rect 12526 -6873 12538 -6837
rect 12572 -6873 12584 -6837
rect 12526 -6907 12584 -6873
rect 12526 -6943 12538 -6907
rect 12572 -6943 12584 -6907
rect 12526 -6955 12584 -6943
rect 5129 -7186 5187 -7174
rect 5129 -7222 5141 -7186
rect 5175 -7222 5187 -7186
rect 5129 -7256 5187 -7222
rect 5129 -7292 5141 -7256
rect 5175 -7292 5187 -7256
rect 5129 -7326 5187 -7292
rect 5129 -7362 5141 -7326
rect 5175 -7362 5187 -7326
rect 5129 -7374 5187 -7362
rect 5387 -7186 5445 -7174
rect 5387 -7222 5399 -7186
rect 5433 -7222 5445 -7186
rect 5387 -7256 5445 -7222
rect 5387 -7292 5399 -7256
rect 5433 -7292 5445 -7256
rect 5387 -7326 5445 -7292
rect 5387 -7362 5399 -7326
rect 5433 -7362 5445 -7326
rect 5387 -7374 5445 -7362
rect 5645 -7186 5703 -7174
rect 5645 -7222 5657 -7186
rect 5691 -7222 5703 -7186
rect 5645 -7256 5703 -7222
rect 5645 -7292 5657 -7256
rect 5691 -7292 5703 -7256
rect 5645 -7327 5703 -7292
rect 5645 -7363 5657 -7327
rect 5691 -7363 5703 -7327
rect 5645 -7374 5703 -7363
rect 5903 -7186 5961 -7174
rect 5903 -7222 5915 -7186
rect 5949 -7222 5961 -7186
rect 5903 -7256 5961 -7222
rect 5903 -7292 5915 -7256
rect 5949 -7292 5961 -7256
rect 5903 -7326 5961 -7292
rect 5903 -7362 5915 -7326
rect 5949 -7362 5961 -7326
rect 5903 -7374 5961 -7362
rect 6161 -7186 6219 -7174
rect 6161 -7222 6173 -7186
rect 6207 -7222 6219 -7186
rect 6161 -7256 6219 -7222
rect 6161 -7292 6173 -7256
rect 6207 -7292 6219 -7256
rect 6161 -7326 6219 -7292
rect 6161 -7362 6173 -7326
rect 6207 -7362 6219 -7326
rect 6161 -7374 6219 -7362
rect 6419 -7186 6477 -7174
rect 6419 -7222 6431 -7186
rect 6465 -7222 6477 -7186
rect 6419 -7256 6477 -7222
rect 6419 -7292 6431 -7256
rect 6465 -7292 6477 -7256
rect 6419 -7326 6477 -7292
rect 6419 -7362 6431 -7326
rect 6465 -7362 6477 -7326
rect 6419 -7374 6477 -7362
rect 6677 -7186 6735 -7174
rect 6677 -7222 6689 -7186
rect 6723 -7222 6735 -7186
rect 6677 -7256 6735 -7222
rect 6677 -7292 6689 -7256
rect 6723 -7292 6735 -7256
rect 6677 -7326 6735 -7292
rect 6677 -7362 6689 -7326
rect 6723 -7362 6735 -7326
rect 6677 -7374 6735 -7362
rect 6935 -7186 6993 -7174
rect 6935 -7222 6947 -7186
rect 6981 -7222 6993 -7186
rect 6935 -7256 6993 -7222
rect 6935 -7292 6947 -7256
rect 6981 -7292 6993 -7256
rect 6935 -7326 6993 -7292
rect 6935 -7362 6947 -7326
rect 6981 -7362 6993 -7326
rect 6935 -7374 6993 -7362
rect 7193 -7186 7251 -7174
rect 7193 -7222 7205 -7186
rect 7239 -7222 7251 -7186
rect 7193 -7256 7251 -7222
rect 7193 -7292 7205 -7256
rect 7239 -7292 7251 -7256
rect 7193 -7326 7251 -7292
rect 7193 -7362 7205 -7326
rect 7239 -7362 7251 -7326
rect 7193 -7374 7251 -7362
rect 7799 -7186 7857 -7174
rect 7799 -7222 7811 -7186
rect 7845 -7222 7857 -7186
rect 7799 -7256 7857 -7222
rect 7799 -7292 7811 -7256
rect 7845 -7292 7857 -7256
rect 7799 -7326 7857 -7292
rect 7799 -7362 7811 -7326
rect 7845 -7362 7857 -7326
rect 7799 -7374 7857 -7362
rect 8057 -7186 8115 -7174
rect 8057 -7222 8069 -7186
rect 8103 -7222 8115 -7186
rect 8057 -7256 8115 -7222
rect 8057 -7292 8069 -7256
rect 8103 -7292 8115 -7256
rect 8057 -7326 8115 -7292
rect 8057 -7362 8069 -7326
rect 8103 -7362 8115 -7326
rect 8057 -7374 8115 -7362
rect 8315 -7186 8373 -7174
rect 8315 -7222 8327 -7186
rect 8361 -7222 8373 -7186
rect 8315 -7256 8373 -7222
rect 8315 -7292 8327 -7256
rect 8361 -7292 8373 -7256
rect 8315 -7327 8373 -7292
rect 8315 -7363 8327 -7327
rect 8361 -7363 8373 -7327
rect 8315 -7374 8373 -7363
rect 8573 -7186 8631 -7174
rect 8573 -7222 8585 -7186
rect 8619 -7222 8631 -7186
rect 8573 -7256 8631 -7222
rect 8573 -7292 8585 -7256
rect 8619 -7292 8631 -7256
rect 8573 -7326 8631 -7292
rect 8573 -7362 8585 -7326
rect 8619 -7362 8631 -7326
rect 8573 -7374 8631 -7362
rect 8831 -7186 8889 -7174
rect 8831 -7222 8843 -7186
rect 8877 -7222 8889 -7186
rect 8831 -7256 8889 -7222
rect 8831 -7292 8843 -7256
rect 8877 -7292 8889 -7256
rect 8831 -7326 8889 -7292
rect 8831 -7362 8843 -7326
rect 8877 -7362 8889 -7326
rect 8831 -7374 8889 -7362
rect 9089 -7186 9147 -7174
rect 9089 -7222 9101 -7186
rect 9135 -7222 9147 -7186
rect 9089 -7256 9147 -7222
rect 9089 -7292 9101 -7256
rect 9135 -7292 9147 -7256
rect 9089 -7326 9147 -7292
rect 9089 -7362 9101 -7326
rect 9135 -7362 9147 -7326
rect 9089 -7374 9147 -7362
rect 9347 -7186 9405 -7174
rect 9347 -7222 9359 -7186
rect 9393 -7222 9405 -7186
rect 9347 -7256 9405 -7222
rect 9347 -7292 9359 -7256
rect 9393 -7292 9405 -7256
rect 9347 -7326 9405 -7292
rect 9347 -7362 9359 -7326
rect 9393 -7362 9405 -7326
rect 9347 -7374 9405 -7362
rect 9605 -7186 9663 -7174
rect 9605 -7222 9617 -7186
rect 9651 -7222 9663 -7186
rect 9605 -7256 9663 -7222
rect 9605 -7292 9617 -7256
rect 9651 -7292 9663 -7256
rect 9605 -7326 9663 -7292
rect 9605 -7362 9617 -7326
rect 9651 -7362 9663 -7326
rect 9605 -7374 9663 -7362
rect 9863 -7186 9921 -7174
rect 9863 -7222 9875 -7186
rect 9909 -7222 9921 -7186
rect 9863 -7256 9921 -7222
rect 9863 -7292 9875 -7256
rect 9909 -7292 9921 -7256
rect 9863 -7326 9921 -7292
rect 9863 -7362 9875 -7326
rect 9909 -7362 9921 -7326
rect 9863 -7374 9921 -7362
rect 10462 -7185 10520 -7173
rect 10462 -7221 10474 -7185
rect 10508 -7221 10520 -7185
rect 10462 -7255 10520 -7221
rect 10462 -7291 10474 -7255
rect 10508 -7291 10520 -7255
rect 10462 -7325 10520 -7291
rect 10462 -7361 10474 -7325
rect 10508 -7361 10520 -7325
rect 10462 -7373 10520 -7361
rect 10720 -7185 10778 -7173
rect 10720 -7221 10732 -7185
rect 10766 -7221 10778 -7185
rect 10720 -7255 10778 -7221
rect 10720 -7291 10732 -7255
rect 10766 -7291 10778 -7255
rect 10720 -7325 10778 -7291
rect 10720 -7361 10732 -7325
rect 10766 -7361 10778 -7325
rect 10720 -7373 10778 -7361
rect 10978 -7185 11036 -7173
rect 10978 -7221 10990 -7185
rect 11024 -7221 11036 -7185
rect 10978 -7255 11036 -7221
rect 10978 -7291 10990 -7255
rect 11024 -7291 11036 -7255
rect 10978 -7326 11036 -7291
rect 10978 -7362 10990 -7326
rect 11024 -7362 11036 -7326
rect 10978 -7373 11036 -7362
rect 11236 -7185 11294 -7173
rect 11236 -7221 11248 -7185
rect 11282 -7221 11294 -7185
rect 11236 -7255 11294 -7221
rect 11236 -7291 11248 -7255
rect 11282 -7291 11294 -7255
rect 11236 -7325 11294 -7291
rect 11236 -7361 11248 -7325
rect 11282 -7361 11294 -7325
rect 11236 -7373 11294 -7361
rect 11494 -7185 11552 -7173
rect 11494 -7221 11506 -7185
rect 11540 -7221 11552 -7185
rect 11494 -7255 11552 -7221
rect 11494 -7291 11506 -7255
rect 11540 -7291 11552 -7255
rect 11494 -7325 11552 -7291
rect 11494 -7361 11506 -7325
rect 11540 -7361 11552 -7325
rect 11494 -7373 11552 -7361
rect 11752 -7185 11810 -7173
rect 11752 -7221 11764 -7185
rect 11798 -7221 11810 -7185
rect 11752 -7255 11810 -7221
rect 11752 -7291 11764 -7255
rect 11798 -7291 11810 -7255
rect 11752 -7325 11810 -7291
rect 11752 -7361 11764 -7325
rect 11798 -7361 11810 -7325
rect 11752 -7373 11810 -7361
rect 12010 -7185 12068 -7173
rect 12010 -7221 12022 -7185
rect 12056 -7221 12068 -7185
rect 12010 -7255 12068 -7221
rect 12010 -7291 12022 -7255
rect 12056 -7291 12068 -7255
rect 12010 -7325 12068 -7291
rect 12010 -7361 12022 -7325
rect 12056 -7361 12068 -7325
rect 12010 -7373 12068 -7361
rect 12268 -7185 12326 -7173
rect 12268 -7221 12280 -7185
rect 12314 -7221 12326 -7185
rect 12268 -7255 12326 -7221
rect 12268 -7291 12280 -7255
rect 12314 -7291 12326 -7255
rect 12268 -7325 12326 -7291
rect 12268 -7361 12280 -7325
rect 12314 -7361 12326 -7325
rect 12268 -7373 12326 -7361
rect 12526 -7185 12584 -7173
rect 12526 -7221 12538 -7185
rect 12572 -7221 12584 -7185
rect 12526 -7255 12584 -7221
rect 12526 -7291 12538 -7255
rect 12572 -7291 12584 -7255
rect 12526 -7325 12584 -7291
rect 12526 -7361 12538 -7325
rect 12572 -7361 12584 -7325
rect 12526 -7373 12584 -7361
rect 5129 -7604 5187 -7592
rect 5129 -7640 5141 -7604
rect 5175 -7640 5187 -7604
rect 5129 -7674 5187 -7640
rect 5129 -7710 5141 -7674
rect 5175 -7710 5187 -7674
rect 5129 -7744 5187 -7710
rect 5129 -7780 5141 -7744
rect 5175 -7780 5187 -7744
rect 5129 -7792 5187 -7780
rect 5387 -7604 5445 -7592
rect 5387 -7640 5399 -7604
rect 5433 -7640 5445 -7604
rect 5387 -7674 5445 -7640
rect 5387 -7710 5399 -7674
rect 5433 -7710 5445 -7674
rect 5387 -7744 5445 -7710
rect 5387 -7780 5399 -7744
rect 5433 -7780 5445 -7744
rect 5387 -7792 5445 -7780
rect 5645 -7604 5703 -7592
rect 5645 -7640 5657 -7604
rect 5691 -7640 5703 -7604
rect 5645 -7674 5703 -7640
rect 5645 -7710 5657 -7674
rect 5691 -7710 5703 -7674
rect 5645 -7745 5703 -7710
rect 5645 -7781 5657 -7745
rect 5691 -7781 5703 -7745
rect 5645 -7792 5703 -7781
rect 5903 -7604 5961 -7592
rect 5903 -7640 5915 -7604
rect 5949 -7640 5961 -7604
rect 5903 -7674 5961 -7640
rect 5903 -7710 5915 -7674
rect 5949 -7710 5961 -7674
rect 5903 -7744 5961 -7710
rect 5903 -7780 5915 -7744
rect 5949 -7780 5961 -7744
rect 5903 -7792 5961 -7780
rect 6161 -7604 6219 -7592
rect 6161 -7640 6173 -7604
rect 6207 -7640 6219 -7604
rect 6161 -7674 6219 -7640
rect 6161 -7710 6173 -7674
rect 6207 -7710 6219 -7674
rect 6161 -7744 6219 -7710
rect 6161 -7780 6173 -7744
rect 6207 -7780 6219 -7744
rect 6161 -7792 6219 -7780
rect 6419 -7604 6477 -7592
rect 6419 -7640 6431 -7604
rect 6465 -7640 6477 -7604
rect 6419 -7674 6477 -7640
rect 6419 -7710 6431 -7674
rect 6465 -7710 6477 -7674
rect 6419 -7744 6477 -7710
rect 6419 -7780 6431 -7744
rect 6465 -7780 6477 -7744
rect 6419 -7792 6477 -7780
rect 6677 -7604 6735 -7592
rect 6677 -7640 6689 -7604
rect 6723 -7640 6735 -7604
rect 6677 -7674 6735 -7640
rect 6677 -7710 6689 -7674
rect 6723 -7710 6735 -7674
rect 6677 -7744 6735 -7710
rect 6677 -7780 6689 -7744
rect 6723 -7780 6735 -7744
rect 6677 -7792 6735 -7780
rect 6935 -7604 6993 -7592
rect 6935 -7640 6947 -7604
rect 6981 -7640 6993 -7604
rect 6935 -7674 6993 -7640
rect 6935 -7710 6947 -7674
rect 6981 -7710 6993 -7674
rect 6935 -7744 6993 -7710
rect 6935 -7780 6947 -7744
rect 6981 -7780 6993 -7744
rect 6935 -7792 6993 -7780
rect 7193 -7604 7251 -7592
rect 7193 -7640 7205 -7604
rect 7239 -7640 7251 -7604
rect 7193 -7674 7251 -7640
rect 7193 -7710 7205 -7674
rect 7239 -7710 7251 -7674
rect 7193 -7744 7251 -7710
rect 7193 -7780 7205 -7744
rect 7239 -7780 7251 -7744
rect 7193 -7792 7251 -7780
rect 7799 -7604 7857 -7592
rect 7799 -7640 7811 -7604
rect 7845 -7640 7857 -7604
rect 7799 -7674 7857 -7640
rect 7799 -7710 7811 -7674
rect 7845 -7710 7857 -7674
rect 7799 -7744 7857 -7710
rect 7799 -7780 7811 -7744
rect 7845 -7780 7857 -7744
rect 7799 -7792 7857 -7780
rect 8057 -7604 8115 -7592
rect 8057 -7640 8069 -7604
rect 8103 -7640 8115 -7604
rect 8057 -7674 8115 -7640
rect 8057 -7710 8069 -7674
rect 8103 -7710 8115 -7674
rect 8057 -7744 8115 -7710
rect 8057 -7780 8069 -7744
rect 8103 -7780 8115 -7744
rect 8057 -7792 8115 -7780
rect 8315 -7604 8373 -7592
rect 8315 -7640 8327 -7604
rect 8361 -7640 8373 -7604
rect 8315 -7674 8373 -7640
rect 8315 -7710 8327 -7674
rect 8361 -7710 8373 -7674
rect 8315 -7745 8373 -7710
rect 8315 -7781 8327 -7745
rect 8361 -7781 8373 -7745
rect 8315 -7792 8373 -7781
rect 8573 -7604 8631 -7592
rect 8573 -7640 8585 -7604
rect 8619 -7640 8631 -7604
rect 8573 -7674 8631 -7640
rect 8573 -7710 8585 -7674
rect 8619 -7710 8631 -7674
rect 8573 -7744 8631 -7710
rect 8573 -7780 8585 -7744
rect 8619 -7780 8631 -7744
rect 8573 -7792 8631 -7780
rect 8831 -7604 8889 -7592
rect 8831 -7640 8843 -7604
rect 8877 -7640 8889 -7604
rect 8831 -7674 8889 -7640
rect 8831 -7710 8843 -7674
rect 8877 -7710 8889 -7674
rect 8831 -7744 8889 -7710
rect 8831 -7780 8843 -7744
rect 8877 -7780 8889 -7744
rect 8831 -7792 8889 -7780
rect 9089 -7604 9147 -7592
rect 9089 -7640 9101 -7604
rect 9135 -7640 9147 -7604
rect 9089 -7674 9147 -7640
rect 9089 -7710 9101 -7674
rect 9135 -7710 9147 -7674
rect 9089 -7744 9147 -7710
rect 9089 -7780 9101 -7744
rect 9135 -7780 9147 -7744
rect 9089 -7792 9147 -7780
rect 9347 -7604 9405 -7592
rect 9347 -7640 9359 -7604
rect 9393 -7640 9405 -7604
rect 9347 -7674 9405 -7640
rect 9347 -7710 9359 -7674
rect 9393 -7710 9405 -7674
rect 9347 -7744 9405 -7710
rect 9347 -7780 9359 -7744
rect 9393 -7780 9405 -7744
rect 9347 -7792 9405 -7780
rect 9605 -7604 9663 -7592
rect 9605 -7640 9617 -7604
rect 9651 -7640 9663 -7604
rect 9605 -7674 9663 -7640
rect 9605 -7710 9617 -7674
rect 9651 -7710 9663 -7674
rect 9605 -7744 9663 -7710
rect 9605 -7780 9617 -7744
rect 9651 -7780 9663 -7744
rect 9605 -7792 9663 -7780
rect 9863 -7604 9921 -7592
rect 9863 -7640 9875 -7604
rect 9909 -7640 9921 -7604
rect 9863 -7674 9921 -7640
rect 9863 -7710 9875 -7674
rect 9909 -7710 9921 -7674
rect 9863 -7744 9921 -7710
rect 9863 -7780 9875 -7744
rect 9909 -7780 9921 -7744
rect 9863 -7792 9921 -7780
rect 10462 -7603 10520 -7591
rect 10462 -7639 10474 -7603
rect 10508 -7639 10520 -7603
rect 10462 -7673 10520 -7639
rect 10462 -7709 10474 -7673
rect 10508 -7709 10520 -7673
rect 10462 -7743 10520 -7709
rect 10462 -7779 10474 -7743
rect 10508 -7779 10520 -7743
rect 10462 -7791 10520 -7779
rect 10720 -7603 10778 -7591
rect 10720 -7639 10732 -7603
rect 10766 -7639 10778 -7603
rect 10720 -7673 10778 -7639
rect 10720 -7709 10732 -7673
rect 10766 -7709 10778 -7673
rect 10720 -7743 10778 -7709
rect 10720 -7779 10732 -7743
rect 10766 -7779 10778 -7743
rect 10720 -7791 10778 -7779
rect 10978 -7603 11036 -7591
rect 10978 -7639 10990 -7603
rect 11024 -7639 11036 -7603
rect 10978 -7673 11036 -7639
rect 10978 -7709 10990 -7673
rect 11024 -7709 11036 -7673
rect 10978 -7744 11036 -7709
rect 10978 -7780 10990 -7744
rect 11024 -7780 11036 -7744
rect 10978 -7791 11036 -7780
rect 11236 -7603 11294 -7591
rect 11236 -7639 11248 -7603
rect 11282 -7639 11294 -7603
rect 11236 -7673 11294 -7639
rect 11236 -7709 11248 -7673
rect 11282 -7709 11294 -7673
rect 11236 -7743 11294 -7709
rect 11236 -7779 11248 -7743
rect 11282 -7779 11294 -7743
rect 11236 -7791 11294 -7779
rect 11494 -7603 11552 -7591
rect 11494 -7639 11506 -7603
rect 11540 -7639 11552 -7603
rect 11494 -7673 11552 -7639
rect 11494 -7709 11506 -7673
rect 11540 -7709 11552 -7673
rect 11494 -7743 11552 -7709
rect 11494 -7779 11506 -7743
rect 11540 -7779 11552 -7743
rect 11494 -7791 11552 -7779
rect 11752 -7603 11810 -7591
rect 11752 -7639 11764 -7603
rect 11798 -7639 11810 -7603
rect 11752 -7673 11810 -7639
rect 11752 -7709 11764 -7673
rect 11798 -7709 11810 -7673
rect 11752 -7743 11810 -7709
rect 11752 -7779 11764 -7743
rect 11798 -7779 11810 -7743
rect 11752 -7791 11810 -7779
rect 12010 -7603 12068 -7591
rect 12010 -7639 12022 -7603
rect 12056 -7639 12068 -7603
rect 12010 -7673 12068 -7639
rect 12010 -7709 12022 -7673
rect 12056 -7709 12068 -7673
rect 12010 -7743 12068 -7709
rect 12010 -7779 12022 -7743
rect 12056 -7779 12068 -7743
rect 12010 -7791 12068 -7779
rect 12268 -7603 12326 -7591
rect 12268 -7639 12280 -7603
rect 12314 -7639 12326 -7603
rect 12268 -7673 12326 -7639
rect 12268 -7709 12280 -7673
rect 12314 -7709 12326 -7673
rect 12268 -7743 12326 -7709
rect 12268 -7779 12280 -7743
rect 12314 -7779 12326 -7743
rect 12268 -7791 12326 -7779
rect 12526 -7603 12584 -7591
rect 12526 -7639 12538 -7603
rect 12572 -7639 12584 -7603
rect 12526 -7673 12584 -7639
rect 12526 -7709 12538 -7673
rect 12572 -7709 12584 -7673
rect 12526 -7743 12584 -7709
rect 12526 -7779 12538 -7743
rect 12572 -7779 12584 -7743
rect 12526 -7791 12584 -7779
rect 5009 -8258 5067 -8244
rect 5009 -8292 5021 -8258
rect 5055 -8292 5067 -8258
rect 5009 -8326 5067 -8292
rect 5009 -8362 5021 -8326
rect 5055 -8362 5067 -8326
rect 5009 -8396 5067 -8362
rect 5009 -8430 5021 -8396
rect 5055 -8430 5067 -8396
rect 5009 -8444 5067 -8430
rect 5267 -8258 5325 -8244
rect 5267 -8292 5279 -8258
rect 5313 -8292 5325 -8258
rect 5267 -8326 5325 -8292
rect 5267 -8362 5279 -8326
rect 5313 -8362 5325 -8326
rect 5267 -8396 5325 -8362
rect 5267 -8430 5279 -8396
rect 5313 -8430 5325 -8396
rect 5267 -8444 5325 -8430
rect 5549 -8258 5607 -8244
rect 5549 -8292 5561 -8258
rect 5595 -8292 5607 -8258
rect 5549 -8326 5607 -8292
rect 5549 -8362 5561 -8326
rect 5595 -8362 5607 -8326
rect 5549 -8396 5607 -8362
rect 5549 -8430 5561 -8396
rect 5595 -8430 5607 -8396
rect 5549 -8444 5607 -8430
rect 5807 -8258 5865 -8244
rect 5807 -8292 5819 -8258
rect 5853 -8292 5865 -8258
rect 5807 -8326 5865 -8292
rect 5807 -8362 5819 -8326
rect 5853 -8362 5865 -8326
rect 5807 -8396 5865 -8362
rect 5807 -8430 5819 -8396
rect 5853 -8430 5865 -8396
rect 5807 -8444 5865 -8430
rect 6029 -8258 6087 -8244
rect 6029 -8292 6041 -8258
rect 6075 -8292 6087 -8258
rect 6029 -8326 6087 -8292
rect 6029 -8362 6041 -8326
rect 6075 -8362 6087 -8326
rect 6029 -8396 6087 -8362
rect 6029 -8430 6041 -8396
rect 6075 -8430 6087 -8396
rect 6029 -8444 6087 -8430
rect 6287 -8258 6345 -8244
rect 6287 -8292 6299 -8258
rect 6333 -8292 6345 -8258
rect 6287 -8326 6345 -8292
rect 6287 -8362 6299 -8326
rect 6333 -8362 6345 -8326
rect 6287 -8396 6345 -8362
rect 6287 -8430 6299 -8396
rect 6333 -8430 6345 -8396
rect 6287 -8444 6345 -8430
rect 6532 -8256 6590 -8242
rect 6532 -8290 6544 -8256
rect 6578 -8290 6590 -8256
rect 6532 -8324 6590 -8290
rect 6532 -8360 6544 -8324
rect 6578 -8360 6590 -8324
rect 6532 -8394 6590 -8360
rect 6532 -8428 6544 -8394
rect 6578 -8428 6590 -8394
rect 6532 -8442 6590 -8428
rect 6790 -8256 6848 -8242
rect 6790 -8290 6802 -8256
rect 6836 -8290 6848 -8256
rect 6790 -8324 6848 -8290
rect 6790 -8360 6802 -8324
rect 6836 -8360 6848 -8324
rect 6790 -8394 6848 -8360
rect 6790 -8428 6802 -8394
rect 6836 -8428 6848 -8394
rect 6790 -8442 6848 -8428
rect 7042 -8246 7100 -8232
rect 7042 -8280 7054 -8246
rect 7088 -8280 7100 -8246
rect 7042 -8314 7100 -8280
rect 7042 -8350 7054 -8314
rect 7088 -8350 7100 -8314
rect 7042 -8384 7100 -8350
rect 7042 -8418 7054 -8384
rect 7088 -8418 7100 -8384
rect 7042 -8432 7100 -8418
rect 7300 -8246 7358 -8232
rect 7300 -8280 7312 -8246
rect 7346 -8280 7358 -8246
rect 7300 -8314 7358 -8280
rect 7300 -8350 7312 -8314
rect 7346 -8350 7358 -8314
rect 7300 -8384 7358 -8350
rect 7300 -8418 7312 -8384
rect 7346 -8418 7358 -8384
rect 7300 -8432 7358 -8418
rect 7679 -8258 7737 -8244
rect 7679 -8292 7691 -8258
rect 7725 -8292 7737 -8258
rect 7679 -8326 7737 -8292
rect 7679 -8362 7691 -8326
rect 7725 -8362 7737 -8326
rect 7679 -8396 7737 -8362
rect 7679 -8430 7691 -8396
rect 7725 -8430 7737 -8396
rect 7679 -8444 7737 -8430
rect 7937 -8258 7995 -8244
rect 7937 -8292 7949 -8258
rect 7983 -8292 7995 -8258
rect 7937 -8326 7995 -8292
rect 7937 -8362 7949 -8326
rect 7983 -8362 7995 -8326
rect 7937 -8396 7995 -8362
rect 7937 -8430 7949 -8396
rect 7983 -8430 7995 -8396
rect 7937 -8444 7995 -8430
rect 8219 -8258 8277 -8244
rect 8219 -8292 8231 -8258
rect 8265 -8292 8277 -8258
rect 8219 -8326 8277 -8292
rect 8219 -8362 8231 -8326
rect 8265 -8362 8277 -8326
rect 8219 -8396 8277 -8362
rect 8219 -8430 8231 -8396
rect 8265 -8430 8277 -8396
rect 8219 -8444 8277 -8430
rect 8477 -8258 8535 -8244
rect 8477 -8292 8489 -8258
rect 8523 -8292 8535 -8258
rect 8477 -8326 8535 -8292
rect 8477 -8362 8489 -8326
rect 8523 -8362 8535 -8326
rect 8477 -8396 8535 -8362
rect 8477 -8430 8489 -8396
rect 8523 -8430 8535 -8396
rect 8477 -8444 8535 -8430
rect 8699 -8258 8757 -8244
rect 8699 -8292 8711 -8258
rect 8745 -8292 8757 -8258
rect 8699 -8326 8757 -8292
rect 8699 -8362 8711 -8326
rect 8745 -8362 8757 -8326
rect 8699 -8396 8757 -8362
rect 8699 -8430 8711 -8396
rect 8745 -8430 8757 -8396
rect 8699 -8444 8757 -8430
rect 8957 -8258 9015 -8244
rect 8957 -8292 8969 -8258
rect 9003 -8292 9015 -8258
rect 8957 -8326 9015 -8292
rect 8957 -8362 8969 -8326
rect 9003 -8362 9015 -8326
rect 8957 -8396 9015 -8362
rect 8957 -8430 8969 -8396
rect 9003 -8430 9015 -8396
rect 8957 -8444 9015 -8430
rect 9202 -8256 9260 -8242
rect 9202 -8290 9214 -8256
rect 9248 -8290 9260 -8256
rect 9202 -8324 9260 -8290
rect 9202 -8360 9214 -8324
rect 9248 -8360 9260 -8324
rect 9202 -8394 9260 -8360
rect 9202 -8428 9214 -8394
rect 9248 -8428 9260 -8394
rect 9202 -8442 9260 -8428
rect 9460 -8256 9518 -8242
rect 9460 -8290 9472 -8256
rect 9506 -8290 9518 -8256
rect 9460 -8324 9518 -8290
rect 9460 -8360 9472 -8324
rect 9506 -8360 9518 -8324
rect 9460 -8394 9518 -8360
rect 9460 -8428 9472 -8394
rect 9506 -8428 9518 -8394
rect 9460 -8442 9518 -8428
rect 9712 -8246 9770 -8232
rect 9712 -8280 9724 -8246
rect 9758 -8280 9770 -8246
rect 9712 -8314 9770 -8280
rect 9712 -8350 9724 -8314
rect 9758 -8350 9770 -8314
rect 9712 -8384 9770 -8350
rect 9712 -8418 9724 -8384
rect 9758 -8418 9770 -8384
rect 9712 -8432 9770 -8418
rect 9970 -8246 10028 -8232
rect 9970 -8280 9982 -8246
rect 10016 -8280 10028 -8246
rect 9970 -8314 10028 -8280
rect 9970 -8350 9982 -8314
rect 10016 -8350 10028 -8314
rect 9970 -8384 10028 -8350
rect 9970 -8418 9982 -8384
rect 10016 -8418 10028 -8384
rect 9970 -8432 10028 -8418
rect 10342 -8257 10400 -8243
rect 10342 -8291 10354 -8257
rect 10388 -8291 10400 -8257
rect 10342 -8325 10400 -8291
rect 10342 -8361 10354 -8325
rect 10388 -8361 10400 -8325
rect 10342 -8395 10400 -8361
rect 10342 -8429 10354 -8395
rect 10388 -8429 10400 -8395
rect 10342 -8443 10400 -8429
rect 10600 -8257 10658 -8243
rect 10600 -8291 10612 -8257
rect 10646 -8291 10658 -8257
rect 10600 -8325 10658 -8291
rect 10600 -8361 10612 -8325
rect 10646 -8361 10658 -8325
rect 10600 -8395 10658 -8361
rect 10600 -8429 10612 -8395
rect 10646 -8429 10658 -8395
rect 10600 -8443 10658 -8429
rect 10882 -8257 10940 -8243
rect 10882 -8291 10894 -8257
rect 10928 -8291 10940 -8257
rect 10882 -8325 10940 -8291
rect 10882 -8361 10894 -8325
rect 10928 -8361 10940 -8325
rect 10882 -8395 10940 -8361
rect 10882 -8429 10894 -8395
rect 10928 -8429 10940 -8395
rect 10882 -8443 10940 -8429
rect 11140 -8257 11198 -8243
rect 11140 -8291 11152 -8257
rect 11186 -8291 11198 -8257
rect 11140 -8325 11198 -8291
rect 11140 -8361 11152 -8325
rect 11186 -8361 11198 -8325
rect 11140 -8395 11198 -8361
rect 11140 -8429 11152 -8395
rect 11186 -8429 11198 -8395
rect 11140 -8443 11198 -8429
rect 11362 -8257 11420 -8243
rect 11362 -8291 11374 -8257
rect 11408 -8291 11420 -8257
rect 11362 -8325 11420 -8291
rect 11362 -8361 11374 -8325
rect 11408 -8361 11420 -8325
rect 11362 -8395 11420 -8361
rect 11362 -8429 11374 -8395
rect 11408 -8429 11420 -8395
rect 11362 -8443 11420 -8429
rect 11620 -8257 11678 -8243
rect 11620 -8291 11632 -8257
rect 11666 -8291 11678 -8257
rect 11620 -8325 11678 -8291
rect 11620 -8361 11632 -8325
rect 11666 -8361 11678 -8325
rect 11620 -8395 11678 -8361
rect 11620 -8429 11632 -8395
rect 11666 -8429 11678 -8395
rect 11620 -8443 11678 -8429
rect 11865 -8255 11923 -8241
rect 11865 -8289 11877 -8255
rect 11911 -8289 11923 -8255
rect 11865 -8323 11923 -8289
rect 11865 -8359 11877 -8323
rect 11911 -8359 11923 -8323
rect 11865 -8393 11923 -8359
rect 11865 -8427 11877 -8393
rect 11911 -8427 11923 -8393
rect 11865 -8441 11923 -8427
rect 12123 -8255 12181 -8241
rect 12123 -8289 12135 -8255
rect 12169 -8289 12181 -8255
rect 12123 -8323 12181 -8289
rect 12123 -8359 12135 -8323
rect 12169 -8359 12181 -8323
rect 12123 -8393 12181 -8359
rect 12123 -8427 12135 -8393
rect 12169 -8427 12181 -8393
rect 12123 -8441 12181 -8427
rect 12375 -8245 12433 -8231
rect 12375 -8279 12387 -8245
rect 12421 -8279 12433 -8245
rect 12375 -8313 12433 -8279
rect 12375 -8349 12387 -8313
rect 12421 -8349 12433 -8313
rect 12375 -8383 12433 -8349
rect 12375 -8417 12387 -8383
rect 12421 -8417 12433 -8383
rect 12375 -8431 12433 -8417
rect 12633 -8245 12691 -8231
rect 12633 -8279 12645 -8245
rect 12679 -8279 12691 -8245
rect 12633 -8313 12691 -8279
rect 12633 -8349 12645 -8313
rect 12679 -8349 12691 -8313
rect 12633 -8383 12691 -8349
rect 12633 -8417 12645 -8383
rect 12679 -8417 12691 -8383
rect 12633 -8431 12691 -8417
rect 14006 8539 14064 8551
rect 14006 7163 14018 8539
rect 14052 7163 14064 8539
rect 14006 7151 14064 7163
rect 15664 8539 15722 8551
rect 15664 7163 15676 8539
rect 15710 7163 15722 8539
rect 15664 7151 15722 7163
rect 17322 8539 17380 8551
rect 17322 7163 17334 8539
rect 17368 7163 17380 8539
rect 17322 7151 17380 7163
rect 14006 7029 14064 7041
rect 14006 5653 14018 7029
rect 14052 5653 14064 7029
rect 14006 5641 14064 5653
rect 15664 7029 15722 7041
rect 15664 5653 15676 7029
rect 15710 5653 15722 7029
rect 15664 5641 15722 5653
rect 17322 7029 17380 7041
rect 17322 5653 17334 7029
rect 17368 5653 17380 7029
rect 17322 5641 17380 5653
rect 14006 5519 14064 5531
rect 14006 4143 14018 5519
rect 14052 4143 14064 5519
rect 14006 4131 14064 4143
rect 15664 5519 15722 5531
rect 15664 4143 15676 5519
rect 15710 4143 15722 5519
rect 15664 4131 15722 4143
rect 17322 5519 17380 5531
rect 17322 4143 17334 5519
rect 17368 4143 17380 5519
rect 17322 4131 17380 4143
rect 14006 4009 14064 4021
rect 14006 2633 14018 4009
rect 14052 2633 14064 4009
rect 14006 2621 14064 2633
rect 15664 4009 15722 4021
rect 15664 2633 15676 4009
rect 15710 2633 15722 4009
rect 15664 2621 15722 2633
rect 17322 4009 17380 4021
rect 17322 2633 17334 4009
rect 17368 2633 17380 4009
rect 17322 2621 17380 2633
rect 14006 2499 14064 2511
rect 14006 1123 14018 2499
rect 14052 1123 14064 2499
rect 14006 1111 14064 1123
rect 15664 2499 15722 2511
rect 15664 1123 15676 2499
rect 15710 1123 15722 2499
rect 15664 1111 15722 1123
rect 17322 2499 17380 2511
rect 17322 1123 17334 2499
rect 17368 1123 17380 2499
rect 17322 1111 17380 1123
rect 14006 989 14064 1001
rect 14006 -387 14018 989
rect 14052 -387 14064 989
rect 14006 -399 14064 -387
rect 15664 989 15722 1001
rect 15664 -387 15676 989
rect 15710 -387 15722 989
rect 15664 -399 15722 -387
rect 17322 989 17380 1001
rect 17322 -387 17334 989
rect 17368 -387 17380 989
rect 17322 -399 17380 -387
rect 14006 -521 14064 -509
rect 14006 -1897 14018 -521
rect 14052 -1897 14064 -521
rect 14006 -1909 14064 -1897
rect 15664 -521 15722 -509
rect 15664 -1897 15676 -521
rect 15710 -1897 15722 -521
rect 15664 -1909 15722 -1897
rect 17322 -521 17380 -509
rect 17322 -1897 17334 -521
rect 17368 -1897 17380 -521
rect 17322 -1909 17380 -1897
rect 14006 -2031 14064 -2019
rect 14006 -3407 14018 -2031
rect 14052 -3407 14064 -2031
rect 14006 -3419 14064 -3407
rect 15664 -2031 15722 -2019
rect 15664 -3407 15676 -2031
rect 15710 -3407 15722 -2031
rect 15664 -3419 15722 -3407
rect 17322 -2031 17380 -2019
rect 17322 -3407 17334 -2031
rect 17368 -3407 17380 -2031
rect 17322 -3419 17380 -3407
rect 14006 -3541 14064 -3529
rect 14006 -4917 14018 -3541
rect 14052 -4917 14064 -3541
rect 14006 -4929 14064 -4917
rect 15664 -3541 15722 -3529
rect 15664 -4917 15676 -3541
rect 15710 -4917 15722 -3541
rect 15664 -4929 15722 -4917
rect 17322 -3541 17380 -3529
rect 17322 -4917 17334 -3541
rect 17368 -4917 17380 -3541
rect 17322 -4929 17380 -4917
rect 14006 -5051 14064 -5039
rect 14006 -6427 14018 -5051
rect 14052 -6427 14064 -5051
rect 14006 -6439 14064 -6427
rect 15664 -5051 15722 -5039
rect 15664 -6427 15676 -5051
rect 15710 -6427 15722 -5051
rect 15664 -6439 15722 -6427
rect 17322 -5051 17380 -5039
rect 17322 -6427 17334 -5051
rect 17368 -6427 17380 -5051
rect 17322 -6439 17380 -6427
rect 14006 -6561 14064 -6549
rect 14006 -7937 14018 -6561
rect 14052 -7937 14064 -6561
rect 14006 -7949 14064 -7937
rect 15664 -6561 15722 -6549
rect 15664 -7937 15676 -6561
rect 15710 -7937 15722 -6561
rect 15664 -7949 15722 -7937
rect 17322 -6561 17380 -6549
rect 17322 -7937 17334 -6561
rect 17368 -7937 17380 -6561
rect 17322 -7949 17380 -7937
rect 14006 -8071 14064 -8059
rect 14006 -9447 14018 -8071
rect 14052 -9447 14064 -8071
rect 14006 -9459 14064 -9447
rect 15664 -8071 15722 -8059
rect 15664 -9447 15676 -8071
rect 15710 -9447 15722 -8071
rect 15664 -9459 15722 -9447
rect 17322 -8071 17380 -8059
rect 17322 -9447 17334 -8071
rect 17368 -9447 17380 -8071
rect 17322 -9459 17380 -9447
<< pdiff >>
rect 5403 8490 5461 8498
rect 5403 8454 5416 8490
rect 5450 8454 5461 8490
rect 5403 8416 5461 8454
rect 5403 8380 5415 8416
rect 5449 8380 5461 8416
rect 5403 8343 5461 8380
rect 5403 8307 5415 8343
rect 5449 8307 5461 8343
rect 5403 8298 5461 8307
rect 5661 8486 5719 8498
rect 5661 8450 5673 8486
rect 5707 8450 5719 8486
rect 5661 8416 5719 8450
rect 5661 8380 5673 8416
rect 5707 8380 5719 8416
rect 5661 8343 5719 8380
rect 5661 8307 5672 8343
rect 5706 8307 5719 8343
rect 5661 8298 5719 8307
rect 6063 8490 6121 8498
rect 6063 8454 6076 8490
rect 6110 8454 6121 8490
rect 6063 8416 6121 8454
rect 6063 8380 6075 8416
rect 6109 8380 6121 8416
rect 6063 8343 6121 8380
rect 6063 8307 6075 8343
rect 6109 8307 6121 8343
rect 6063 8298 6121 8307
rect 6321 8486 6379 8498
rect 6321 8450 6333 8486
rect 6367 8450 6379 8486
rect 6321 8416 6379 8450
rect 6321 8380 6333 8416
rect 6367 8380 6379 8416
rect 6321 8343 6379 8380
rect 6321 8307 6332 8343
rect 6366 8307 6379 8343
rect 6321 8298 6379 8307
rect 6533 8490 6591 8498
rect 6533 8454 6546 8490
rect 6580 8454 6591 8490
rect 6533 8416 6591 8454
rect 6533 8380 6545 8416
rect 6579 8380 6591 8416
rect 6533 8343 6591 8380
rect 6533 8307 6545 8343
rect 6579 8307 6591 8343
rect 6533 8298 6591 8307
rect 6791 8486 6849 8498
rect 6791 8450 6803 8486
rect 6837 8450 6849 8486
rect 6791 8416 6849 8450
rect 6791 8380 6803 8416
rect 6837 8380 6849 8416
rect 6791 8343 6849 8380
rect 6791 8307 6802 8343
rect 6836 8307 6849 8343
rect 6791 8298 6849 8307
rect 7136 8486 7194 8497
rect 7136 8450 7148 8486
rect 7182 8450 7194 8486
rect 7136 8415 7194 8450
rect 7136 8379 7148 8415
rect 7182 8379 7194 8415
rect 7136 8344 7194 8379
rect 7136 8308 7148 8344
rect 7182 8308 7194 8344
rect 7136 8297 7194 8308
rect 7394 8486 7452 8497
rect 7394 8450 7406 8486
rect 7440 8450 7452 8486
rect 7394 8415 7452 8450
rect 7394 8379 7406 8415
rect 7440 8379 7452 8415
rect 7394 8344 7452 8379
rect 7394 8308 7406 8344
rect 7440 8308 7452 8344
rect 7394 8297 7452 8308
rect 7652 8486 7710 8497
rect 7652 8450 7664 8486
rect 7698 8450 7710 8486
rect 7652 8415 7710 8450
rect 7652 8379 7664 8415
rect 7698 8379 7710 8415
rect 7652 8344 7710 8379
rect 7652 8308 7664 8344
rect 7698 8308 7710 8344
rect 7652 8297 7710 8308
rect 7910 8486 7968 8497
rect 7910 8450 7922 8486
rect 7956 8450 7968 8486
rect 7910 8415 7968 8450
rect 7910 8379 7922 8415
rect 7956 8379 7968 8415
rect 7910 8344 7968 8379
rect 7910 8308 7922 8344
rect 7956 8308 7968 8344
rect 7910 8297 7968 8308
rect 8168 8486 8226 8497
rect 8168 8450 8180 8486
rect 8214 8450 8226 8486
rect 8168 8415 8226 8450
rect 8168 8379 8180 8415
rect 8214 8379 8226 8415
rect 8168 8344 8226 8379
rect 8168 8308 8180 8344
rect 8214 8308 8226 8344
rect 8168 8297 8226 8308
rect 8426 8486 8484 8497
rect 8426 8450 8438 8486
rect 8472 8450 8484 8486
rect 8426 8415 8484 8450
rect 8426 8379 8438 8415
rect 8472 8379 8484 8415
rect 8426 8344 8484 8379
rect 8426 8308 8438 8344
rect 8472 8308 8484 8344
rect 8426 8297 8484 8308
rect 8951 8486 9009 8497
rect 8951 8450 8963 8486
rect 8997 8450 9009 8486
rect 8951 8415 9009 8450
rect 8951 8379 8963 8415
rect 8997 8379 9009 8415
rect 8951 8344 9009 8379
rect 8951 8308 8963 8344
rect 8997 8308 9009 8344
rect 8951 8297 9009 8308
rect 9209 8486 9267 8497
rect 9209 8450 9221 8486
rect 9255 8450 9267 8486
rect 9209 8415 9267 8450
rect 9209 8379 9221 8415
rect 9255 8379 9267 8415
rect 9209 8344 9267 8379
rect 9209 8308 9221 8344
rect 9255 8308 9267 8344
rect 9209 8297 9267 8308
rect 9467 8486 9525 8497
rect 9467 8450 9479 8486
rect 9513 8450 9525 8486
rect 9467 8415 9525 8450
rect 9467 8379 9479 8415
rect 9513 8379 9525 8415
rect 9467 8344 9525 8379
rect 9467 8308 9479 8344
rect 9513 8308 9525 8344
rect 9467 8297 9525 8308
rect 9725 8486 9783 8497
rect 9725 8450 9737 8486
rect 9771 8450 9783 8486
rect 9725 8415 9783 8450
rect 9725 8379 9737 8415
rect 9771 8379 9783 8415
rect 9725 8344 9783 8379
rect 9725 8308 9737 8344
rect 9771 8308 9783 8344
rect 9725 8297 9783 8308
rect 9983 8486 10041 8497
rect 9983 8450 9995 8486
rect 10029 8450 10041 8486
rect 9983 8415 10041 8450
rect 9983 8379 9995 8415
rect 10029 8379 10041 8415
rect 9983 8344 10041 8379
rect 9983 8308 9995 8344
rect 10029 8308 10041 8344
rect 9983 8297 10041 8308
rect 10241 8486 10299 8497
rect 10241 8450 10253 8486
rect 10287 8450 10299 8486
rect 10241 8415 10299 8450
rect 10241 8379 10253 8415
rect 10287 8379 10299 8415
rect 10241 8344 10299 8379
rect 10241 8308 10253 8344
rect 10287 8308 10299 8344
rect 10241 8297 10299 8308
rect 10757 8486 10815 8497
rect 10757 8450 10769 8486
rect 10803 8450 10815 8486
rect 10757 8415 10815 8450
rect 10757 8379 10769 8415
rect 10803 8379 10815 8415
rect 10757 8344 10815 8379
rect 10757 8308 10769 8344
rect 10803 8308 10815 8344
rect 10757 8297 10815 8308
rect 11015 8486 11073 8497
rect 11015 8450 11027 8486
rect 11061 8450 11073 8486
rect 11015 8415 11073 8450
rect 11015 8379 11027 8415
rect 11061 8379 11073 8415
rect 11015 8344 11073 8379
rect 11015 8308 11027 8344
rect 11061 8308 11073 8344
rect 11015 8297 11073 8308
rect 11273 8486 11331 8497
rect 11273 8450 11285 8486
rect 11319 8450 11331 8486
rect 11273 8415 11331 8450
rect 11273 8379 11285 8415
rect 11319 8379 11331 8415
rect 11273 8344 11331 8379
rect 11273 8308 11285 8344
rect 11319 8308 11331 8344
rect 11273 8297 11331 8308
rect 11531 8486 11589 8497
rect 11531 8450 11543 8486
rect 11577 8450 11589 8486
rect 11531 8415 11589 8450
rect 11531 8379 11543 8415
rect 11577 8379 11589 8415
rect 11531 8344 11589 8379
rect 11531 8308 11543 8344
rect 11577 8308 11589 8344
rect 11531 8297 11589 8308
rect 11789 8486 11847 8497
rect 11789 8450 11801 8486
rect 11835 8450 11847 8486
rect 11789 8415 11847 8450
rect 11789 8379 11801 8415
rect 11835 8379 11847 8415
rect 11789 8344 11847 8379
rect 11789 8308 11801 8344
rect 11835 8308 11847 8344
rect 11789 8297 11847 8308
rect 12047 8486 12105 8497
rect 12047 8450 12059 8486
rect 12093 8450 12105 8486
rect 12047 8415 12105 8450
rect 12047 8379 12059 8415
rect 12093 8379 12105 8415
rect 12047 8344 12105 8379
rect 12047 8308 12059 8344
rect 12093 8308 12105 8344
rect 12047 8297 12105 8308
rect 5338 7486 5412 7524
rect 5338 7450 5358 7486
rect 5396 7450 5412 7486
rect 5338 7414 5412 7450
rect 5528 7488 5602 7524
rect 5528 7452 5544 7488
rect 5582 7452 5602 7488
rect 5528 7414 5602 7452
rect 5707 7486 5765 7524
rect 5707 7452 5719 7486
rect 5753 7452 5765 7486
rect 5707 7414 5765 7452
rect 6565 7486 6623 7524
rect 6565 7452 6577 7486
rect 6611 7452 6623 7486
rect 6565 7414 6623 7452
rect 6724 7486 6798 7524
rect 6724 7450 6744 7486
rect 6782 7450 6798 7486
rect 6724 7414 6798 7450
rect 6914 7488 6988 7524
rect 6914 7452 6930 7488
rect 6968 7452 6988 7488
rect 6914 7414 6988 7452
rect 7094 7486 7168 7524
rect 7094 7450 7114 7486
rect 7152 7450 7168 7486
rect 7094 7414 7168 7450
rect 7284 7488 7358 7524
rect 7284 7452 7300 7488
rect 7338 7452 7358 7488
rect 7284 7414 7358 7452
rect 7516 7486 7590 7524
rect 7516 7450 7536 7486
rect 7574 7450 7590 7486
rect 7516 7414 7590 7450
rect 7706 7488 7780 7524
rect 7706 7452 7722 7488
rect 7760 7452 7780 7488
rect 7706 7414 7780 7452
rect 7938 7486 8012 7524
rect 7938 7450 7958 7486
rect 7996 7450 8012 7486
rect 7938 7414 8012 7450
rect 8128 7488 8202 7524
rect 8128 7452 8144 7488
rect 8182 7452 8202 7488
rect 8128 7414 8202 7452
rect 8377 7486 8435 7524
rect 8377 7452 8389 7486
rect 8423 7452 8435 7486
rect 8377 7414 8435 7452
rect 9235 7486 9293 7524
rect 9235 7452 9247 7486
rect 9281 7452 9293 7486
rect 9235 7414 9293 7452
rect 9438 7486 9512 7524
rect 9438 7450 9458 7486
rect 9496 7450 9512 7486
rect 9438 7414 9512 7450
rect 9628 7488 9702 7524
rect 9628 7452 9644 7488
rect 9682 7452 9702 7488
rect 9628 7414 9702 7452
rect 9808 7486 9882 7524
rect 9808 7450 9828 7486
rect 9866 7450 9882 7486
rect 9808 7414 9882 7450
rect 9998 7488 10072 7524
rect 9998 7452 10014 7488
rect 10052 7452 10072 7488
rect 9998 7414 10072 7452
rect 10230 7486 10304 7524
rect 10230 7450 10250 7486
rect 10288 7450 10304 7486
rect 10230 7414 10304 7450
rect 10420 7488 10494 7524
rect 10420 7452 10436 7488
rect 10474 7452 10494 7488
rect 10420 7414 10494 7452
rect 10652 7486 10726 7524
rect 10652 7450 10672 7486
rect 10710 7450 10726 7486
rect 10652 7414 10726 7450
rect 10842 7488 10916 7524
rect 10842 7452 10858 7488
rect 10896 7452 10916 7488
rect 10842 7414 10916 7452
rect 11040 7487 11098 7525
rect 11040 7453 11052 7487
rect 11086 7453 11098 7487
rect 11040 7415 11098 7453
rect 11898 7487 11956 7525
rect 11898 7453 11910 7487
rect 11944 7453 11956 7487
rect 11898 7415 11956 7453
rect 12092 7486 12166 7524
rect 12092 7450 12112 7486
rect 12150 7450 12166 7486
rect 12092 7414 12166 7450
rect 12282 7488 12356 7524
rect 12282 7452 12298 7488
rect 12336 7452 12356 7488
rect 12282 7414 12356 7452
rect 5338 1804 5412 1842
rect 5338 1768 5358 1804
rect 5396 1768 5412 1804
rect 5338 1732 5412 1768
rect 5528 1806 5602 1842
rect 5528 1770 5544 1806
rect 5582 1770 5602 1806
rect 5528 1732 5602 1770
rect 5699 1804 5757 1842
rect 5699 1770 5711 1804
rect 5745 1770 5757 1804
rect 5699 1732 5757 1770
rect 6557 1804 6615 1842
rect 6557 1770 6569 1804
rect 6603 1770 6615 1804
rect 6557 1732 6615 1770
rect 6724 1803 6798 1841
rect 6724 1767 6744 1803
rect 6782 1767 6798 1803
rect 6724 1731 6798 1767
rect 6914 1805 6988 1841
rect 6914 1769 6930 1805
rect 6968 1769 6988 1805
rect 6914 1731 6988 1769
rect 7094 1803 7168 1841
rect 7094 1767 7114 1803
rect 7152 1767 7168 1803
rect 7094 1731 7168 1767
rect 7284 1805 7358 1841
rect 7284 1769 7300 1805
rect 7338 1769 7358 1805
rect 7284 1731 7358 1769
rect 7516 1803 7590 1841
rect 7516 1767 7536 1803
rect 7574 1767 7590 1803
rect 7516 1731 7590 1767
rect 7706 1805 7780 1841
rect 7706 1769 7722 1805
rect 7760 1769 7780 1805
rect 7706 1731 7780 1769
rect 7938 1803 8012 1841
rect 7938 1767 7958 1803
rect 7996 1767 8012 1803
rect 7938 1731 8012 1767
rect 8128 1805 8202 1841
rect 8128 1769 8144 1805
rect 8182 1769 8202 1805
rect 8128 1731 8202 1769
rect 8375 1804 8434 1842
rect 8375 1770 8388 1804
rect 8422 1770 8434 1804
rect 8375 1735 8434 1770
rect 8376 1732 8434 1735
rect 9234 1804 9292 1842
rect 9234 1770 9246 1804
rect 9280 1770 9292 1804
rect 9234 1732 9292 1770
rect 9438 1807 9512 1845
rect 9438 1771 9458 1807
rect 9496 1771 9512 1807
rect 9438 1735 9512 1771
rect 9628 1809 9702 1845
rect 9628 1773 9644 1809
rect 9682 1773 9702 1809
rect 9628 1735 9702 1773
rect 9808 1807 9882 1845
rect 9808 1771 9828 1807
rect 9866 1771 9882 1807
rect 9808 1735 9882 1771
rect 9998 1809 10072 1845
rect 9998 1773 10014 1809
rect 10052 1773 10072 1809
rect 9998 1735 10072 1773
rect 10230 1807 10304 1845
rect 10230 1771 10250 1807
rect 10288 1771 10304 1807
rect 10230 1735 10304 1771
rect 10420 1809 10494 1845
rect 10420 1773 10436 1809
rect 10474 1773 10494 1809
rect 10420 1735 10494 1773
rect 10652 1807 10726 1845
rect 10652 1771 10672 1807
rect 10710 1771 10726 1807
rect 10652 1735 10726 1771
rect 10842 1809 10916 1845
rect 10842 1773 10858 1809
rect 10896 1773 10916 1809
rect 10842 1735 10916 1773
rect 11040 1805 11098 1843
rect 11040 1771 11052 1805
rect 11086 1771 11098 1805
rect 11040 1733 11098 1771
rect 11898 1805 11956 1843
rect 11898 1771 11910 1805
rect 11944 1771 11956 1805
rect 11898 1733 11956 1771
rect 12036 1804 12110 1842
rect 12036 1768 12056 1804
rect 12094 1768 12110 1804
rect 12036 1732 12110 1768
rect 12226 1806 12300 1842
rect 12226 1770 12242 1806
rect 12280 1770 12300 1806
rect 12226 1732 12300 1770
rect 12670 -3461 12728 -3449
rect 5383 -4120 5457 -4082
rect 5383 -4156 5403 -4120
rect 5441 -4156 5457 -4120
rect 5383 -4192 5457 -4156
rect 5573 -4118 5647 -4082
rect 5573 -4154 5589 -4118
rect 5627 -4154 5647 -4118
rect 5573 -4192 5647 -4154
rect 5707 -4121 5765 -4083
rect 5707 -4155 5719 -4121
rect 5753 -4155 5765 -4121
rect 5707 -4193 5765 -4155
rect 6565 -4121 6623 -4083
rect 6565 -4155 6577 -4121
rect 6611 -4155 6623 -4121
rect 6565 -4193 6623 -4155
rect 6724 -4122 6798 -4084
rect 6724 -4158 6744 -4122
rect 6782 -4158 6798 -4122
rect 6724 -4194 6798 -4158
rect 6914 -4120 6988 -4084
rect 6914 -4156 6930 -4120
rect 6968 -4156 6988 -4120
rect 6914 -4194 6988 -4156
rect 7094 -4122 7168 -4084
rect 7094 -4158 7114 -4122
rect 7152 -4158 7168 -4122
rect 7094 -4194 7168 -4158
rect 7284 -4120 7358 -4084
rect 7284 -4156 7300 -4120
rect 7338 -4156 7358 -4120
rect 7284 -4194 7358 -4156
rect 7516 -4122 7590 -4084
rect 7516 -4158 7536 -4122
rect 7574 -4158 7590 -4122
rect 7516 -4194 7590 -4158
rect 7706 -4120 7780 -4084
rect 7706 -4156 7722 -4120
rect 7760 -4156 7780 -4120
rect 7706 -4194 7780 -4156
rect 7938 -4122 8012 -4084
rect 7938 -4158 7958 -4122
rect 7996 -4158 8012 -4122
rect 7938 -4194 8012 -4158
rect 8128 -4120 8202 -4084
rect 8128 -4156 8144 -4120
rect 8182 -4156 8202 -4120
rect 8128 -4194 8202 -4156
rect 8377 -4121 8435 -4083
rect 8377 -4155 8389 -4121
rect 8423 -4155 8435 -4121
rect 8377 -4193 8435 -4155
rect 9235 -4121 9293 -4083
rect 9235 -4155 9247 -4121
rect 9281 -4155 9293 -4121
rect 9235 -4193 9293 -4155
rect 9425 -4122 9499 -4084
rect 9425 -4158 9445 -4122
rect 9483 -4158 9499 -4122
rect 9425 -4194 9499 -4158
rect 9615 -4120 9689 -4084
rect 9615 -4156 9631 -4120
rect 9669 -4156 9689 -4120
rect 9615 -4194 9689 -4156
rect 9795 -4122 9869 -4084
rect 9795 -4158 9815 -4122
rect 9853 -4158 9869 -4122
rect 9795 -4194 9869 -4158
rect 9985 -4120 10059 -4084
rect 9985 -4156 10001 -4120
rect 10039 -4156 10059 -4120
rect 9985 -4194 10059 -4156
rect 10217 -4122 10291 -4084
rect 10217 -4158 10237 -4122
rect 10275 -4158 10291 -4122
rect 10217 -4194 10291 -4158
rect 10407 -4120 10481 -4084
rect 10407 -4156 10423 -4120
rect 10461 -4156 10481 -4120
rect 10407 -4194 10481 -4156
rect 10639 -4122 10713 -4084
rect 10639 -4158 10659 -4122
rect 10697 -4158 10713 -4122
rect 10639 -4194 10713 -4158
rect 10829 -4120 10903 -4084
rect 10829 -4156 10845 -4120
rect 10883 -4156 10903 -4120
rect 10829 -4194 10903 -4156
rect 11040 -4120 11098 -4082
rect 11040 -4154 11052 -4120
rect 11086 -4154 11098 -4120
rect 11040 -4192 11098 -4154
rect 11898 -4120 11956 -4082
rect 11898 -4154 11910 -4120
rect 11944 -4154 11956 -4120
rect 11898 -4192 11956 -4154
rect 12670 -3773 12682 -3461
rect 12716 -3773 12728 -3461
rect 12670 -3785 12728 -3773
rect 12758 -3461 12816 -3449
rect 12758 -3773 12770 -3461
rect 12804 -3773 12816 -3461
rect 12758 -3785 12816 -3773
rect 13060 -3463 13118 -3451
rect 13060 -3775 13072 -3463
rect 13106 -3775 13118 -3463
rect 13060 -3787 13118 -3775
rect 13148 -3463 13206 -3451
rect 13148 -3775 13160 -3463
rect 13194 -3775 13206 -3463
rect 13148 -3787 13206 -3775
<< ndiffc >>
rect 397 7162 431 8538
rect 2055 7162 2089 8538
rect 3713 7162 3747 8538
rect 397 5652 431 7028
rect 2055 5652 2089 7028
rect 3713 5652 3747 7028
rect 397 4142 431 5518
rect 2055 4142 2089 5518
rect 3713 4142 3747 5518
rect 397 2632 431 4008
rect 2055 2632 2089 4008
rect 3713 2632 3747 4008
rect 397 1122 431 2498
rect 2055 1122 2089 2498
rect 3713 1122 3747 2498
rect 397 -388 431 988
rect 2055 -388 2089 988
rect 3713 -388 3747 988
rect 397 -1898 431 -522
rect 2055 -1898 2089 -522
rect 3713 -1898 3747 -522
rect 397 -3408 431 -2032
rect 2055 -3408 2089 -2032
rect 3713 -3408 3747 -2032
rect 397 -4918 431 -3542
rect 2055 -4918 2089 -3542
rect 3713 -4918 3747 -3542
rect 397 -6428 431 -5052
rect 2055 -6428 2089 -5052
rect 3713 -6428 3747 -5052
rect 397 -7938 431 -6562
rect 2055 -7938 2089 -6562
rect 3713 -7938 3747 -6562
rect 397 -9448 431 -8072
rect 2055 -9448 2089 -8072
rect 3713 -9448 3747 -8072
rect 5141 6489 5175 6525
rect 5141 6419 5175 6455
rect 5141 6349 5175 6385
rect 5399 6489 5433 6525
rect 5399 6419 5433 6455
rect 5399 6349 5433 6385
rect 5657 6489 5691 6525
rect 5657 6419 5691 6455
rect 5657 6348 5691 6384
rect 5915 6489 5949 6525
rect 5915 6419 5949 6455
rect 5915 6349 5949 6385
rect 6173 6489 6207 6525
rect 6173 6419 6207 6455
rect 6173 6349 6207 6385
rect 6431 6489 6465 6525
rect 6431 6419 6465 6455
rect 6431 6349 6465 6385
rect 6689 6489 6723 6525
rect 6689 6419 6723 6455
rect 6689 6349 6723 6385
rect 6947 6489 6981 6525
rect 6947 6419 6981 6455
rect 6947 6349 6981 6385
rect 7205 6489 7239 6525
rect 7205 6419 7239 6455
rect 7205 6349 7239 6385
rect 7811 6489 7845 6525
rect 7811 6419 7845 6455
rect 7811 6349 7845 6385
rect 8069 6489 8103 6525
rect 8069 6419 8103 6455
rect 8069 6349 8103 6385
rect 8327 6489 8361 6525
rect 8327 6419 8361 6455
rect 8327 6348 8361 6384
rect 8585 6489 8619 6525
rect 8585 6419 8619 6455
rect 8585 6349 8619 6385
rect 8843 6489 8877 6525
rect 8843 6419 8877 6455
rect 8843 6349 8877 6385
rect 9101 6489 9135 6525
rect 9101 6419 9135 6455
rect 9101 6349 9135 6385
rect 9359 6489 9393 6525
rect 9359 6419 9393 6455
rect 9359 6349 9393 6385
rect 9617 6489 9651 6525
rect 9617 6419 9651 6455
rect 9617 6349 9651 6385
rect 9875 6489 9909 6525
rect 9875 6419 9909 6455
rect 9875 6349 9909 6385
rect 10474 6490 10508 6526
rect 10474 6420 10508 6456
rect 10474 6350 10508 6386
rect 10732 6490 10766 6526
rect 10732 6420 10766 6456
rect 10732 6350 10766 6386
rect 10990 6490 11024 6526
rect 10990 6420 11024 6456
rect 10990 6349 11024 6385
rect 11248 6490 11282 6526
rect 11248 6420 11282 6456
rect 11248 6350 11282 6386
rect 11506 6490 11540 6526
rect 11506 6420 11540 6456
rect 11506 6350 11540 6386
rect 11764 6490 11798 6526
rect 11764 6420 11798 6456
rect 11764 6350 11798 6386
rect 12022 6490 12056 6526
rect 12022 6420 12056 6456
rect 12022 6350 12056 6386
rect 12280 6490 12314 6526
rect 12280 6420 12314 6456
rect 12280 6350 12314 6386
rect 12538 6490 12572 6526
rect 12538 6420 12572 6456
rect 12538 6350 12572 6386
rect 5141 6071 5175 6107
rect 5141 6001 5175 6037
rect 5141 5931 5175 5967
rect 5399 6071 5433 6107
rect 5399 6001 5433 6037
rect 5399 5931 5433 5967
rect 5657 6071 5691 6107
rect 5657 6001 5691 6037
rect 5657 5930 5691 5966
rect 5915 6071 5949 6107
rect 5915 6001 5949 6037
rect 5915 5931 5949 5967
rect 6173 6071 6207 6107
rect 6173 6001 6207 6037
rect 6173 5931 6207 5967
rect 6431 6071 6465 6107
rect 6431 6001 6465 6037
rect 6431 5931 6465 5967
rect 6689 6071 6723 6107
rect 6689 6001 6723 6037
rect 6689 5931 6723 5967
rect 6947 6071 6981 6107
rect 6947 6001 6981 6037
rect 6947 5931 6981 5967
rect 7205 6071 7239 6107
rect 7205 6001 7239 6037
rect 7205 5931 7239 5967
rect 7811 6071 7845 6107
rect 7811 6001 7845 6037
rect 7811 5931 7845 5967
rect 8069 6071 8103 6107
rect 8069 6001 8103 6037
rect 8069 5931 8103 5967
rect 8327 6071 8361 6107
rect 8327 6001 8361 6037
rect 8327 5930 8361 5966
rect 8585 6071 8619 6107
rect 8585 6001 8619 6037
rect 8585 5931 8619 5967
rect 8843 6071 8877 6107
rect 8843 6001 8877 6037
rect 8843 5931 8877 5967
rect 9101 6071 9135 6107
rect 9101 6001 9135 6037
rect 9101 5931 9135 5967
rect 9359 6071 9393 6107
rect 9359 6001 9393 6037
rect 9359 5931 9393 5967
rect 9617 6071 9651 6107
rect 9617 6001 9651 6037
rect 9617 5931 9651 5967
rect 9875 6071 9909 6107
rect 9875 6001 9909 6037
rect 9875 5931 9909 5967
rect 10474 6072 10508 6108
rect 10474 6002 10508 6038
rect 10474 5932 10508 5968
rect 10732 6072 10766 6108
rect 10732 6002 10766 6038
rect 10732 5932 10766 5968
rect 10990 6072 11024 6108
rect 10990 6002 11024 6038
rect 10990 5931 11024 5967
rect 11248 6072 11282 6108
rect 11248 6002 11282 6038
rect 11248 5932 11282 5968
rect 11506 6072 11540 6108
rect 11506 6002 11540 6038
rect 11506 5932 11540 5968
rect 11764 6072 11798 6108
rect 11764 6002 11798 6038
rect 11764 5932 11798 5968
rect 12022 6072 12056 6108
rect 12022 6002 12056 6038
rect 12022 5932 12056 5968
rect 12280 6072 12314 6108
rect 12280 6002 12314 6038
rect 12280 5932 12314 5968
rect 12538 6072 12572 6108
rect 12538 6002 12572 6038
rect 12538 5932 12572 5968
rect 5141 5653 5175 5689
rect 5141 5583 5175 5619
rect 5141 5513 5175 5549
rect 5399 5653 5433 5689
rect 5399 5583 5433 5619
rect 5399 5513 5433 5549
rect 5657 5653 5691 5689
rect 5657 5583 5691 5619
rect 5657 5512 5691 5548
rect 5915 5653 5949 5689
rect 5915 5583 5949 5619
rect 5915 5513 5949 5549
rect 6173 5653 6207 5689
rect 6173 5583 6207 5619
rect 6173 5513 6207 5549
rect 6431 5653 6465 5689
rect 6431 5583 6465 5619
rect 6431 5513 6465 5549
rect 6689 5653 6723 5689
rect 6689 5583 6723 5619
rect 6689 5513 6723 5549
rect 6947 5653 6981 5689
rect 6947 5583 6981 5619
rect 6947 5513 6981 5549
rect 7205 5653 7239 5689
rect 7205 5583 7239 5619
rect 7205 5513 7239 5549
rect 7811 5653 7845 5689
rect 7811 5583 7845 5619
rect 7811 5513 7845 5549
rect 8069 5653 8103 5689
rect 8069 5583 8103 5619
rect 8069 5513 8103 5549
rect 8327 5653 8361 5689
rect 8327 5583 8361 5619
rect 8327 5512 8361 5548
rect 8585 5653 8619 5689
rect 8585 5583 8619 5619
rect 8585 5513 8619 5549
rect 8843 5653 8877 5689
rect 8843 5583 8877 5619
rect 8843 5513 8877 5549
rect 9101 5653 9135 5689
rect 9101 5583 9135 5619
rect 9101 5513 9135 5549
rect 9359 5653 9393 5689
rect 9359 5583 9393 5619
rect 9359 5513 9393 5549
rect 9617 5653 9651 5689
rect 9617 5583 9651 5619
rect 9617 5513 9651 5549
rect 9875 5653 9909 5689
rect 9875 5583 9909 5619
rect 9875 5513 9909 5549
rect 10474 5654 10508 5690
rect 10474 5584 10508 5620
rect 10474 5514 10508 5550
rect 10732 5654 10766 5690
rect 10732 5584 10766 5620
rect 10732 5514 10766 5550
rect 10990 5654 11024 5690
rect 10990 5584 11024 5620
rect 10990 5513 11024 5549
rect 11248 5654 11282 5690
rect 11248 5584 11282 5620
rect 11248 5514 11282 5550
rect 11506 5654 11540 5690
rect 11506 5584 11540 5620
rect 11506 5514 11540 5550
rect 11764 5654 11798 5690
rect 11764 5584 11798 5620
rect 11764 5514 11798 5550
rect 12022 5654 12056 5690
rect 12022 5584 12056 5620
rect 12022 5514 12056 5550
rect 12280 5654 12314 5690
rect 12280 5584 12314 5620
rect 12280 5514 12314 5550
rect 12538 5654 12572 5690
rect 12538 5584 12572 5620
rect 12538 5514 12572 5550
rect 5141 5235 5175 5271
rect 5141 5165 5175 5201
rect 5141 5095 5175 5131
rect 5399 5235 5433 5271
rect 5399 5165 5433 5201
rect 5399 5095 5433 5131
rect 5657 5235 5691 5271
rect 5657 5165 5691 5201
rect 5657 5094 5691 5130
rect 5915 5235 5949 5271
rect 5915 5165 5949 5201
rect 5915 5095 5949 5131
rect 6173 5235 6207 5271
rect 6173 5165 6207 5201
rect 6173 5095 6207 5131
rect 6431 5235 6465 5271
rect 6431 5165 6465 5201
rect 6431 5095 6465 5131
rect 6689 5235 6723 5271
rect 6689 5165 6723 5201
rect 6689 5095 6723 5131
rect 6947 5235 6981 5271
rect 6947 5165 6981 5201
rect 6947 5095 6981 5131
rect 7205 5235 7239 5271
rect 7205 5165 7239 5201
rect 7205 5095 7239 5131
rect 7811 5235 7845 5271
rect 7811 5165 7845 5201
rect 7811 5095 7845 5131
rect 8069 5235 8103 5271
rect 8069 5165 8103 5201
rect 8069 5095 8103 5131
rect 8327 5235 8361 5271
rect 8327 5165 8361 5201
rect 8327 5094 8361 5130
rect 8585 5235 8619 5271
rect 8585 5165 8619 5201
rect 8585 5095 8619 5131
rect 8843 5235 8877 5271
rect 8843 5165 8877 5201
rect 8843 5095 8877 5131
rect 9101 5235 9135 5271
rect 9101 5165 9135 5201
rect 9101 5095 9135 5131
rect 9359 5235 9393 5271
rect 9359 5165 9393 5201
rect 9359 5095 9393 5131
rect 9617 5235 9651 5271
rect 9617 5165 9651 5201
rect 9617 5095 9651 5131
rect 9875 5235 9909 5271
rect 9875 5165 9909 5201
rect 9875 5095 9909 5131
rect 10474 5236 10508 5272
rect 10474 5166 10508 5202
rect 10474 5096 10508 5132
rect 10732 5236 10766 5272
rect 10732 5166 10766 5202
rect 10732 5096 10766 5132
rect 10990 5236 11024 5272
rect 10990 5166 11024 5202
rect 10990 5095 11024 5131
rect 11248 5236 11282 5272
rect 11248 5166 11282 5202
rect 11248 5096 11282 5132
rect 11506 5236 11540 5272
rect 11506 5166 11540 5202
rect 11506 5096 11540 5132
rect 11764 5236 11798 5272
rect 11764 5166 11798 5202
rect 11764 5096 11798 5132
rect 12022 5236 12056 5272
rect 12022 5166 12056 5202
rect 12022 5096 12056 5132
rect 12280 5236 12314 5272
rect 12280 5166 12314 5202
rect 12280 5096 12314 5132
rect 12538 5236 12572 5272
rect 12538 5166 12572 5202
rect 12538 5096 12572 5132
rect 5141 4817 5175 4853
rect 5141 4747 5175 4783
rect 5141 4677 5175 4713
rect 5399 4817 5433 4853
rect 5399 4747 5433 4783
rect 5399 4677 5433 4713
rect 5657 4817 5691 4853
rect 5657 4747 5691 4783
rect 5657 4676 5691 4712
rect 5915 4817 5949 4853
rect 5915 4747 5949 4783
rect 5915 4677 5949 4713
rect 6173 4817 6207 4853
rect 6173 4747 6207 4783
rect 6173 4677 6207 4713
rect 6431 4817 6465 4853
rect 6431 4747 6465 4783
rect 6431 4677 6465 4713
rect 6689 4817 6723 4853
rect 6689 4747 6723 4783
rect 6689 4677 6723 4713
rect 6947 4817 6981 4853
rect 6947 4747 6981 4783
rect 6947 4677 6981 4713
rect 7205 4817 7239 4853
rect 7205 4747 7239 4783
rect 7205 4677 7239 4713
rect 7811 4817 7845 4853
rect 7811 4747 7845 4783
rect 7811 4677 7845 4713
rect 8069 4817 8103 4853
rect 8069 4747 8103 4783
rect 8069 4677 8103 4713
rect 8327 4817 8361 4853
rect 8327 4747 8361 4783
rect 8327 4676 8361 4712
rect 8585 4817 8619 4853
rect 8585 4747 8619 4783
rect 8585 4677 8619 4713
rect 8843 4817 8877 4853
rect 8843 4747 8877 4783
rect 8843 4677 8877 4713
rect 9101 4817 9135 4853
rect 9101 4747 9135 4783
rect 9101 4677 9135 4713
rect 9359 4817 9393 4853
rect 9359 4747 9393 4783
rect 9359 4677 9393 4713
rect 9617 4817 9651 4853
rect 9617 4747 9651 4783
rect 9617 4677 9651 4713
rect 9875 4817 9909 4853
rect 9875 4747 9909 4783
rect 9875 4677 9909 4713
rect 10474 4818 10508 4854
rect 10474 4748 10508 4784
rect 10474 4678 10508 4714
rect 10732 4818 10766 4854
rect 10732 4748 10766 4784
rect 10732 4678 10766 4714
rect 10990 4818 11024 4854
rect 10990 4748 11024 4784
rect 10990 4677 11024 4713
rect 11248 4818 11282 4854
rect 11248 4748 11282 4784
rect 11248 4678 11282 4714
rect 11506 4818 11540 4854
rect 11506 4748 11540 4784
rect 11506 4678 11540 4714
rect 11764 4818 11798 4854
rect 11764 4748 11798 4784
rect 11764 4678 11798 4714
rect 12022 4818 12056 4854
rect 12022 4748 12056 4784
rect 12022 4678 12056 4714
rect 12280 4818 12314 4854
rect 12280 4748 12314 4784
rect 12280 4678 12314 4714
rect 12538 4818 12572 4854
rect 12538 4748 12572 4784
rect 12538 4678 12572 4714
rect 5141 4399 5175 4435
rect 5141 4329 5175 4365
rect 5141 4259 5175 4295
rect 5399 4399 5433 4435
rect 5399 4329 5433 4365
rect 5399 4259 5433 4295
rect 5657 4399 5691 4435
rect 5657 4329 5691 4365
rect 5657 4258 5691 4294
rect 5915 4399 5949 4435
rect 5915 4329 5949 4365
rect 5915 4259 5949 4295
rect 6173 4399 6207 4435
rect 6173 4329 6207 4365
rect 6173 4259 6207 4295
rect 6431 4399 6465 4435
rect 6431 4329 6465 4365
rect 6431 4259 6465 4295
rect 6689 4399 6723 4435
rect 6689 4329 6723 4365
rect 6689 4259 6723 4295
rect 6947 4399 6981 4435
rect 6947 4329 6981 4365
rect 6947 4259 6981 4295
rect 7205 4399 7239 4435
rect 7205 4329 7239 4365
rect 7205 4259 7239 4295
rect 7811 4399 7845 4435
rect 7811 4329 7845 4365
rect 7811 4259 7845 4295
rect 8069 4399 8103 4435
rect 8069 4329 8103 4365
rect 8069 4259 8103 4295
rect 8327 4399 8361 4435
rect 8327 4329 8361 4365
rect 8327 4258 8361 4294
rect 8585 4399 8619 4435
rect 8585 4329 8619 4365
rect 8585 4259 8619 4295
rect 8843 4399 8877 4435
rect 8843 4329 8877 4365
rect 8843 4259 8877 4295
rect 9101 4399 9135 4435
rect 9101 4329 9135 4365
rect 9101 4259 9135 4295
rect 9359 4399 9393 4435
rect 9359 4329 9393 4365
rect 9359 4259 9393 4295
rect 9617 4399 9651 4435
rect 9617 4329 9651 4365
rect 9617 4259 9651 4295
rect 9875 4399 9909 4435
rect 9875 4329 9909 4365
rect 9875 4259 9909 4295
rect 10474 4400 10508 4436
rect 10474 4330 10508 4366
rect 10474 4260 10508 4296
rect 10732 4400 10766 4436
rect 10732 4330 10766 4366
rect 10732 4260 10766 4296
rect 10990 4400 11024 4436
rect 10990 4330 11024 4366
rect 10990 4259 11024 4295
rect 11248 4400 11282 4436
rect 11248 4330 11282 4366
rect 11248 4260 11282 4296
rect 11506 4400 11540 4436
rect 11506 4330 11540 4366
rect 11506 4260 11540 4296
rect 11764 4400 11798 4436
rect 11764 4330 11798 4366
rect 11764 4260 11798 4296
rect 12022 4400 12056 4436
rect 12022 4330 12056 4366
rect 12022 4260 12056 4296
rect 12280 4400 12314 4436
rect 12280 4330 12314 4366
rect 12280 4260 12314 4296
rect 12538 4400 12572 4436
rect 12538 4330 12572 4366
rect 12538 4260 12572 4296
rect 5141 3981 5175 4017
rect 5141 3911 5175 3947
rect 5141 3841 5175 3877
rect 5399 3981 5433 4017
rect 5399 3911 5433 3947
rect 5399 3841 5433 3877
rect 5657 3981 5691 4017
rect 5657 3911 5691 3947
rect 5657 3840 5691 3876
rect 5915 3981 5949 4017
rect 5915 3911 5949 3947
rect 5915 3841 5949 3877
rect 6173 3981 6207 4017
rect 6173 3911 6207 3947
rect 6173 3841 6207 3877
rect 6431 3981 6465 4017
rect 6431 3911 6465 3947
rect 6431 3841 6465 3877
rect 6689 3981 6723 4017
rect 6689 3911 6723 3947
rect 6689 3841 6723 3877
rect 6947 3981 6981 4017
rect 6947 3911 6981 3947
rect 6947 3841 6981 3877
rect 7205 3981 7239 4017
rect 7205 3911 7239 3947
rect 7205 3841 7239 3877
rect 7811 3981 7845 4017
rect 7811 3911 7845 3947
rect 7811 3841 7845 3877
rect 8069 3981 8103 4017
rect 8069 3911 8103 3947
rect 8069 3841 8103 3877
rect 8327 3981 8361 4017
rect 8327 3911 8361 3947
rect 8327 3840 8361 3876
rect 8585 3981 8619 4017
rect 8585 3911 8619 3947
rect 8585 3841 8619 3877
rect 8843 3981 8877 4017
rect 8843 3911 8877 3947
rect 8843 3841 8877 3877
rect 9101 3981 9135 4017
rect 9101 3911 9135 3947
rect 9101 3841 9135 3877
rect 9359 3981 9393 4017
rect 9359 3911 9393 3947
rect 9359 3841 9393 3877
rect 9617 3981 9651 4017
rect 9617 3911 9651 3947
rect 9617 3841 9651 3877
rect 9875 3981 9909 4017
rect 9875 3911 9909 3947
rect 9875 3841 9909 3877
rect 10474 3982 10508 4018
rect 10474 3912 10508 3948
rect 10474 3842 10508 3878
rect 10732 3982 10766 4018
rect 10732 3912 10766 3948
rect 10732 3842 10766 3878
rect 10990 3982 11024 4018
rect 10990 3912 11024 3948
rect 10990 3841 11024 3877
rect 11248 3982 11282 4018
rect 11248 3912 11282 3948
rect 11248 3842 11282 3878
rect 11506 3982 11540 4018
rect 11506 3912 11540 3948
rect 11506 3842 11540 3878
rect 11764 3982 11798 4018
rect 11764 3912 11798 3948
rect 11764 3842 11798 3878
rect 12022 3982 12056 4018
rect 12022 3912 12056 3948
rect 12022 3842 12056 3878
rect 12280 3982 12314 4018
rect 12280 3912 12314 3948
rect 12280 3842 12314 3878
rect 12538 3982 12572 4018
rect 12538 3912 12572 3948
rect 12538 3842 12572 3878
rect 5021 3329 5055 3363
rect 5021 3259 5055 3295
rect 5021 3191 5055 3225
rect 5279 3329 5313 3363
rect 5279 3259 5313 3295
rect 5279 3191 5313 3225
rect 5561 3329 5595 3363
rect 5561 3259 5595 3295
rect 5561 3191 5595 3225
rect 5819 3329 5853 3363
rect 5819 3259 5853 3295
rect 5819 3191 5853 3225
rect 6041 3329 6075 3363
rect 6041 3259 6075 3295
rect 6041 3191 6075 3225
rect 6299 3329 6333 3363
rect 6299 3259 6333 3295
rect 6299 3191 6333 3225
rect 6544 3331 6578 3365
rect 6544 3261 6578 3297
rect 6544 3193 6578 3227
rect 6802 3331 6836 3365
rect 6802 3261 6836 3297
rect 6802 3193 6836 3227
rect 7054 3341 7088 3375
rect 7054 3271 7088 3307
rect 7054 3203 7088 3237
rect 7312 3341 7346 3375
rect 7312 3271 7346 3307
rect 7312 3203 7346 3237
rect 7691 3329 7725 3363
rect 7691 3259 7725 3295
rect 7691 3191 7725 3225
rect 7949 3329 7983 3363
rect 7949 3259 7983 3295
rect 7949 3191 7983 3225
rect 8231 3329 8265 3363
rect 8231 3259 8265 3295
rect 8231 3191 8265 3225
rect 8489 3329 8523 3363
rect 8489 3259 8523 3295
rect 8489 3191 8523 3225
rect 8711 3329 8745 3363
rect 8711 3259 8745 3295
rect 8711 3191 8745 3225
rect 8969 3329 9003 3363
rect 8969 3259 9003 3295
rect 8969 3191 9003 3225
rect 9214 3331 9248 3365
rect 9214 3261 9248 3297
rect 9214 3193 9248 3227
rect 9472 3331 9506 3365
rect 9472 3261 9506 3297
rect 9472 3193 9506 3227
rect 9724 3341 9758 3375
rect 9724 3271 9758 3307
rect 9724 3203 9758 3237
rect 9982 3341 10016 3375
rect 9982 3271 10016 3307
rect 9982 3203 10016 3237
rect 10354 3330 10388 3364
rect 10354 3260 10388 3296
rect 10354 3192 10388 3226
rect 10612 3330 10646 3364
rect 10612 3260 10646 3296
rect 10612 3192 10646 3226
rect 10894 3330 10928 3364
rect 10894 3260 10928 3296
rect 10894 3192 10928 3226
rect 11152 3330 11186 3364
rect 11152 3260 11186 3296
rect 11152 3192 11186 3226
rect 11374 3330 11408 3364
rect 11374 3260 11408 3296
rect 11374 3192 11408 3226
rect 11632 3330 11666 3364
rect 11632 3260 11666 3296
rect 11632 3192 11666 3226
rect 11877 3332 11911 3366
rect 11877 3262 11911 3298
rect 11877 3194 11911 3228
rect 12135 3332 12169 3366
rect 12135 3262 12169 3298
rect 12135 3194 12169 3228
rect 12387 3342 12421 3376
rect 12387 3272 12421 3308
rect 12387 3204 12421 3238
rect 12645 3342 12679 3376
rect 12645 3272 12679 3308
rect 12645 3204 12679 3238
rect 5141 772 5175 808
rect 5141 702 5175 738
rect 5141 632 5175 668
rect 5399 772 5433 808
rect 5399 702 5433 738
rect 5399 632 5433 668
rect 5657 772 5691 808
rect 5657 702 5691 738
rect 5657 631 5691 667
rect 5915 772 5949 808
rect 5915 702 5949 738
rect 5915 632 5949 668
rect 6173 772 6207 808
rect 6173 702 6207 738
rect 6173 632 6207 668
rect 6431 772 6465 808
rect 6431 702 6465 738
rect 6431 632 6465 668
rect 6689 772 6723 808
rect 6689 702 6723 738
rect 6689 632 6723 668
rect 6947 772 6981 808
rect 6947 702 6981 738
rect 6947 632 6981 668
rect 7205 772 7239 808
rect 7205 702 7239 738
rect 7205 632 7239 668
rect 7811 772 7845 808
rect 7811 702 7845 738
rect 7811 632 7845 668
rect 8069 772 8103 808
rect 8069 702 8103 738
rect 8069 632 8103 668
rect 8327 772 8361 808
rect 8327 702 8361 738
rect 8327 631 8361 667
rect 8585 772 8619 808
rect 8585 702 8619 738
rect 8585 632 8619 668
rect 8843 772 8877 808
rect 8843 702 8877 738
rect 8843 632 8877 668
rect 9101 772 9135 808
rect 9101 702 9135 738
rect 9101 632 9135 668
rect 9359 772 9393 808
rect 9359 702 9393 738
rect 9359 632 9393 668
rect 9617 772 9651 808
rect 9617 702 9651 738
rect 9617 632 9651 668
rect 9875 772 9909 808
rect 9875 702 9909 738
rect 9875 632 9909 668
rect 10474 773 10508 809
rect 10474 703 10508 739
rect 10474 633 10508 669
rect 10732 773 10766 809
rect 10732 703 10766 739
rect 10732 633 10766 669
rect 10990 773 11024 809
rect 10990 703 11024 739
rect 10990 632 11024 668
rect 11248 773 11282 809
rect 11248 703 11282 739
rect 11248 633 11282 669
rect 11506 773 11540 809
rect 11506 703 11540 739
rect 11506 633 11540 669
rect 11764 773 11798 809
rect 11764 703 11798 739
rect 11764 633 11798 669
rect 12022 773 12056 809
rect 12022 703 12056 739
rect 12022 633 12056 669
rect 12280 773 12314 809
rect 12280 703 12314 739
rect 12280 633 12314 669
rect 12538 773 12572 809
rect 12538 703 12572 739
rect 12538 633 12572 669
rect 5141 354 5175 390
rect 5141 284 5175 320
rect 5141 214 5175 250
rect 5399 354 5433 390
rect 5399 284 5433 320
rect 5399 214 5433 250
rect 5657 354 5691 390
rect 5657 284 5691 320
rect 5657 213 5691 249
rect 5915 354 5949 390
rect 5915 284 5949 320
rect 5915 214 5949 250
rect 6173 354 6207 390
rect 6173 284 6207 320
rect 6173 214 6207 250
rect 6431 354 6465 390
rect 6431 284 6465 320
rect 6431 214 6465 250
rect 6689 354 6723 390
rect 6689 284 6723 320
rect 6689 214 6723 250
rect 6947 354 6981 390
rect 6947 284 6981 320
rect 6947 214 6981 250
rect 7205 354 7239 390
rect 7205 284 7239 320
rect 7205 214 7239 250
rect 7811 354 7845 390
rect 7811 284 7845 320
rect 7811 214 7845 250
rect 8069 354 8103 390
rect 8069 284 8103 320
rect 8069 214 8103 250
rect 8327 354 8361 390
rect 8327 284 8361 320
rect 8327 213 8361 249
rect 8585 354 8619 390
rect 8585 284 8619 320
rect 8585 214 8619 250
rect 8843 354 8877 390
rect 8843 284 8877 320
rect 8843 214 8877 250
rect 9101 354 9135 390
rect 9101 284 9135 320
rect 9101 214 9135 250
rect 9359 354 9393 390
rect 9359 284 9393 320
rect 9359 214 9393 250
rect 9617 354 9651 390
rect 9617 284 9651 320
rect 9617 214 9651 250
rect 9875 354 9909 390
rect 9875 284 9909 320
rect 9875 214 9909 250
rect 10474 355 10508 391
rect 10474 285 10508 321
rect 10474 215 10508 251
rect 10732 355 10766 391
rect 10732 285 10766 321
rect 10732 215 10766 251
rect 10990 355 11024 391
rect 10990 285 11024 321
rect 10990 214 11024 250
rect 11248 355 11282 391
rect 11248 285 11282 321
rect 11248 215 11282 251
rect 11506 355 11540 391
rect 11506 285 11540 321
rect 11506 215 11540 251
rect 11764 355 11798 391
rect 11764 285 11798 321
rect 11764 215 11798 251
rect 12022 355 12056 391
rect 12022 285 12056 321
rect 12022 215 12056 251
rect 12280 355 12314 391
rect 12280 285 12314 321
rect 12280 215 12314 251
rect 12538 355 12572 391
rect 12538 285 12572 321
rect 12538 215 12572 251
rect 5141 -64 5175 -28
rect 5141 -134 5175 -98
rect 5141 -204 5175 -168
rect 5399 -64 5433 -28
rect 5399 -134 5433 -98
rect 5399 -204 5433 -168
rect 5657 -64 5691 -28
rect 5657 -134 5691 -98
rect 5657 -205 5691 -169
rect 5915 -64 5949 -28
rect 5915 -134 5949 -98
rect 5915 -204 5949 -168
rect 6173 -64 6207 -28
rect 6173 -134 6207 -98
rect 6173 -204 6207 -168
rect 6431 -64 6465 -28
rect 6431 -134 6465 -98
rect 6431 -204 6465 -168
rect 6689 -64 6723 -28
rect 6689 -134 6723 -98
rect 6689 -204 6723 -168
rect 6947 -64 6981 -28
rect 6947 -134 6981 -98
rect 6947 -204 6981 -168
rect 7205 -64 7239 -28
rect 7205 -134 7239 -98
rect 7205 -204 7239 -168
rect 7811 -64 7845 -28
rect 7811 -134 7845 -98
rect 7811 -204 7845 -168
rect 8069 -64 8103 -28
rect 8069 -134 8103 -98
rect 8069 -204 8103 -168
rect 8327 -64 8361 -28
rect 8327 -134 8361 -98
rect 8327 -205 8361 -169
rect 8585 -64 8619 -28
rect 8585 -134 8619 -98
rect 8585 -204 8619 -168
rect 8843 -64 8877 -28
rect 8843 -134 8877 -98
rect 8843 -204 8877 -168
rect 9101 -64 9135 -28
rect 9101 -134 9135 -98
rect 9101 -204 9135 -168
rect 9359 -64 9393 -28
rect 9359 -134 9393 -98
rect 9359 -204 9393 -168
rect 9617 -64 9651 -28
rect 9617 -134 9651 -98
rect 9617 -204 9651 -168
rect 9875 -64 9909 -28
rect 9875 -134 9909 -98
rect 9875 -204 9909 -168
rect 10474 -63 10508 -27
rect 10474 -133 10508 -97
rect 10474 -203 10508 -167
rect 10732 -63 10766 -27
rect 10732 -133 10766 -97
rect 10732 -203 10766 -167
rect 10990 -63 11024 -27
rect 10990 -133 11024 -97
rect 10990 -204 11024 -168
rect 11248 -63 11282 -27
rect 11248 -133 11282 -97
rect 11248 -203 11282 -167
rect 11506 -63 11540 -27
rect 11506 -133 11540 -97
rect 11506 -203 11540 -167
rect 11764 -63 11798 -27
rect 11764 -133 11798 -97
rect 11764 -203 11798 -167
rect 12022 -63 12056 -27
rect 12022 -133 12056 -97
rect 12022 -203 12056 -167
rect 12280 -63 12314 -27
rect 12280 -133 12314 -97
rect 12280 -203 12314 -167
rect 12538 -63 12572 -27
rect 12538 -133 12572 -97
rect 12538 -203 12572 -167
rect 5141 -482 5175 -446
rect 5141 -552 5175 -516
rect 5141 -622 5175 -586
rect 5399 -482 5433 -446
rect 5399 -552 5433 -516
rect 5399 -622 5433 -586
rect 5657 -482 5691 -446
rect 5657 -552 5691 -516
rect 5657 -623 5691 -587
rect 5915 -482 5949 -446
rect 5915 -552 5949 -516
rect 5915 -622 5949 -586
rect 6173 -482 6207 -446
rect 6173 -552 6207 -516
rect 6173 -622 6207 -586
rect 6431 -482 6465 -446
rect 6431 -552 6465 -516
rect 6431 -622 6465 -586
rect 6689 -482 6723 -446
rect 6689 -552 6723 -516
rect 6689 -622 6723 -586
rect 6947 -482 6981 -446
rect 6947 -552 6981 -516
rect 6947 -622 6981 -586
rect 7205 -482 7239 -446
rect 7205 -552 7239 -516
rect 7205 -622 7239 -586
rect 7811 -482 7845 -446
rect 7811 -552 7845 -516
rect 7811 -622 7845 -586
rect 8069 -482 8103 -446
rect 8069 -552 8103 -516
rect 8069 -622 8103 -586
rect 8327 -482 8361 -446
rect 8327 -552 8361 -516
rect 8327 -623 8361 -587
rect 8585 -482 8619 -446
rect 8585 -552 8619 -516
rect 8585 -622 8619 -586
rect 8843 -482 8877 -446
rect 8843 -552 8877 -516
rect 8843 -622 8877 -586
rect 9101 -482 9135 -446
rect 9101 -552 9135 -516
rect 9101 -622 9135 -586
rect 9359 -482 9393 -446
rect 9359 -552 9393 -516
rect 9359 -622 9393 -586
rect 9617 -482 9651 -446
rect 9617 -552 9651 -516
rect 9617 -622 9651 -586
rect 9875 -482 9909 -446
rect 9875 -552 9909 -516
rect 9875 -622 9909 -586
rect 10474 -481 10508 -445
rect 10474 -551 10508 -515
rect 10474 -621 10508 -585
rect 10732 -481 10766 -445
rect 10732 -551 10766 -515
rect 10732 -621 10766 -585
rect 10990 -481 11024 -445
rect 10990 -551 11024 -515
rect 10990 -622 11024 -586
rect 11248 -481 11282 -445
rect 11248 -551 11282 -515
rect 11248 -621 11282 -585
rect 11506 -481 11540 -445
rect 11506 -551 11540 -515
rect 11506 -621 11540 -585
rect 11764 -481 11798 -445
rect 11764 -551 11798 -515
rect 11764 -621 11798 -585
rect 12022 -481 12056 -445
rect 12022 -551 12056 -515
rect 12022 -621 12056 -585
rect 12280 -481 12314 -445
rect 12280 -551 12314 -515
rect 12280 -621 12314 -585
rect 12538 -481 12572 -445
rect 12538 -551 12572 -515
rect 12538 -621 12572 -585
rect 5141 -900 5175 -864
rect 5141 -970 5175 -934
rect 5141 -1040 5175 -1004
rect 5399 -900 5433 -864
rect 5399 -970 5433 -934
rect 5399 -1040 5433 -1004
rect 5657 -900 5691 -864
rect 5657 -970 5691 -934
rect 5657 -1041 5691 -1005
rect 5915 -900 5949 -864
rect 5915 -970 5949 -934
rect 5915 -1040 5949 -1004
rect 6173 -900 6207 -864
rect 6173 -970 6207 -934
rect 6173 -1040 6207 -1004
rect 6431 -900 6465 -864
rect 6431 -970 6465 -934
rect 6431 -1040 6465 -1004
rect 6689 -900 6723 -864
rect 6689 -970 6723 -934
rect 6689 -1040 6723 -1004
rect 6947 -900 6981 -864
rect 6947 -970 6981 -934
rect 6947 -1040 6981 -1004
rect 7205 -900 7239 -864
rect 7205 -970 7239 -934
rect 7205 -1040 7239 -1004
rect 7811 -900 7845 -864
rect 7811 -970 7845 -934
rect 7811 -1040 7845 -1004
rect 8069 -900 8103 -864
rect 8069 -970 8103 -934
rect 8069 -1040 8103 -1004
rect 8327 -900 8361 -864
rect 8327 -970 8361 -934
rect 8327 -1041 8361 -1005
rect 8585 -900 8619 -864
rect 8585 -970 8619 -934
rect 8585 -1040 8619 -1004
rect 8843 -900 8877 -864
rect 8843 -970 8877 -934
rect 8843 -1040 8877 -1004
rect 9101 -900 9135 -864
rect 9101 -970 9135 -934
rect 9101 -1040 9135 -1004
rect 9359 -900 9393 -864
rect 9359 -970 9393 -934
rect 9359 -1040 9393 -1004
rect 9617 -900 9651 -864
rect 9617 -970 9651 -934
rect 9617 -1040 9651 -1004
rect 9875 -900 9909 -864
rect 9875 -970 9909 -934
rect 9875 -1040 9909 -1004
rect 10474 -899 10508 -863
rect 10474 -969 10508 -933
rect 10474 -1039 10508 -1003
rect 10732 -899 10766 -863
rect 10732 -969 10766 -933
rect 10732 -1039 10766 -1003
rect 10990 -899 11024 -863
rect 10990 -969 11024 -933
rect 10990 -1040 11024 -1004
rect 11248 -899 11282 -863
rect 11248 -969 11282 -933
rect 11248 -1039 11282 -1003
rect 11506 -899 11540 -863
rect 11506 -969 11540 -933
rect 11506 -1039 11540 -1003
rect 11764 -899 11798 -863
rect 11764 -969 11798 -933
rect 11764 -1039 11798 -1003
rect 12022 -899 12056 -863
rect 12022 -969 12056 -933
rect 12022 -1039 12056 -1003
rect 12280 -899 12314 -863
rect 12280 -969 12314 -933
rect 12280 -1039 12314 -1003
rect 12538 -899 12572 -863
rect 12538 -969 12572 -933
rect 12538 -1039 12572 -1003
rect 5141 -1318 5175 -1282
rect 5141 -1388 5175 -1352
rect 5141 -1458 5175 -1422
rect 5399 -1318 5433 -1282
rect 5399 -1388 5433 -1352
rect 5399 -1458 5433 -1422
rect 5657 -1318 5691 -1282
rect 5657 -1388 5691 -1352
rect 5657 -1459 5691 -1423
rect 5915 -1318 5949 -1282
rect 5915 -1388 5949 -1352
rect 5915 -1458 5949 -1422
rect 6173 -1318 6207 -1282
rect 6173 -1388 6207 -1352
rect 6173 -1458 6207 -1422
rect 6431 -1318 6465 -1282
rect 6431 -1388 6465 -1352
rect 6431 -1458 6465 -1422
rect 6689 -1318 6723 -1282
rect 6689 -1388 6723 -1352
rect 6689 -1458 6723 -1422
rect 6947 -1318 6981 -1282
rect 6947 -1388 6981 -1352
rect 6947 -1458 6981 -1422
rect 7205 -1318 7239 -1282
rect 7205 -1388 7239 -1352
rect 7205 -1458 7239 -1422
rect 7811 -1318 7845 -1282
rect 7811 -1388 7845 -1352
rect 7811 -1458 7845 -1422
rect 8069 -1318 8103 -1282
rect 8069 -1388 8103 -1352
rect 8069 -1458 8103 -1422
rect 8327 -1318 8361 -1282
rect 8327 -1388 8361 -1352
rect 8327 -1459 8361 -1423
rect 8585 -1318 8619 -1282
rect 8585 -1388 8619 -1352
rect 8585 -1458 8619 -1422
rect 8843 -1318 8877 -1282
rect 8843 -1388 8877 -1352
rect 8843 -1458 8877 -1422
rect 9101 -1318 9135 -1282
rect 9101 -1388 9135 -1352
rect 9101 -1458 9135 -1422
rect 9359 -1318 9393 -1282
rect 9359 -1388 9393 -1352
rect 9359 -1458 9393 -1422
rect 9617 -1318 9651 -1282
rect 9617 -1388 9651 -1352
rect 9617 -1458 9651 -1422
rect 9875 -1318 9909 -1282
rect 9875 -1388 9909 -1352
rect 9875 -1458 9909 -1422
rect 10474 -1317 10508 -1281
rect 10474 -1387 10508 -1351
rect 10474 -1457 10508 -1421
rect 10732 -1317 10766 -1281
rect 10732 -1387 10766 -1351
rect 10732 -1457 10766 -1421
rect 10990 -1317 11024 -1281
rect 10990 -1387 11024 -1351
rect 10990 -1458 11024 -1422
rect 11248 -1317 11282 -1281
rect 11248 -1387 11282 -1351
rect 11248 -1457 11282 -1421
rect 11506 -1317 11540 -1281
rect 11506 -1387 11540 -1351
rect 11506 -1457 11540 -1421
rect 11764 -1317 11798 -1281
rect 11764 -1387 11798 -1351
rect 11764 -1457 11798 -1421
rect 12022 -1317 12056 -1281
rect 12022 -1387 12056 -1351
rect 12022 -1457 12056 -1421
rect 12280 -1317 12314 -1281
rect 12280 -1387 12314 -1351
rect 12280 -1457 12314 -1421
rect 12538 -1317 12572 -1281
rect 12538 -1387 12572 -1351
rect 12538 -1457 12572 -1421
rect 5141 -1736 5175 -1700
rect 5141 -1806 5175 -1770
rect 5141 -1876 5175 -1840
rect 5399 -1736 5433 -1700
rect 5399 -1806 5433 -1770
rect 5399 -1876 5433 -1840
rect 5657 -1736 5691 -1700
rect 5657 -1806 5691 -1770
rect 5657 -1877 5691 -1841
rect 5915 -1736 5949 -1700
rect 5915 -1806 5949 -1770
rect 5915 -1876 5949 -1840
rect 6173 -1736 6207 -1700
rect 6173 -1806 6207 -1770
rect 6173 -1876 6207 -1840
rect 6431 -1736 6465 -1700
rect 6431 -1806 6465 -1770
rect 6431 -1876 6465 -1840
rect 6689 -1736 6723 -1700
rect 6689 -1806 6723 -1770
rect 6689 -1876 6723 -1840
rect 6947 -1736 6981 -1700
rect 6947 -1806 6981 -1770
rect 6947 -1876 6981 -1840
rect 7205 -1736 7239 -1700
rect 7205 -1806 7239 -1770
rect 7205 -1876 7239 -1840
rect 7811 -1736 7845 -1700
rect 7811 -1806 7845 -1770
rect 7811 -1876 7845 -1840
rect 8069 -1736 8103 -1700
rect 8069 -1806 8103 -1770
rect 8069 -1876 8103 -1840
rect 8327 -1736 8361 -1700
rect 8327 -1806 8361 -1770
rect 8327 -1877 8361 -1841
rect 8585 -1736 8619 -1700
rect 8585 -1806 8619 -1770
rect 8585 -1876 8619 -1840
rect 8843 -1736 8877 -1700
rect 8843 -1806 8877 -1770
rect 8843 -1876 8877 -1840
rect 9101 -1736 9135 -1700
rect 9101 -1806 9135 -1770
rect 9101 -1876 9135 -1840
rect 9359 -1736 9393 -1700
rect 9359 -1806 9393 -1770
rect 9359 -1876 9393 -1840
rect 9617 -1736 9651 -1700
rect 9617 -1806 9651 -1770
rect 9617 -1876 9651 -1840
rect 9875 -1736 9909 -1700
rect 9875 -1806 9909 -1770
rect 9875 -1876 9909 -1840
rect 10474 -1735 10508 -1699
rect 10474 -1805 10508 -1769
rect 10474 -1875 10508 -1839
rect 10732 -1735 10766 -1699
rect 10732 -1805 10766 -1769
rect 10732 -1875 10766 -1839
rect 10990 -1735 11024 -1699
rect 10990 -1805 11024 -1769
rect 10990 -1876 11024 -1840
rect 11248 -1735 11282 -1699
rect 11248 -1805 11282 -1769
rect 11248 -1875 11282 -1839
rect 11506 -1735 11540 -1699
rect 11506 -1805 11540 -1769
rect 11506 -1875 11540 -1839
rect 11764 -1735 11798 -1699
rect 11764 -1805 11798 -1769
rect 11764 -1875 11798 -1839
rect 12022 -1735 12056 -1699
rect 12022 -1805 12056 -1769
rect 12022 -1875 12056 -1839
rect 12280 -1735 12314 -1699
rect 12280 -1805 12314 -1769
rect 12280 -1875 12314 -1839
rect 12538 -1735 12572 -1699
rect 12538 -1805 12572 -1769
rect 12538 -1875 12572 -1839
rect 5021 -2388 5055 -2354
rect 5021 -2458 5055 -2422
rect 5021 -2526 5055 -2492
rect 5279 -2388 5313 -2354
rect 5279 -2458 5313 -2422
rect 5279 -2526 5313 -2492
rect 5561 -2388 5595 -2354
rect 5561 -2458 5595 -2422
rect 5561 -2526 5595 -2492
rect 5819 -2388 5853 -2354
rect 5819 -2458 5853 -2422
rect 5819 -2526 5853 -2492
rect 6041 -2388 6075 -2354
rect 6041 -2458 6075 -2422
rect 6041 -2526 6075 -2492
rect 6299 -2388 6333 -2354
rect 6299 -2458 6333 -2422
rect 6299 -2526 6333 -2492
rect 6544 -2386 6578 -2352
rect 6544 -2456 6578 -2420
rect 6544 -2524 6578 -2490
rect 6802 -2386 6836 -2352
rect 6802 -2456 6836 -2420
rect 6802 -2524 6836 -2490
rect 7054 -2376 7088 -2342
rect 7054 -2446 7088 -2410
rect 7054 -2514 7088 -2480
rect 7312 -2376 7346 -2342
rect 7312 -2446 7346 -2410
rect 7312 -2514 7346 -2480
rect 7691 -2388 7725 -2354
rect 7691 -2458 7725 -2422
rect 7691 -2526 7725 -2492
rect 7949 -2388 7983 -2354
rect 7949 -2458 7983 -2422
rect 7949 -2526 7983 -2492
rect 8231 -2388 8265 -2354
rect 8231 -2458 8265 -2422
rect 8231 -2526 8265 -2492
rect 8489 -2388 8523 -2354
rect 8489 -2458 8523 -2422
rect 8489 -2526 8523 -2492
rect 8711 -2388 8745 -2354
rect 8711 -2458 8745 -2422
rect 8711 -2526 8745 -2492
rect 8969 -2388 9003 -2354
rect 8969 -2458 9003 -2422
rect 8969 -2526 9003 -2492
rect 9214 -2386 9248 -2352
rect 9214 -2456 9248 -2420
rect 9214 -2524 9248 -2490
rect 9472 -2386 9506 -2352
rect 9472 -2456 9506 -2420
rect 9472 -2524 9506 -2490
rect 9724 -2376 9758 -2342
rect 9724 -2446 9758 -2410
rect 9724 -2514 9758 -2480
rect 9982 -2376 10016 -2342
rect 9982 -2446 10016 -2410
rect 9982 -2514 10016 -2480
rect 10354 -2387 10388 -2353
rect 10354 -2457 10388 -2421
rect 10354 -2525 10388 -2491
rect 10612 -2387 10646 -2353
rect 10612 -2457 10646 -2421
rect 10612 -2525 10646 -2491
rect 10894 -2387 10928 -2353
rect 10894 -2457 10928 -2421
rect 10894 -2525 10928 -2491
rect 11152 -2387 11186 -2353
rect 11152 -2457 11186 -2421
rect 11152 -2525 11186 -2491
rect 11374 -2387 11408 -2353
rect 11374 -2457 11408 -2421
rect 11374 -2525 11408 -2491
rect 11632 -2387 11666 -2353
rect 11632 -2457 11666 -2421
rect 11632 -2525 11666 -2491
rect 11877 -2385 11911 -2351
rect 11877 -2455 11911 -2419
rect 11877 -2523 11911 -2489
rect 12135 -2385 12169 -2351
rect 12135 -2455 12169 -2419
rect 12135 -2523 12169 -2489
rect 12387 -2375 12421 -2341
rect 12387 -2445 12421 -2409
rect 12387 -2513 12421 -2479
rect 12645 -2375 12679 -2341
rect 12645 -2445 12679 -2409
rect 12645 -2513 12679 -2479
rect 12686 -4308 12720 -4248
rect 12774 -4308 12808 -4248
rect 13076 -4308 13110 -4248
rect 13164 -4308 13198 -4248
rect 5141 -5132 5175 -5096
rect 5141 -5202 5175 -5166
rect 5141 -5272 5175 -5236
rect 5399 -5132 5433 -5096
rect 5399 -5202 5433 -5166
rect 5399 -5272 5433 -5236
rect 5657 -5132 5691 -5096
rect 5657 -5202 5691 -5166
rect 5657 -5273 5691 -5237
rect 5915 -5132 5949 -5096
rect 5915 -5202 5949 -5166
rect 5915 -5272 5949 -5236
rect 6173 -5132 6207 -5096
rect 6173 -5202 6207 -5166
rect 6173 -5272 6207 -5236
rect 6431 -5132 6465 -5096
rect 6431 -5202 6465 -5166
rect 6431 -5272 6465 -5236
rect 6689 -5132 6723 -5096
rect 6689 -5202 6723 -5166
rect 6689 -5272 6723 -5236
rect 6947 -5132 6981 -5096
rect 6947 -5202 6981 -5166
rect 6947 -5272 6981 -5236
rect 7205 -5132 7239 -5096
rect 7205 -5202 7239 -5166
rect 7205 -5272 7239 -5236
rect 7811 -5132 7845 -5096
rect 7811 -5202 7845 -5166
rect 7811 -5272 7845 -5236
rect 8069 -5132 8103 -5096
rect 8069 -5202 8103 -5166
rect 8069 -5272 8103 -5236
rect 8327 -5132 8361 -5096
rect 8327 -5202 8361 -5166
rect 8327 -5273 8361 -5237
rect 8585 -5132 8619 -5096
rect 8585 -5202 8619 -5166
rect 8585 -5272 8619 -5236
rect 8843 -5132 8877 -5096
rect 8843 -5202 8877 -5166
rect 8843 -5272 8877 -5236
rect 9101 -5132 9135 -5096
rect 9101 -5202 9135 -5166
rect 9101 -5272 9135 -5236
rect 9359 -5132 9393 -5096
rect 9359 -5202 9393 -5166
rect 9359 -5272 9393 -5236
rect 9617 -5132 9651 -5096
rect 9617 -5202 9651 -5166
rect 9617 -5272 9651 -5236
rect 9875 -5132 9909 -5096
rect 9875 -5202 9909 -5166
rect 9875 -5272 9909 -5236
rect 10474 -5131 10508 -5095
rect 10474 -5201 10508 -5165
rect 10474 -5271 10508 -5235
rect 10732 -5131 10766 -5095
rect 10732 -5201 10766 -5165
rect 10732 -5271 10766 -5235
rect 10990 -5131 11024 -5095
rect 10990 -5201 11024 -5165
rect 10990 -5272 11024 -5236
rect 11248 -5131 11282 -5095
rect 11248 -5201 11282 -5165
rect 11248 -5271 11282 -5235
rect 11506 -5131 11540 -5095
rect 11506 -5201 11540 -5165
rect 11506 -5271 11540 -5235
rect 11764 -5131 11798 -5095
rect 11764 -5201 11798 -5165
rect 11764 -5271 11798 -5235
rect 12022 -5131 12056 -5095
rect 12022 -5201 12056 -5165
rect 12022 -5271 12056 -5235
rect 12280 -5131 12314 -5095
rect 12280 -5201 12314 -5165
rect 12280 -5271 12314 -5235
rect 12538 -5131 12572 -5095
rect 12538 -5201 12572 -5165
rect 12538 -5271 12572 -5235
rect 5141 -5550 5175 -5514
rect 5141 -5620 5175 -5584
rect 5141 -5690 5175 -5654
rect 5399 -5550 5433 -5514
rect 5399 -5620 5433 -5584
rect 5399 -5690 5433 -5654
rect 5657 -5550 5691 -5514
rect 5657 -5620 5691 -5584
rect 5657 -5691 5691 -5655
rect 5915 -5550 5949 -5514
rect 5915 -5620 5949 -5584
rect 5915 -5690 5949 -5654
rect 6173 -5550 6207 -5514
rect 6173 -5620 6207 -5584
rect 6173 -5690 6207 -5654
rect 6431 -5550 6465 -5514
rect 6431 -5620 6465 -5584
rect 6431 -5690 6465 -5654
rect 6689 -5550 6723 -5514
rect 6689 -5620 6723 -5584
rect 6689 -5690 6723 -5654
rect 6947 -5550 6981 -5514
rect 6947 -5620 6981 -5584
rect 6947 -5690 6981 -5654
rect 7205 -5550 7239 -5514
rect 7205 -5620 7239 -5584
rect 7205 -5690 7239 -5654
rect 7811 -5550 7845 -5514
rect 7811 -5620 7845 -5584
rect 7811 -5690 7845 -5654
rect 8069 -5550 8103 -5514
rect 8069 -5620 8103 -5584
rect 8069 -5690 8103 -5654
rect 8327 -5550 8361 -5514
rect 8327 -5620 8361 -5584
rect 8327 -5691 8361 -5655
rect 8585 -5550 8619 -5514
rect 8585 -5620 8619 -5584
rect 8585 -5690 8619 -5654
rect 8843 -5550 8877 -5514
rect 8843 -5620 8877 -5584
rect 8843 -5690 8877 -5654
rect 9101 -5550 9135 -5514
rect 9101 -5620 9135 -5584
rect 9101 -5690 9135 -5654
rect 9359 -5550 9393 -5514
rect 9359 -5620 9393 -5584
rect 9359 -5690 9393 -5654
rect 9617 -5550 9651 -5514
rect 9617 -5620 9651 -5584
rect 9617 -5690 9651 -5654
rect 9875 -5550 9909 -5514
rect 9875 -5620 9909 -5584
rect 9875 -5690 9909 -5654
rect 10474 -5549 10508 -5513
rect 10474 -5619 10508 -5583
rect 10474 -5689 10508 -5653
rect 10732 -5549 10766 -5513
rect 10732 -5619 10766 -5583
rect 10732 -5689 10766 -5653
rect 10990 -5549 11024 -5513
rect 10990 -5619 11024 -5583
rect 10990 -5690 11024 -5654
rect 11248 -5549 11282 -5513
rect 11248 -5619 11282 -5583
rect 11248 -5689 11282 -5653
rect 11506 -5549 11540 -5513
rect 11506 -5619 11540 -5583
rect 11506 -5689 11540 -5653
rect 11764 -5549 11798 -5513
rect 11764 -5619 11798 -5583
rect 11764 -5689 11798 -5653
rect 12022 -5549 12056 -5513
rect 12022 -5619 12056 -5583
rect 12022 -5689 12056 -5653
rect 12280 -5549 12314 -5513
rect 12280 -5619 12314 -5583
rect 12280 -5689 12314 -5653
rect 12538 -5549 12572 -5513
rect 12538 -5619 12572 -5583
rect 12538 -5689 12572 -5653
rect 5141 -5968 5175 -5932
rect 5141 -6038 5175 -6002
rect 5141 -6108 5175 -6072
rect 5399 -5968 5433 -5932
rect 5399 -6038 5433 -6002
rect 5399 -6108 5433 -6072
rect 5657 -5968 5691 -5932
rect 5657 -6038 5691 -6002
rect 5657 -6109 5691 -6073
rect 5915 -5968 5949 -5932
rect 5915 -6038 5949 -6002
rect 5915 -6108 5949 -6072
rect 6173 -5968 6207 -5932
rect 6173 -6038 6207 -6002
rect 6173 -6108 6207 -6072
rect 6431 -5968 6465 -5932
rect 6431 -6038 6465 -6002
rect 6431 -6108 6465 -6072
rect 6689 -5968 6723 -5932
rect 6689 -6038 6723 -6002
rect 6689 -6108 6723 -6072
rect 6947 -5968 6981 -5932
rect 6947 -6038 6981 -6002
rect 6947 -6108 6981 -6072
rect 7205 -5968 7239 -5932
rect 7205 -6038 7239 -6002
rect 7205 -6108 7239 -6072
rect 7811 -5968 7845 -5932
rect 7811 -6038 7845 -6002
rect 7811 -6108 7845 -6072
rect 8069 -5968 8103 -5932
rect 8069 -6038 8103 -6002
rect 8069 -6108 8103 -6072
rect 8327 -5968 8361 -5932
rect 8327 -6038 8361 -6002
rect 8327 -6109 8361 -6073
rect 8585 -5968 8619 -5932
rect 8585 -6038 8619 -6002
rect 8585 -6108 8619 -6072
rect 8843 -5968 8877 -5932
rect 8843 -6038 8877 -6002
rect 8843 -6108 8877 -6072
rect 9101 -5968 9135 -5932
rect 9101 -6038 9135 -6002
rect 9101 -6108 9135 -6072
rect 9359 -5968 9393 -5932
rect 9359 -6038 9393 -6002
rect 9359 -6108 9393 -6072
rect 9617 -5968 9651 -5932
rect 9617 -6038 9651 -6002
rect 9617 -6108 9651 -6072
rect 9875 -5968 9909 -5932
rect 9875 -6038 9909 -6002
rect 9875 -6108 9909 -6072
rect 10474 -5967 10508 -5931
rect 10474 -6037 10508 -6001
rect 10474 -6107 10508 -6071
rect 10732 -5967 10766 -5931
rect 10732 -6037 10766 -6001
rect 10732 -6107 10766 -6071
rect 10990 -5967 11024 -5931
rect 10990 -6037 11024 -6001
rect 10990 -6108 11024 -6072
rect 11248 -5967 11282 -5931
rect 11248 -6037 11282 -6001
rect 11248 -6107 11282 -6071
rect 11506 -5967 11540 -5931
rect 11506 -6037 11540 -6001
rect 11506 -6107 11540 -6071
rect 11764 -5967 11798 -5931
rect 11764 -6037 11798 -6001
rect 11764 -6107 11798 -6071
rect 12022 -5967 12056 -5931
rect 12022 -6037 12056 -6001
rect 12022 -6107 12056 -6071
rect 12280 -5967 12314 -5931
rect 12280 -6037 12314 -6001
rect 12280 -6107 12314 -6071
rect 12538 -5967 12572 -5931
rect 12538 -6037 12572 -6001
rect 12538 -6107 12572 -6071
rect 5141 -6386 5175 -6350
rect 5141 -6456 5175 -6420
rect 5141 -6526 5175 -6490
rect 5399 -6386 5433 -6350
rect 5399 -6456 5433 -6420
rect 5399 -6526 5433 -6490
rect 5657 -6386 5691 -6350
rect 5657 -6456 5691 -6420
rect 5657 -6527 5691 -6491
rect 5915 -6386 5949 -6350
rect 5915 -6456 5949 -6420
rect 5915 -6526 5949 -6490
rect 6173 -6386 6207 -6350
rect 6173 -6456 6207 -6420
rect 6173 -6526 6207 -6490
rect 6431 -6386 6465 -6350
rect 6431 -6456 6465 -6420
rect 6431 -6526 6465 -6490
rect 6689 -6386 6723 -6350
rect 6689 -6456 6723 -6420
rect 6689 -6526 6723 -6490
rect 6947 -6386 6981 -6350
rect 6947 -6456 6981 -6420
rect 6947 -6526 6981 -6490
rect 7205 -6386 7239 -6350
rect 7205 -6456 7239 -6420
rect 7205 -6526 7239 -6490
rect 7811 -6386 7845 -6350
rect 7811 -6456 7845 -6420
rect 7811 -6526 7845 -6490
rect 8069 -6386 8103 -6350
rect 8069 -6456 8103 -6420
rect 8069 -6526 8103 -6490
rect 8327 -6386 8361 -6350
rect 8327 -6456 8361 -6420
rect 8327 -6527 8361 -6491
rect 8585 -6386 8619 -6350
rect 8585 -6456 8619 -6420
rect 8585 -6526 8619 -6490
rect 8843 -6386 8877 -6350
rect 8843 -6456 8877 -6420
rect 8843 -6526 8877 -6490
rect 9101 -6386 9135 -6350
rect 9101 -6456 9135 -6420
rect 9101 -6526 9135 -6490
rect 9359 -6386 9393 -6350
rect 9359 -6456 9393 -6420
rect 9359 -6526 9393 -6490
rect 9617 -6386 9651 -6350
rect 9617 -6456 9651 -6420
rect 9617 -6526 9651 -6490
rect 9875 -6386 9909 -6350
rect 9875 -6456 9909 -6420
rect 9875 -6526 9909 -6490
rect 10474 -6385 10508 -6349
rect 10474 -6455 10508 -6419
rect 10474 -6525 10508 -6489
rect 10732 -6385 10766 -6349
rect 10732 -6455 10766 -6419
rect 10732 -6525 10766 -6489
rect 10990 -6385 11024 -6349
rect 10990 -6455 11024 -6419
rect 10990 -6526 11024 -6490
rect 11248 -6385 11282 -6349
rect 11248 -6455 11282 -6419
rect 11248 -6525 11282 -6489
rect 11506 -6385 11540 -6349
rect 11506 -6455 11540 -6419
rect 11506 -6525 11540 -6489
rect 11764 -6385 11798 -6349
rect 11764 -6455 11798 -6419
rect 11764 -6525 11798 -6489
rect 12022 -6385 12056 -6349
rect 12022 -6455 12056 -6419
rect 12022 -6525 12056 -6489
rect 12280 -6385 12314 -6349
rect 12280 -6455 12314 -6419
rect 12280 -6525 12314 -6489
rect 12538 -6385 12572 -6349
rect 12538 -6455 12572 -6419
rect 12538 -6525 12572 -6489
rect 5141 -6804 5175 -6768
rect 5141 -6874 5175 -6838
rect 5141 -6944 5175 -6908
rect 5399 -6804 5433 -6768
rect 5399 -6874 5433 -6838
rect 5399 -6944 5433 -6908
rect 5657 -6804 5691 -6768
rect 5657 -6874 5691 -6838
rect 5657 -6945 5691 -6909
rect 5915 -6804 5949 -6768
rect 5915 -6874 5949 -6838
rect 5915 -6944 5949 -6908
rect 6173 -6804 6207 -6768
rect 6173 -6874 6207 -6838
rect 6173 -6944 6207 -6908
rect 6431 -6804 6465 -6768
rect 6431 -6874 6465 -6838
rect 6431 -6944 6465 -6908
rect 6689 -6804 6723 -6768
rect 6689 -6874 6723 -6838
rect 6689 -6944 6723 -6908
rect 6947 -6804 6981 -6768
rect 6947 -6874 6981 -6838
rect 6947 -6944 6981 -6908
rect 7205 -6804 7239 -6768
rect 7205 -6874 7239 -6838
rect 7205 -6944 7239 -6908
rect 7811 -6804 7845 -6768
rect 7811 -6874 7845 -6838
rect 7811 -6944 7845 -6908
rect 8069 -6804 8103 -6768
rect 8069 -6874 8103 -6838
rect 8069 -6944 8103 -6908
rect 8327 -6804 8361 -6768
rect 8327 -6874 8361 -6838
rect 8327 -6945 8361 -6909
rect 8585 -6804 8619 -6768
rect 8585 -6874 8619 -6838
rect 8585 -6944 8619 -6908
rect 8843 -6804 8877 -6768
rect 8843 -6874 8877 -6838
rect 8843 -6944 8877 -6908
rect 9101 -6804 9135 -6768
rect 9101 -6874 9135 -6838
rect 9101 -6944 9135 -6908
rect 9359 -6804 9393 -6768
rect 9359 -6874 9393 -6838
rect 9359 -6944 9393 -6908
rect 9617 -6804 9651 -6768
rect 9617 -6874 9651 -6838
rect 9617 -6944 9651 -6908
rect 9875 -6804 9909 -6768
rect 9875 -6874 9909 -6838
rect 9875 -6944 9909 -6908
rect 10474 -6803 10508 -6767
rect 10474 -6873 10508 -6837
rect 10474 -6943 10508 -6907
rect 10732 -6803 10766 -6767
rect 10732 -6873 10766 -6837
rect 10732 -6943 10766 -6907
rect 10990 -6803 11024 -6767
rect 10990 -6873 11024 -6837
rect 10990 -6944 11024 -6908
rect 11248 -6803 11282 -6767
rect 11248 -6873 11282 -6837
rect 11248 -6943 11282 -6907
rect 11506 -6803 11540 -6767
rect 11506 -6873 11540 -6837
rect 11506 -6943 11540 -6907
rect 11764 -6803 11798 -6767
rect 11764 -6873 11798 -6837
rect 11764 -6943 11798 -6907
rect 12022 -6803 12056 -6767
rect 12022 -6873 12056 -6837
rect 12022 -6943 12056 -6907
rect 12280 -6803 12314 -6767
rect 12280 -6873 12314 -6837
rect 12280 -6943 12314 -6907
rect 12538 -6803 12572 -6767
rect 12538 -6873 12572 -6837
rect 12538 -6943 12572 -6907
rect 5141 -7222 5175 -7186
rect 5141 -7292 5175 -7256
rect 5141 -7362 5175 -7326
rect 5399 -7222 5433 -7186
rect 5399 -7292 5433 -7256
rect 5399 -7362 5433 -7326
rect 5657 -7222 5691 -7186
rect 5657 -7292 5691 -7256
rect 5657 -7363 5691 -7327
rect 5915 -7222 5949 -7186
rect 5915 -7292 5949 -7256
rect 5915 -7362 5949 -7326
rect 6173 -7222 6207 -7186
rect 6173 -7292 6207 -7256
rect 6173 -7362 6207 -7326
rect 6431 -7222 6465 -7186
rect 6431 -7292 6465 -7256
rect 6431 -7362 6465 -7326
rect 6689 -7222 6723 -7186
rect 6689 -7292 6723 -7256
rect 6689 -7362 6723 -7326
rect 6947 -7222 6981 -7186
rect 6947 -7292 6981 -7256
rect 6947 -7362 6981 -7326
rect 7205 -7222 7239 -7186
rect 7205 -7292 7239 -7256
rect 7205 -7362 7239 -7326
rect 7811 -7222 7845 -7186
rect 7811 -7292 7845 -7256
rect 7811 -7362 7845 -7326
rect 8069 -7222 8103 -7186
rect 8069 -7292 8103 -7256
rect 8069 -7362 8103 -7326
rect 8327 -7222 8361 -7186
rect 8327 -7292 8361 -7256
rect 8327 -7363 8361 -7327
rect 8585 -7222 8619 -7186
rect 8585 -7292 8619 -7256
rect 8585 -7362 8619 -7326
rect 8843 -7222 8877 -7186
rect 8843 -7292 8877 -7256
rect 8843 -7362 8877 -7326
rect 9101 -7222 9135 -7186
rect 9101 -7292 9135 -7256
rect 9101 -7362 9135 -7326
rect 9359 -7222 9393 -7186
rect 9359 -7292 9393 -7256
rect 9359 -7362 9393 -7326
rect 9617 -7222 9651 -7186
rect 9617 -7292 9651 -7256
rect 9617 -7362 9651 -7326
rect 9875 -7222 9909 -7186
rect 9875 -7292 9909 -7256
rect 9875 -7362 9909 -7326
rect 10474 -7221 10508 -7185
rect 10474 -7291 10508 -7255
rect 10474 -7361 10508 -7325
rect 10732 -7221 10766 -7185
rect 10732 -7291 10766 -7255
rect 10732 -7361 10766 -7325
rect 10990 -7221 11024 -7185
rect 10990 -7291 11024 -7255
rect 10990 -7362 11024 -7326
rect 11248 -7221 11282 -7185
rect 11248 -7291 11282 -7255
rect 11248 -7361 11282 -7325
rect 11506 -7221 11540 -7185
rect 11506 -7291 11540 -7255
rect 11506 -7361 11540 -7325
rect 11764 -7221 11798 -7185
rect 11764 -7291 11798 -7255
rect 11764 -7361 11798 -7325
rect 12022 -7221 12056 -7185
rect 12022 -7291 12056 -7255
rect 12022 -7361 12056 -7325
rect 12280 -7221 12314 -7185
rect 12280 -7291 12314 -7255
rect 12280 -7361 12314 -7325
rect 12538 -7221 12572 -7185
rect 12538 -7291 12572 -7255
rect 12538 -7361 12572 -7325
rect 5141 -7640 5175 -7604
rect 5141 -7710 5175 -7674
rect 5141 -7780 5175 -7744
rect 5399 -7640 5433 -7604
rect 5399 -7710 5433 -7674
rect 5399 -7780 5433 -7744
rect 5657 -7640 5691 -7604
rect 5657 -7710 5691 -7674
rect 5657 -7781 5691 -7745
rect 5915 -7640 5949 -7604
rect 5915 -7710 5949 -7674
rect 5915 -7780 5949 -7744
rect 6173 -7640 6207 -7604
rect 6173 -7710 6207 -7674
rect 6173 -7780 6207 -7744
rect 6431 -7640 6465 -7604
rect 6431 -7710 6465 -7674
rect 6431 -7780 6465 -7744
rect 6689 -7640 6723 -7604
rect 6689 -7710 6723 -7674
rect 6689 -7780 6723 -7744
rect 6947 -7640 6981 -7604
rect 6947 -7710 6981 -7674
rect 6947 -7780 6981 -7744
rect 7205 -7640 7239 -7604
rect 7205 -7710 7239 -7674
rect 7205 -7780 7239 -7744
rect 7811 -7640 7845 -7604
rect 7811 -7710 7845 -7674
rect 7811 -7780 7845 -7744
rect 8069 -7640 8103 -7604
rect 8069 -7710 8103 -7674
rect 8069 -7780 8103 -7744
rect 8327 -7640 8361 -7604
rect 8327 -7710 8361 -7674
rect 8327 -7781 8361 -7745
rect 8585 -7640 8619 -7604
rect 8585 -7710 8619 -7674
rect 8585 -7780 8619 -7744
rect 8843 -7640 8877 -7604
rect 8843 -7710 8877 -7674
rect 8843 -7780 8877 -7744
rect 9101 -7640 9135 -7604
rect 9101 -7710 9135 -7674
rect 9101 -7780 9135 -7744
rect 9359 -7640 9393 -7604
rect 9359 -7710 9393 -7674
rect 9359 -7780 9393 -7744
rect 9617 -7640 9651 -7604
rect 9617 -7710 9651 -7674
rect 9617 -7780 9651 -7744
rect 9875 -7640 9909 -7604
rect 9875 -7710 9909 -7674
rect 9875 -7780 9909 -7744
rect 10474 -7639 10508 -7603
rect 10474 -7709 10508 -7673
rect 10474 -7779 10508 -7743
rect 10732 -7639 10766 -7603
rect 10732 -7709 10766 -7673
rect 10732 -7779 10766 -7743
rect 10990 -7639 11024 -7603
rect 10990 -7709 11024 -7673
rect 10990 -7780 11024 -7744
rect 11248 -7639 11282 -7603
rect 11248 -7709 11282 -7673
rect 11248 -7779 11282 -7743
rect 11506 -7639 11540 -7603
rect 11506 -7709 11540 -7673
rect 11506 -7779 11540 -7743
rect 11764 -7639 11798 -7603
rect 11764 -7709 11798 -7673
rect 11764 -7779 11798 -7743
rect 12022 -7639 12056 -7603
rect 12022 -7709 12056 -7673
rect 12022 -7779 12056 -7743
rect 12280 -7639 12314 -7603
rect 12280 -7709 12314 -7673
rect 12280 -7779 12314 -7743
rect 12538 -7639 12572 -7603
rect 12538 -7709 12572 -7673
rect 12538 -7779 12572 -7743
rect 5021 -8292 5055 -8258
rect 5021 -8362 5055 -8326
rect 5021 -8430 5055 -8396
rect 5279 -8292 5313 -8258
rect 5279 -8362 5313 -8326
rect 5279 -8430 5313 -8396
rect 5561 -8292 5595 -8258
rect 5561 -8362 5595 -8326
rect 5561 -8430 5595 -8396
rect 5819 -8292 5853 -8258
rect 5819 -8362 5853 -8326
rect 5819 -8430 5853 -8396
rect 6041 -8292 6075 -8258
rect 6041 -8362 6075 -8326
rect 6041 -8430 6075 -8396
rect 6299 -8292 6333 -8258
rect 6299 -8362 6333 -8326
rect 6299 -8430 6333 -8396
rect 6544 -8290 6578 -8256
rect 6544 -8360 6578 -8324
rect 6544 -8428 6578 -8394
rect 6802 -8290 6836 -8256
rect 6802 -8360 6836 -8324
rect 6802 -8428 6836 -8394
rect 7054 -8280 7088 -8246
rect 7054 -8350 7088 -8314
rect 7054 -8418 7088 -8384
rect 7312 -8280 7346 -8246
rect 7312 -8350 7346 -8314
rect 7312 -8418 7346 -8384
rect 7691 -8292 7725 -8258
rect 7691 -8362 7725 -8326
rect 7691 -8430 7725 -8396
rect 7949 -8292 7983 -8258
rect 7949 -8362 7983 -8326
rect 7949 -8430 7983 -8396
rect 8231 -8292 8265 -8258
rect 8231 -8362 8265 -8326
rect 8231 -8430 8265 -8396
rect 8489 -8292 8523 -8258
rect 8489 -8362 8523 -8326
rect 8489 -8430 8523 -8396
rect 8711 -8292 8745 -8258
rect 8711 -8362 8745 -8326
rect 8711 -8430 8745 -8396
rect 8969 -8292 9003 -8258
rect 8969 -8362 9003 -8326
rect 8969 -8430 9003 -8396
rect 9214 -8290 9248 -8256
rect 9214 -8360 9248 -8324
rect 9214 -8428 9248 -8394
rect 9472 -8290 9506 -8256
rect 9472 -8360 9506 -8324
rect 9472 -8428 9506 -8394
rect 9724 -8280 9758 -8246
rect 9724 -8350 9758 -8314
rect 9724 -8418 9758 -8384
rect 9982 -8280 10016 -8246
rect 9982 -8350 10016 -8314
rect 9982 -8418 10016 -8384
rect 10354 -8291 10388 -8257
rect 10354 -8361 10388 -8325
rect 10354 -8429 10388 -8395
rect 10612 -8291 10646 -8257
rect 10612 -8361 10646 -8325
rect 10612 -8429 10646 -8395
rect 10894 -8291 10928 -8257
rect 10894 -8361 10928 -8325
rect 10894 -8429 10928 -8395
rect 11152 -8291 11186 -8257
rect 11152 -8361 11186 -8325
rect 11152 -8429 11186 -8395
rect 11374 -8291 11408 -8257
rect 11374 -8361 11408 -8325
rect 11374 -8429 11408 -8395
rect 11632 -8291 11666 -8257
rect 11632 -8361 11666 -8325
rect 11632 -8429 11666 -8395
rect 11877 -8289 11911 -8255
rect 11877 -8359 11911 -8323
rect 11877 -8427 11911 -8393
rect 12135 -8289 12169 -8255
rect 12135 -8359 12169 -8323
rect 12135 -8427 12169 -8393
rect 12387 -8279 12421 -8245
rect 12387 -8349 12421 -8313
rect 12387 -8417 12421 -8383
rect 12645 -8279 12679 -8245
rect 12645 -8349 12679 -8313
rect 12645 -8417 12679 -8383
rect 14018 7163 14052 8539
rect 15676 7163 15710 8539
rect 17334 7163 17368 8539
rect 14018 5653 14052 7029
rect 15676 5653 15710 7029
rect 17334 5653 17368 7029
rect 14018 4143 14052 5519
rect 15676 4143 15710 5519
rect 17334 4143 17368 5519
rect 14018 2633 14052 4009
rect 15676 2633 15710 4009
rect 17334 2633 17368 4009
rect 14018 1123 14052 2499
rect 15676 1123 15710 2499
rect 17334 1123 17368 2499
rect 14018 -387 14052 989
rect 15676 -387 15710 989
rect 17334 -387 17368 989
rect 14018 -1897 14052 -521
rect 15676 -1897 15710 -521
rect 17334 -1897 17368 -521
rect 14018 -3407 14052 -2031
rect 15676 -3407 15710 -2031
rect 17334 -3407 17368 -2031
rect 14018 -4917 14052 -3541
rect 15676 -4917 15710 -3541
rect 17334 -4917 17368 -3541
rect 14018 -6427 14052 -5051
rect 15676 -6427 15710 -5051
rect 17334 -6427 17368 -5051
rect 14018 -7937 14052 -6561
rect 15676 -7937 15710 -6561
rect 17334 -7937 17368 -6561
rect 14018 -9447 14052 -8071
rect 15676 -9447 15710 -8071
rect 17334 -9447 17368 -8071
<< pdiffc >>
rect 5416 8454 5450 8490
rect 5415 8380 5449 8416
rect 5415 8307 5449 8343
rect 5673 8450 5707 8486
rect 5673 8380 5707 8416
rect 5672 8307 5706 8343
rect 6076 8454 6110 8490
rect 6075 8380 6109 8416
rect 6075 8307 6109 8343
rect 6333 8450 6367 8486
rect 6333 8380 6367 8416
rect 6332 8307 6366 8343
rect 6546 8454 6580 8490
rect 6545 8380 6579 8416
rect 6545 8307 6579 8343
rect 6803 8450 6837 8486
rect 6803 8380 6837 8416
rect 6802 8307 6836 8343
rect 7148 8450 7182 8486
rect 7148 8379 7182 8415
rect 7148 8308 7182 8344
rect 7406 8450 7440 8486
rect 7406 8379 7440 8415
rect 7406 8308 7440 8344
rect 7664 8450 7698 8486
rect 7664 8379 7698 8415
rect 7664 8308 7698 8344
rect 7922 8450 7956 8486
rect 7922 8379 7956 8415
rect 7922 8308 7956 8344
rect 8180 8450 8214 8486
rect 8180 8379 8214 8415
rect 8180 8308 8214 8344
rect 8438 8450 8472 8486
rect 8438 8379 8472 8415
rect 8438 8308 8472 8344
rect 8963 8450 8997 8486
rect 8963 8379 8997 8415
rect 8963 8308 8997 8344
rect 9221 8450 9255 8486
rect 9221 8379 9255 8415
rect 9221 8308 9255 8344
rect 9479 8450 9513 8486
rect 9479 8379 9513 8415
rect 9479 8308 9513 8344
rect 9737 8450 9771 8486
rect 9737 8379 9771 8415
rect 9737 8308 9771 8344
rect 9995 8450 10029 8486
rect 9995 8379 10029 8415
rect 9995 8308 10029 8344
rect 10253 8450 10287 8486
rect 10253 8379 10287 8415
rect 10253 8308 10287 8344
rect 10769 8450 10803 8486
rect 10769 8379 10803 8415
rect 10769 8308 10803 8344
rect 11027 8450 11061 8486
rect 11027 8379 11061 8415
rect 11027 8308 11061 8344
rect 11285 8450 11319 8486
rect 11285 8379 11319 8415
rect 11285 8308 11319 8344
rect 11543 8450 11577 8486
rect 11543 8379 11577 8415
rect 11543 8308 11577 8344
rect 11801 8450 11835 8486
rect 11801 8379 11835 8415
rect 11801 8308 11835 8344
rect 12059 8450 12093 8486
rect 12059 8379 12093 8415
rect 12059 8308 12093 8344
rect 5358 7450 5396 7486
rect 5544 7452 5582 7488
rect 5719 7452 5753 7486
rect 6577 7452 6611 7486
rect 6744 7450 6782 7486
rect 6930 7452 6968 7488
rect 7114 7450 7152 7486
rect 7300 7452 7338 7488
rect 7536 7450 7574 7486
rect 7722 7452 7760 7488
rect 7958 7450 7996 7486
rect 8144 7452 8182 7488
rect 8389 7452 8423 7486
rect 9247 7452 9281 7486
rect 9458 7450 9496 7486
rect 9644 7452 9682 7488
rect 9828 7450 9866 7486
rect 10014 7452 10052 7488
rect 10250 7450 10288 7486
rect 10436 7452 10474 7488
rect 10672 7450 10710 7486
rect 10858 7452 10896 7488
rect 11052 7453 11086 7487
rect 11910 7453 11944 7487
rect 12112 7450 12150 7486
rect 12298 7452 12336 7488
rect 5358 1768 5396 1804
rect 5544 1770 5582 1806
rect 5711 1770 5745 1804
rect 6569 1770 6603 1804
rect 6744 1767 6782 1803
rect 6930 1769 6968 1805
rect 7114 1767 7152 1803
rect 7300 1769 7338 1805
rect 7536 1767 7574 1803
rect 7722 1769 7760 1805
rect 7958 1767 7996 1803
rect 8144 1769 8182 1805
rect 8388 1770 8422 1804
rect 9246 1770 9280 1804
rect 9458 1771 9496 1807
rect 9644 1773 9682 1809
rect 9828 1771 9866 1807
rect 10014 1773 10052 1809
rect 10250 1771 10288 1807
rect 10436 1773 10474 1809
rect 10672 1771 10710 1807
rect 10858 1773 10896 1809
rect 11052 1771 11086 1805
rect 11910 1771 11944 1805
rect 12056 1768 12094 1804
rect 12242 1770 12280 1806
rect 5403 -4156 5441 -4120
rect 5589 -4154 5627 -4118
rect 5719 -4155 5753 -4121
rect 6577 -4155 6611 -4121
rect 6744 -4158 6782 -4122
rect 6930 -4156 6968 -4120
rect 7114 -4158 7152 -4122
rect 7300 -4156 7338 -4120
rect 7536 -4158 7574 -4122
rect 7722 -4156 7760 -4120
rect 7958 -4158 7996 -4122
rect 8144 -4156 8182 -4120
rect 8389 -4155 8423 -4121
rect 9247 -4155 9281 -4121
rect 9445 -4158 9483 -4122
rect 9631 -4156 9669 -4120
rect 9815 -4158 9853 -4122
rect 10001 -4156 10039 -4120
rect 10237 -4158 10275 -4122
rect 10423 -4156 10461 -4120
rect 10659 -4158 10697 -4122
rect 10845 -4156 10883 -4120
rect 11052 -4154 11086 -4120
rect 11910 -4154 11944 -4120
rect 12682 -3773 12716 -3461
rect 12770 -3773 12804 -3461
rect 13072 -3775 13106 -3463
rect 13160 -3775 13194 -3463
<< psubdiff >>
rect 283 8628 317 8653
rect 3827 8628 3861 8653
rect 283 -9600 317 -9538
rect 13904 8629 13938 8654
rect 4744 6666 12908 6796
rect 4744 3024 4954 6666
rect 12756 3024 12906 6666
rect 4744 3012 12906 3024
rect 4744 2906 5998 3012
rect 6104 2906 8662 3012
rect 8768 2906 11324 3012
rect 11430 2906 12906 3012
rect 4744 2870 12906 2906
rect 4744 2866 4954 2870
rect 4698 1138 12958 1144
rect 4698 956 12964 1138
rect 4698 -2692 4890 956
rect 12786 -2692 12964 956
rect 4698 -2712 12964 -2692
rect 4698 -2806 6000 -2712
rect 6092 -2806 8668 -2712
rect 8760 -2806 11334 -2712
rect 11426 -2806 12964 -2712
rect 4698 -2840 12964 -2806
rect 12548 -4096 13340 -4062
rect 12548 -4242 12606 -4096
rect 12548 -4314 12554 -4242
rect 12598 -4314 12606 -4242
rect 12548 -4460 12606 -4314
rect 12874 -4242 12996 -4096
rect 12874 -4314 12944 -4242
rect 12988 -4314 12996 -4242
rect 12874 -4460 12996 -4314
rect 13264 -4460 13340 -4096
rect 12548 -4494 13340 -4460
rect 4542 -4742 13080 -4740
rect 4542 -4940 13082 -4742
rect 4542 -8574 4846 -4940
rect 12814 -8574 13082 -4940
rect 4542 -8608 13084 -8574
rect 4542 -8702 6000 -8608
rect 6092 -8702 8670 -8608
rect 8762 -8702 11336 -8608
rect 11428 -8702 13084 -8608
rect 4542 -8868 13084 -8702
rect 3827 -9600 3861 -9538
rect 283 -9634 379 -9600
rect 3765 -9634 3861 -9600
rect 17448 8629 17482 8654
rect 13904 -9599 13938 -9537
rect 17448 -9599 17482 -9537
rect 13904 -9633 14000 -9599
rect 17386 -9633 17482 -9599
<< nsubdiff >>
rect 5034 8860 5266 8864
rect 5024 8794 12718 8860
rect 5024 8699 6194 8794
rect 6822 8790 12718 8794
rect 6822 8699 8974 8790
rect 5024 8695 8974 8699
rect 9602 8695 12718 8790
rect 5024 8680 12718 8695
rect 5034 7498 5266 8680
rect 12090 8678 12718 8680
rect 12434 8038 12718 8678
rect 5034 7236 5083 7498
rect 5220 7236 5266 7498
rect 12432 7479 12718 8038
rect 5034 7140 5266 7236
rect 12432 7217 12502 7479
rect 12639 7217 12718 7479
rect 12432 7140 12718 7217
rect 5032 6904 12718 7140
rect 5032 6900 12586 6904
rect 12090 6898 12586 6900
rect 5024 2344 12636 2348
rect 5018 2338 12636 2344
rect 5018 2196 12686 2338
rect 5018 1932 5234 2196
rect 5018 1670 5042 1932
rect 5179 1670 5234 1932
rect 5018 1464 5234 1670
rect 12386 1925 12686 2196
rect 12386 1663 12456 1925
rect 12593 1663 12686 1925
rect 12386 1464 12686 1663
rect 5018 1324 12686 1464
rect 5024 1318 12686 1324
rect 12528 -3268 12918 -3266
rect 12528 -3300 13308 -3268
rect 4717 -3364 5194 -3354
rect 4717 -3370 5338 -3364
rect 4717 -3372 12402 -3370
rect 12528 -3372 12602 -3300
rect 12872 -3302 13308 -3300
rect 4717 -3406 12602 -3372
rect 4717 -3550 12276 -3406
rect 4717 -3951 5301 -3550
rect 4717 -4212 5001 -3951
rect 5137 -4212 5301 -3951
rect 12132 -3720 12276 -3550
rect 12478 -3408 12602 -3406
rect 12478 -3576 12616 -3408
rect 12478 -3638 12538 -3576
rect 12594 -3638 12616 -3576
rect 12478 -3720 12616 -3638
rect 12132 -3722 12616 -3720
rect 12132 -3760 12602 -3722
rect 4717 -4392 5301 -4212
rect 12132 -4392 12402 -3760
rect 12528 -3930 12602 -3760
rect 12872 -3578 12992 -3302
rect 12872 -3640 12928 -3578
rect 12984 -3640 12992 -3578
rect 12872 -3930 12992 -3640
rect 13262 -3930 13308 -3302
rect 12528 -3960 13308 -3930
rect 12528 -3968 12828 -3960
rect 12528 -3970 12600 -3968
rect 12996 -3970 13308 -3960
rect 4717 -4571 12402 -4392
rect 5084 -4572 12402 -4571
<< psubdiffcont >>
rect 283 -9538 317 8628
rect 3827 -9538 3861 8628
rect 5998 2906 6104 3012
rect 8662 2906 8768 3012
rect 11324 2906 11430 3012
rect 6000 -2806 6092 -2712
rect 8668 -2806 8760 -2712
rect 11334 -2806 11426 -2712
rect 12554 -4314 12598 -4242
rect 12944 -4314 12988 -4242
rect 6000 -8702 6092 -8608
rect 8670 -8702 8762 -8608
rect 11336 -8702 11428 -8608
rect 379 -9634 3765 -9600
rect 13904 -9537 13938 8629
rect 17448 -9537 17482 8629
rect 14000 -9633 17386 -9599
<< nsubdiffcont >>
rect 6194 8699 6822 8794
rect 8974 8695 9602 8790
rect 5083 7236 5220 7498
rect 12502 7217 12639 7479
rect 5042 1670 5179 1932
rect 12456 1663 12593 1925
rect 5001 -4212 5137 -3951
rect 12276 -3720 12478 -3406
rect 12538 -3638 12594 -3576
rect 12928 -3640 12984 -3578
<< poly >>
rect 443 8622 2043 8638
rect 443 8588 459 8622
rect 1824 8588 2043 8622
rect 443 8550 2043 8588
rect 2101 8622 3701 8638
rect 2101 8588 2318 8622
rect 3685 8588 3701 8622
rect 2101 8550 3701 8588
rect 443 7112 2043 7150
rect 443 7078 459 7112
rect 1824 7078 2043 7112
rect 443 7040 2043 7078
rect 2101 7112 3701 7150
rect 2101 7078 2318 7112
rect 3685 7078 3701 7112
rect 2101 7040 3701 7078
rect 443 5602 2043 5640
rect 443 5568 459 5602
rect 1824 5568 2043 5602
rect 443 5530 2043 5568
rect 2101 5602 3701 5640
rect 2101 5568 2318 5602
rect 3685 5568 3701 5602
rect 2101 5530 3701 5568
rect 443 4092 2043 4130
rect 443 4058 459 4092
rect 1824 4058 2043 4092
rect 443 4020 2043 4058
rect 2101 4092 3701 4130
rect 2101 4058 2318 4092
rect 3685 4058 3701 4092
rect 2101 4020 3701 4058
rect 443 2582 2043 2620
rect 443 2548 459 2582
rect 1824 2548 2043 2582
rect 443 2510 2043 2548
rect 2101 2582 3701 2620
rect 2101 2548 2318 2582
rect 3685 2548 3701 2582
rect 2101 2510 3701 2548
rect 443 1072 2043 1110
rect 443 1038 459 1072
rect 1824 1038 2043 1072
rect 443 1000 2043 1038
rect 2101 1072 3701 1110
rect 2101 1038 2318 1072
rect 3685 1038 3701 1072
rect 2101 1000 3701 1038
rect 443 -438 2043 -400
rect 443 -472 459 -438
rect 1824 -472 2043 -438
rect 443 -510 2043 -472
rect 2101 -438 3701 -400
rect 2101 -472 2318 -438
rect 3685 -472 3701 -438
rect 2101 -510 3701 -472
rect 443 -1948 2043 -1910
rect 443 -1982 459 -1948
rect 1824 -1982 2043 -1948
rect 443 -2020 2043 -1982
rect 2101 -1948 3701 -1910
rect 2101 -1982 2318 -1948
rect 3685 -1982 3701 -1948
rect 2101 -2020 3701 -1982
rect 443 -3458 2043 -3420
rect 443 -3492 459 -3458
rect 1824 -3492 2043 -3458
rect 443 -3530 2043 -3492
rect 2101 -3458 3701 -3420
rect 2101 -3492 2318 -3458
rect 3685 -3492 3701 -3458
rect 2101 -3530 3701 -3492
rect 443 -4968 2043 -4930
rect 443 -5002 459 -4968
rect 1824 -5002 2043 -4968
rect 443 -5040 2043 -5002
rect 2101 -4968 3701 -4930
rect 2101 -5002 2318 -4968
rect 3685 -5002 3701 -4968
rect 2101 -5040 3701 -5002
rect 443 -6478 2043 -6440
rect 443 -6512 459 -6478
rect 1824 -6512 2043 -6478
rect 443 -6550 2043 -6512
rect 2101 -6478 3701 -6440
rect 2101 -6512 2318 -6478
rect 3685 -6512 3701 -6478
rect 2101 -6550 3701 -6512
rect 443 -7988 2043 -7950
rect 443 -8022 459 -7988
rect 1824 -8022 2043 -7988
rect 443 -8060 2043 -8022
rect 2101 -7988 3701 -7950
rect 2101 -8022 2318 -7988
rect 3685 -8022 3701 -7988
rect 2101 -8060 3701 -8022
rect 443 -9498 2043 -9460
rect 443 -9532 459 -9498
rect 1824 -9532 2043 -9498
rect 443 -9548 2043 -9532
rect 2101 -9498 3701 -9460
rect 2101 -9532 2318 -9498
rect 3685 -9532 3701 -9498
rect 2101 -9548 3701 -9532
rect 5528 8579 5594 8595
rect 5528 8562 5544 8579
rect 5461 8545 5544 8562
rect 5578 8562 5594 8579
rect 6188 8579 6254 8595
rect 6188 8562 6204 8579
rect 5578 8545 5661 8562
rect 5461 8498 5661 8545
rect 6121 8545 6204 8562
rect 6238 8562 6254 8579
rect 6658 8579 6724 8595
rect 6658 8562 6674 8579
rect 6238 8545 6321 8562
rect 6121 8498 6321 8545
rect 6591 8545 6674 8562
rect 6708 8562 6724 8579
rect 7261 8578 7327 8594
rect 6708 8545 6791 8562
rect 7261 8561 7277 8578
rect 6591 8498 6791 8545
rect 7194 8544 7277 8561
rect 7311 8561 7327 8578
rect 7519 8578 7585 8594
rect 7519 8561 7535 8578
rect 7311 8544 7394 8561
rect 7194 8497 7394 8544
rect 7452 8544 7535 8561
rect 7569 8561 7585 8578
rect 7777 8578 7843 8594
rect 7777 8561 7793 8578
rect 7569 8544 7652 8561
rect 7452 8497 7652 8544
rect 7710 8544 7793 8561
rect 7827 8561 7843 8578
rect 8035 8578 8101 8594
rect 8035 8561 8051 8578
rect 7827 8544 7910 8561
rect 7710 8497 7910 8544
rect 7968 8544 8051 8561
rect 8085 8561 8101 8578
rect 8293 8578 8359 8594
rect 8293 8561 8309 8578
rect 8085 8544 8168 8561
rect 7968 8497 8168 8544
rect 8226 8544 8309 8561
rect 8343 8561 8359 8578
rect 9076 8578 9142 8594
rect 9076 8561 9092 8578
rect 8343 8544 8426 8561
rect 8226 8497 8426 8544
rect 9009 8544 9092 8561
rect 9126 8561 9142 8578
rect 9334 8578 9400 8594
rect 9334 8561 9350 8578
rect 9126 8544 9209 8561
rect 9009 8497 9209 8544
rect 9267 8544 9350 8561
rect 9384 8561 9400 8578
rect 9592 8578 9658 8594
rect 9592 8561 9608 8578
rect 9384 8544 9467 8561
rect 9267 8497 9467 8544
rect 9525 8544 9608 8561
rect 9642 8561 9658 8578
rect 9850 8578 9916 8594
rect 9850 8561 9866 8578
rect 9642 8544 9725 8561
rect 9525 8497 9725 8544
rect 9783 8544 9866 8561
rect 9900 8561 9916 8578
rect 10108 8578 10174 8594
rect 10108 8561 10124 8578
rect 9900 8544 9983 8561
rect 9783 8497 9983 8544
rect 10041 8544 10124 8561
rect 10158 8561 10174 8578
rect 10882 8578 10948 8594
rect 10882 8561 10898 8578
rect 10158 8544 10241 8561
rect 10041 8497 10241 8544
rect 10815 8544 10898 8561
rect 10932 8561 10948 8578
rect 11140 8578 11206 8594
rect 11140 8561 11156 8578
rect 10932 8544 11015 8561
rect 10815 8497 11015 8544
rect 11073 8544 11156 8561
rect 11190 8561 11206 8578
rect 11398 8578 11464 8594
rect 11398 8561 11414 8578
rect 11190 8544 11273 8561
rect 11073 8497 11273 8544
rect 11331 8544 11414 8561
rect 11448 8561 11464 8578
rect 11656 8578 11722 8594
rect 11656 8561 11672 8578
rect 11448 8544 11531 8561
rect 11331 8497 11531 8544
rect 11589 8544 11672 8561
rect 11706 8561 11722 8578
rect 11914 8578 11980 8594
rect 11914 8561 11930 8578
rect 11706 8544 11789 8561
rect 11589 8497 11789 8544
rect 11847 8544 11930 8561
rect 11964 8561 11980 8578
rect 11964 8544 12047 8561
rect 11847 8497 12047 8544
rect 5461 8251 5661 8298
rect 5461 8234 5544 8251
rect 5528 8217 5544 8234
rect 5578 8234 5661 8251
rect 6121 8251 6321 8298
rect 6121 8234 6204 8251
rect 5578 8217 5594 8234
rect 5528 8201 5594 8217
rect 6188 8217 6204 8234
rect 6238 8234 6321 8251
rect 6591 8251 6791 8298
rect 6591 8234 6674 8251
rect 6238 8217 6254 8234
rect 6188 8201 6254 8217
rect 6658 8217 6674 8234
rect 6708 8234 6791 8251
rect 7194 8250 7394 8297
rect 6708 8217 6724 8234
rect 7194 8233 7277 8250
rect 6658 8201 6724 8217
rect 7261 8216 7277 8233
rect 7311 8233 7394 8250
rect 7452 8250 7652 8297
rect 7452 8233 7535 8250
rect 7311 8216 7327 8233
rect 7261 8200 7327 8216
rect 7519 8216 7535 8233
rect 7569 8233 7652 8250
rect 7710 8250 7910 8297
rect 7710 8233 7793 8250
rect 7569 8216 7585 8233
rect 7519 8200 7585 8216
rect 7777 8216 7793 8233
rect 7827 8233 7910 8250
rect 7968 8250 8168 8297
rect 7968 8233 8051 8250
rect 7827 8216 7843 8233
rect 7777 8200 7843 8216
rect 8035 8216 8051 8233
rect 8085 8233 8168 8250
rect 8226 8250 8426 8297
rect 8226 8233 8309 8250
rect 8085 8216 8101 8233
rect 8035 8200 8101 8216
rect 8293 8216 8309 8233
rect 8343 8233 8426 8250
rect 9009 8250 9209 8297
rect 9009 8233 9092 8250
rect 8343 8216 8359 8233
rect 8293 8200 8359 8216
rect 9076 8216 9092 8233
rect 9126 8233 9209 8250
rect 9267 8250 9467 8297
rect 9267 8233 9350 8250
rect 9126 8216 9142 8233
rect 9076 8200 9142 8216
rect 9334 8216 9350 8233
rect 9384 8233 9467 8250
rect 9525 8250 9725 8297
rect 9525 8233 9608 8250
rect 9384 8216 9400 8233
rect 9334 8200 9400 8216
rect 9592 8216 9608 8233
rect 9642 8233 9725 8250
rect 9783 8250 9983 8297
rect 9783 8233 9866 8250
rect 9642 8216 9658 8233
rect 9592 8200 9658 8216
rect 9850 8216 9866 8233
rect 9900 8233 9983 8250
rect 10041 8250 10241 8297
rect 10041 8233 10124 8250
rect 9900 8216 9916 8233
rect 9850 8200 9916 8216
rect 10108 8216 10124 8233
rect 10158 8233 10241 8250
rect 10815 8250 11015 8297
rect 10815 8233 10898 8250
rect 10158 8216 10174 8233
rect 10108 8200 10174 8216
rect 10882 8216 10898 8233
rect 10932 8233 11015 8250
rect 11073 8250 11273 8297
rect 11073 8233 11156 8250
rect 10932 8216 10948 8233
rect 10882 8200 10948 8216
rect 11140 8216 11156 8233
rect 11190 8233 11273 8250
rect 11331 8250 11531 8297
rect 11331 8233 11414 8250
rect 11190 8216 11206 8233
rect 11140 8200 11206 8216
rect 11398 8216 11414 8233
rect 11448 8233 11531 8250
rect 11589 8250 11789 8297
rect 11589 8233 11672 8250
rect 11448 8216 11464 8233
rect 11398 8200 11464 8216
rect 11656 8216 11672 8233
rect 11706 8233 11789 8250
rect 11847 8250 12047 8297
rect 11847 8233 11930 8250
rect 11706 8216 11722 8233
rect 11656 8200 11722 8216
rect 11914 8216 11930 8233
rect 11964 8233 12047 8250
rect 11964 8216 11980 8233
rect 11914 8200 11980 8216
rect 5412 7612 5528 7640
rect 5412 7574 5436 7612
rect 5502 7574 5528 7612
rect 6072 7605 6258 7621
rect 6072 7588 6088 7605
rect 5412 7524 5528 7574
rect 5765 7571 6088 7588
rect 6242 7588 6258 7605
rect 6798 7612 6914 7640
rect 6242 7571 6565 7588
rect 5765 7524 6565 7571
rect 6798 7574 6822 7612
rect 6888 7574 6914 7612
rect 6798 7524 6914 7574
rect 7168 7612 7284 7640
rect 7168 7574 7192 7612
rect 7258 7574 7284 7612
rect 7168 7524 7284 7574
rect 7590 7612 7706 7640
rect 7590 7574 7614 7612
rect 7680 7574 7706 7612
rect 7590 7524 7706 7574
rect 8012 7612 8128 7640
rect 8012 7574 8036 7612
rect 8102 7574 8128 7612
rect 8742 7605 8928 7621
rect 8742 7588 8758 7605
rect 8012 7524 8128 7574
rect 8435 7571 8758 7588
rect 8912 7588 8928 7605
rect 9512 7612 9628 7640
rect 8912 7571 9235 7588
rect 8435 7524 9235 7571
rect 9512 7574 9536 7612
rect 9602 7574 9628 7612
rect 9512 7524 9628 7574
rect 9882 7612 9998 7640
rect 9882 7574 9906 7612
rect 9972 7574 9998 7612
rect 9882 7524 9998 7574
rect 10304 7612 10420 7640
rect 10304 7574 10328 7612
rect 10394 7574 10420 7612
rect 10304 7524 10420 7574
rect 10726 7612 10842 7640
rect 10726 7574 10750 7612
rect 10816 7574 10842 7612
rect 11405 7606 11591 7622
rect 11405 7589 11421 7606
rect 10726 7524 10842 7574
rect 11098 7572 11421 7589
rect 11575 7589 11591 7606
rect 12166 7612 12282 7640
rect 11575 7572 11898 7589
rect 11098 7525 11898 7572
rect 12166 7574 12190 7612
rect 12256 7574 12282 7612
rect 12166 7524 12282 7574
rect 5412 7350 5528 7414
rect 5765 7367 6565 7414
rect 5765 7350 6088 7367
rect 6072 7333 6088 7350
rect 6242 7350 6565 7367
rect 6798 7350 6914 7414
rect 7168 7350 7284 7414
rect 7590 7350 7706 7414
rect 8012 7350 8128 7414
rect 8435 7367 9235 7414
rect 8435 7350 8758 7367
rect 6242 7333 6258 7350
rect 6072 7317 6258 7333
rect 8742 7333 8758 7350
rect 8912 7350 9235 7367
rect 9512 7350 9628 7414
rect 9882 7350 9998 7414
rect 10304 7350 10420 7414
rect 10726 7350 10842 7414
rect 11098 7368 11898 7415
rect 11098 7351 11421 7368
rect 8912 7333 8928 7350
rect 8742 7317 8928 7333
rect 11405 7334 11421 7351
rect 11575 7351 11898 7368
rect 11575 7334 11591 7351
rect 12166 7350 12282 7414
rect 11405 7318 11591 7334
rect 5254 6609 5320 6625
rect 5254 6592 5270 6609
rect 5187 6575 5270 6592
rect 5304 6592 5320 6609
rect 5512 6609 5578 6625
rect 5512 6592 5528 6609
rect 5304 6575 5387 6592
rect 5187 6537 5387 6575
rect 5445 6575 5528 6592
rect 5562 6592 5578 6609
rect 5770 6609 5836 6625
rect 5770 6592 5786 6609
rect 5562 6575 5645 6592
rect 5445 6537 5645 6575
rect 5703 6575 5786 6592
rect 5820 6592 5836 6609
rect 6028 6609 6094 6625
rect 6028 6592 6044 6609
rect 5820 6575 5903 6592
rect 5703 6537 5903 6575
rect 5961 6575 6044 6592
rect 6078 6592 6094 6609
rect 6286 6609 6352 6625
rect 6286 6592 6302 6609
rect 6078 6575 6161 6592
rect 5961 6537 6161 6575
rect 6219 6575 6302 6592
rect 6336 6592 6352 6609
rect 6544 6609 6610 6625
rect 6544 6592 6560 6609
rect 6336 6575 6419 6592
rect 6219 6537 6419 6575
rect 6477 6575 6560 6592
rect 6594 6592 6610 6609
rect 6802 6609 6868 6625
rect 6802 6592 6818 6609
rect 6594 6575 6677 6592
rect 6477 6537 6677 6575
rect 6735 6575 6818 6592
rect 6852 6592 6868 6609
rect 7060 6609 7126 6625
rect 7060 6592 7076 6609
rect 6852 6575 6935 6592
rect 6735 6537 6935 6575
rect 6993 6575 7076 6592
rect 7110 6592 7126 6609
rect 7924 6609 7990 6625
rect 7924 6592 7940 6609
rect 7110 6575 7193 6592
rect 6993 6537 7193 6575
rect 7857 6575 7940 6592
rect 7974 6592 7990 6609
rect 8182 6609 8248 6625
rect 8182 6592 8198 6609
rect 7974 6575 8057 6592
rect 7857 6537 8057 6575
rect 8115 6575 8198 6592
rect 8232 6592 8248 6609
rect 8440 6609 8506 6625
rect 8440 6592 8456 6609
rect 8232 6575 8315 6592
rect 8115 6537 8315 6575
rect 8373 6575 8456 6592
rect 8490 6592 8506 6609
rect 8698 6609 8764 6625
rect 8698 6592 8714 6609
rect 8490 6575 8573 6592
rect 8373 6537 8573 6575
rect 8631 6575 8714 6592
rect 8748 6592 8764 6609
rect 8956 6609 9022 6625
rect 8956 6592 8972 6609
rect 8748 6575 8831 6592
rect 8631 6537 8831 6575
rect 8889 6575 8972 6592
rect 9006 6592 9022 6609
rect 9214 6609 9280 6625
rect 9214 6592 9230 6609
rect 9006 6575 9089 6592
rect 8889 6537 9089 6575
rect 9147 6575 9230 6592
rect 9264 6592 9280 6609
rect 9472 6609 9538 6625
rect 9472 6592 9488 6609
rect 9264 6575 9347 6592
rect 9147 6537 9347 6575
rect 9405 6575 9488 6592
rect 9522 6592 9538 6609
rect 9730 6609 9796 6625
rect 9730 6592 9746 6609
rect 9522 6575 9605 6592
rect 9405 6537 9605 6575
rect 9663 6575 9746 6592
rect 9780 6592 9796 6609
rect 10587 6610 10653 6626
rect 10587 6593 10603 6610
rect 9780 6575 9863 6592
rect 9663 6537 9863 6575
rect 10520 6576 10603 6593
rect 10637 6593 10653 6610
rect 10845 6610 10911 6626
rect 10845 6593 10861 6610
rect 10637 6576 10720 6593
rect 10520 6538 10720 6576
rect 10778 6576 10861 6593
rect 10895 6593 10911 6610
rect 11103 6610 11169 6626
rect 11103 6593 11119 6610
rect 10895 6576 10978 6593
rect 10778 6538 10978 6576
rect 11036 6576 11119 6593
rect 11153 6593 11169 6610
rect 11361 6610 11427 6626
rect 11361 6593 11377 6610
rect 11153 6576 11236 6593
rect 11036 6538 11236 6576
rect 11294 6576 11377 6593
rect 11411 6593 11427 6610
rect 11619 6610 11685 6626
rect 11619 6593 11635 6610
rect 11411 6576 11494 6593
rect 11294 6538 11494 6576
rect 11552 6576 11635 6593
rect 11669 6593 11685 6610
rect 11877 6610 11943 6626
rect 11877 6593 11893 6610
rect 11669 6576 11752 6593
rect 11552 6538 11752 6576
rect 11810 6576 11893 6593
rect 11927 6593 11943 6610
rect 12135 6610 12201 6626
rect 12135 6593 12151 6610
rect 11927 6576 12010 6593
rect 11810 6538 12010 6576
rect 12068 6576 12151 6593
rect 12185 6593 12201 6610
rect 12393 6610 12459 6626
rect 12393 6593 12409 6610
rect 12185 6576 12268 6593
rect 12068 6538 12268 6576
rect 12326 6576 12409 6593
rect 12443 6593 12459 6610
rect 12443 6576 12526 6593
rect 12326 6538 12526 6576
rect 5187 6299 5387 6337
rect 5187 6282 5270 6299
rect 5254 6265 5270 6282
rect 5304 6282 5387 6299
rect 5445 6299 5645 6337
rect 5445 6282 5528 6299
rect 5304 6265 5320 6282
rect 5254 6249 5320 6265
rect 5512 6265 5528 6282
rect 5562 6282 5645 6299
rect 5703 6299 5903 6337
rect 5703 6282 5786 6299
rect 5562 6265 5578 6282
rect 5512 6249 5578 6265
rect 5770 6265 5786 6282
rect 5820 6282 5903 6299
rect 5961 6299 6161 6337
rect 5961 6282 6044 6299
rect 5820 6265 5836 6282
rect 5770 6249 5836 6265
rect 6028 6265 6044 6282
rect 6078 6282 6161 6299
rect 6219 6299 6419 6337
rect 6219 6282 6302 6299
rect 6078 6265 6094 6282
rect 6028 6249 6094 6265
rect 6286 6265 6302 6282
rect 6336 6282 6419 6299
rect 6477 6299 6677 6337
rect 6477 6282 6560 6299
rect 6336 6265 6352 6282
rect 6286 6249 6352 6265
rect 6544 6265 6560 6282
rect 6594 6282 6677 6299
rect 6735 6299 6935 6337
rect 6735 6282 6818 6299
rect 6594 6265 6610 6282
rect 6544 6249 6610 6265
rect 6802 6265 6818 6282
rect 6852 6282 6935 6299
rect 6993 6299 7193 6337
rect 6993 6282 7076 6299
rect 6852 6265 6868 6282
rect 6802 6249 6868 6265
rect 7060 6265 7076 6282
rect 7110 6282 7193 6299
rect 7857 6299 8057 6337
rect 7857 6282 7940 6299
rect 7110 6265 7126 6282
rect 7060 6249 7126 6265
rect 7924 6265 7940 6282
rect 7974 6282 8057 6299
rect 8115 6299 8315 6337
rect 8115 6282 8198 6299
rect 7974 6265 7990 6282
rect 7924 6249 7990 6265
rect 8182 6265 8198 6282
rect 8232 6282 8315 6299
rect 8373 6299 8573 6337
rect 8373 6282 8456 6299
rect 8232 6265 8248 6282
rect 8182 6249 8248 6265
rect 8440 6265 8456 6282
rect 8490 6282 8573 6299
rect 8631 6299 8831 6337
rect 8631 6282 8714 6299
rect 8490 6265 8506 6282
rect 8440 6249 8506 6265
rect 8698 6265 8714 6282
rect 8748 6282 8831 6299
rect 8889 6299 9089 6337
rect 8889 6282 8972 6299
rect 8748 6265 8764 6282
rect 8698 6249 8764 6265
rect 8956 6265 8972 6282
rect 9006 6282 9089 6299
rect 9147 6299 9347 6337
rect 9147 6282 9230 6299
rect 9006 6265 9022 6282
rect 8956 6249 9022 6265
rect 9214 6265 9230 6282
rect 9264 6282 9347 6299
rect 9405 6299 9605 6337
rect 9405 6282 9488 6299
rect 9264 6265 9280 6282
rect 9214 6249 9280 6265
rect 9472 6265 9488 6282
rect 9522 6282 9605 6299
rect 9663 6299 9863 6337
rect 9663 6282 9746 6299
rect 9522 6265 9538 6282
rect 9472 6249 9538 6265
rect 9730 6265 9746 6282
rect 9780 6282 9863 6299
rect 10520 6300 10720 6338
rect 10520 6283 10603 6300
rect 9780 6265 9796 6282
rect 9730 6249 9796 6265
rect 10587 6266 10603 6283
rect 10637 6283 10720 6300
rect 10778 6300 10978 6338
rect 10778 6283 10861 6300
rect 10637 6266 10653 6283
rect 10587 6250 10653 6266
rect 10845 6266 10861 6283
rect 10895 6283 10978 6300
rect 11036 6300 11236 6338
rect 11036 6283 11119 6300
rect 10895 6266 10911 6283
rect 10845 6250 10911 6266
rect 11103 6266 11119 6283
rect 11153 6283 11236 6300
rect 11294 6300 11494 6338
rect 11294 6283 11377 6300
rect 11153 6266 11169 6283
rect 11103 6250 11169 6266
rect 11361 6266 11377 6283
rect 11411 6283 11494 6300
rect 11552 6300 11752 6338
rect 11552 6283 11635 6300
rect 11411 6266 11427 6283
rect 11361 6250 11427 6266
rect 11619 6266 11635 6283
rect 11669 6283 11752 6300
rect 11810 6300 12010 6338
rect 11810 6283 11893 6300
rect 11669 6266 11685 6283
rect 11619 6250 11685 6266
rect 11877 6266 11893 6283
rect 11927 6283 12010 6300
rect 12068 6300 12268 6338
rect 12068 6283 12151 6300
rect 11927 6266 11943 6283
rect 11877 6250 11943 6266
rect 12135 6266 12151 6283
rect 12185 6283 12268 6300
rect 12326 6300 12526 6338
rect 12326 6283 12409 6300
rect 12185 6266 12201 6283
rect 12135 6250 12201 6266
rect 12393 6266 12409 6283
rect 12443 6283 12526 6300
rect 12443 6266 12459 6283
rect 12393 6250 12459 6266
rect 5254 6191 5320 6207
rect 5254 6174 5270 6191
rect 5187 6157 5270 6174
rect 5304 6174 5320 6191
rect 5512 6191 5578 6207
rect 5512 6174 5528 6191
rect 5304 6157 5387 6174
rect 5187 6119 5387 6157
rect 5445 6157 5528 6174
rect 5562 6174 5578 6191
rect 5770 6191 5836 6207
rect 5770 6174 5786 6191
rect 5562 6157 5645 6174
rect 5445 6119 5645 6157
rect 5703 6157 5786 6174
rect 5820 6174 5836 6191
rect 6028 6191 6094 6207
rect 6028 6174 6044 6191
rect 5820 6157 5903 6174
rect 5703 6119 5903 6157
rect 5961 6157 6044 6174
rect 6078 6174 6094 6191
rect 6286 6191 6352 6207
rect 6286 6174 6302 6191
rect 6078 6157 6161 6174
rect 5961 6119 6161 6157
rect 6219 6157 6302 6174
rect 6336 6174 6352 6191
rect 6544 6191 6610 6207
rect 6544 6174 6560 6191
rect 6336 6157 6419 6174
rect 6219 6119 6419 6157
rect 6477 6157 6560 6174
rect 6594 6174 6610 6191
rect 6802 6191 6868 6207
rect 6802 6174 6818 6191
rect 6594 6157 6677 6174
rect 6477 6119 6677 6157
rect 6735 6157 6818 6174
rect 6852 6174 6868 6191
rect 7060 6191 7126 6207
rect 7060 6174 7076 6191
rect 6852 6157 6935 6174
rect 6735 6119 6935 6157
rect 6993 6157 7076 6174
rect 7110 6174 7126 6191
rect 7924 6191 7990 6207
rect 7924 6174 7940 6191
rect 7110 6157 7193 6174
rect 6993 6119 7193 6157
rect 7857 6157 7940 6174
rect 7974 6174 7990 6191
rect 8182 6191 8248 6207
rect 8182 6174 8198 6191
rect 7974 6157 8057 6174
rect 7857 6119 8057 6157
rect 8115 6157 8198 6174
rect 8232 6174 8248 6191
rect 8440 6191 8506 6207
rect 8440 6174 8456 6191
rect 8232 6157 8315 6174
rect 8115 6119 8315 6157
rect 8373 6157 8456 6174
rect 8490 6174 8506 6191
rect 8698 6191 8764 6207
rect 8698 6174 8714 6191
rect 8490 6157 8573 6174
rect 8373 6119 8573 6157
rect 8631 6157 8714 6174
rect 8748 6174 8764 6191
rect 8956 6191 9022 6207
rect 8956 6174 8972 6191
rect 8748 6157 8831 6174
rect 8631 6119 8831 6157
rect 8889 6157 8972 6174
rect 9006 6174 9022 6191
rect 9214 6191 9280 6207
rect 9214 6174 9230 6191
rect 9006 6157 9089 6174
rect 8889 6119 9089 6157
rect 9147 6157 9230 6174
rect 9264 6174 9280 6191
rect 9472 6191 9538 6207
rect 9472 6174 9488 6191
rect 9264 6157 9347 6174
rect 9147 6119 9347 6157
rect 9405 6157 9488 6174
rect 9522 6174 9538 6191
rect 9730 6191 9796 6207
rect 9730 6174 9746 6191
rect 9522 6157 9605 6174
rect 9405 6119 9605 6157
rect 9663 6157 9746 6174
rect 9780 6174 9796 6191
rect 10587 6192 10653 6208
rect 10587 6175 10603 6192
rect 9780 6157 9863 6174
rect 9663 6119 9863 6157
rect 10520 6158 10603 6175
rect 10637 6175 10653 6192
rect 10845 6192 10911 6208
rect 10845 6175 10861 6192
rect 10637 6158 10720 6175
rect 10520 6120 10720 6158
rect 10778 6158 10861 6175
rect 10895 6175 10911 6192
rect 11103 6192 11169 6208
rect 11103 6175 11119 6192
rect 10895 6158 10978 6175
rect 10778 6120 10978 6158
rect 11036 6158 11119 6175
rect 11153 6175 11169 6192
rect 11361 6192 11427 6208
rect 11361 6175 11377 6192
rect 11153 6158 11236 6175
rect 11036 6120 11236 6158
rect 11294 6158 11377 6175
rect 11411 6175 11427 6192
rect 11619 6192 11685 6208
rect 11619 6175 11635 6192
rect 11411 6158 11494 6175
rect 11294 6120 11494 6158
rect 11552 6158 11635 6175
rect 11669 6175 11685 6192
rect 11877 6192 11943 6208
rect 11877 6175 11893 6192
rect 11669 6158 11752 6175
rect 11552 6120 11752 6158
rect 11810 6158 11893 6175
rect 11927 6175 11943 6192
rect 12135 6192 12201 6208
rect 12135 6175 12151 6192
rect 11927 6158 12010 6175
rect 11810 6120 12010 6158
rect 12068 6158 12151 6175
rect 12185 6175 12201 6192
rect 12393 6192 12459 6208
rect 12393 6175 12409 6192
rect 12185 6158 12268 6175
rect 12068 6120 12268 6158
rect 12326 6158 12409 6175
rect 12443 6175 12459 6192
rect 12443 6158 12526 6175
rect 12326 6120 12526 6158
rect 5187 5881 5387 5919
rect 5187 5864 5270 5881
rect 5254 5847 5270 5864
rect 5304 5864 5387 5881
rect 5445 5881 5645 5919
rect 5445 5864 5528 5881
rect 5304 5847 5320 5864
rect 5254 5831 5320 5847
rect 5512 5847 5528 5864
rect 5562 5864 5645 5881
rect 5703 5881 5903 5919
rect 5703 5864 5786 5881
rect 5562 5847 5578 5864
rect 5512 5831 5578 5847
rect 5770 5847 5786 5864
rect 5820 5864 5903 5881
rect 5961 5881 6161 5919
rect 5961 5864 6044 5881
rect 5820 5847 5836 5864
rect 5770 5831 5836 5847
rect 6028 5847 6044 5864
rect 6078 5864 6161 5881
rect 6219 5881 6419 5919
rect 6219 5864 6302 5881
rect 6078 5847 6094 5864
rect 6028 5831 6094 5847
rect 6286 5847 6302 5864
rect 6336 5864 6419 5881
rect 6477 5881 6677 5919
rect 6477 5864 6560 5881
rect 6336 5847 6352 5864
rect 6286 5831 6352 5847
rect 6544 5847 6560 5864
rect 6594 5864 6677 5881
rect 6735 5881 6935 5919
rect 6735 5864 6818 5881
rect 6594 5847 6610 5864
rect 6544 5831 6610 5847
rect 6802 5847 6818 5864
rect 6852 5864 6935 5881
rect 6993 5881 7193 5919
rect 6993 5864 7076 5881
rect 6852 5847 6868 5864
rect 6802 5831 6868 5847
rect 7060 5847 7076 5864
rect 7110 5864 7193 5881
rect 7857 5881 8057 5919
rect 7857 5864 7940 5881
rect 7110 5847 7126 5864
rect 7060 5831 7126 5847
rect 7924 5847 7940 5864
rect 7974 5864 8057 5881
rect 8115 5881 8315 5919
rect 8115 5864 8198 5881
rect 7974 5847 7990 5864
rect 7924 5831 7990 5847
rect 8182 5847 8198 5864
rect 8232 5864 8315 5881
rect 8373 5881 8573 5919
rect 8373 5864 8456 5881
rect 8232 5847 8248 5864
rect 8182 5831 8248 5847
rect 8440 5847 8456 5864
rect 8490 5864 8573 5881
rect 8631 5881 8831 5919
rect 8631 5864 8714 5881
rect 8490 5847 8506 5864
rect 8440 5831 8506 5847
rect 8698 5847 8714 5864
rect 8748 5864 8831 5881
rect 8889 5881 9089 5919
rect 8889 5864 8972 5881
rect 8748 5847 8764 5864
rect 8698 5831 8764 5847
rect 8956 5847 8972 5864
rect 9006 5864 9089 5881
rect 9147 5881 9347 5919
rect 9147 5864 9230 5881
rect 9006 5847 9022 5864
rect 8956 5831 9022 5847
rect 9214 5847 9230 5864
rect 9264 5864 9347 5881
rect 9405 5881 9605 5919
rect 9405 5864 9488 5881
rect 9264 5847 9280 5864
rect 9214 5831 9280 5847
rect 9472 5847 9488 5864
rect 9522 5864 9605 5881
rect 9663 5881 9863 5919
rect 9663 5864 9746 5881
rect 9522 5847 9538 5864
rect 9472 5831 9538 5847
rect 9730 5847 9746 5864
rect 9780 5864 9863 5881
rect 10520 5882 10720 5920
rect 10520 5865 10603 5882
rect 9780 5847 9796 5864
rect 9730 5831 9796 5847
rect 10587 5848 10603 5865
rect 10637 5865 10720 5882
rect 10778 5882 10978 5920
rect 10778 5865 10861 5882
rect 10637 5848 10653 5865
rect 10587 5832 10653 5848
rect 10845 5848 10861 5865
rect 10895 5865 10978 5882
rect 11036 5882 11236 5920
rect 11036 5865 11119 5882
rect 10895 5848 10911 5865
rect 10845 5832 10911 5848
rect 11103 5848 11119 5865
rect 11153 5865 11236 5882
rect 11294 5882 11494 5920
rect 11294 5865 11377 5882
rect 11153 5848 11169 5865
rect 11103 5832 11169 5848
rect 11361 5848 11377 5865
rect 11411 5865 11494 5882
rect 11552 5882 11752 5920
rect 11552 5865 11635 5882
rect 11411 5848 11427 5865
rect 11361 5832 11427 5848
rect 11619 5848 11635 5865
rect 11669 5865 11752 5882
rect 11810 5882 12010 5920
rect 11810 5865 11893 5882
rect 11669 5848 11685 5865
rect 11619 5832 11685 5848
rect 11877 5848 11893 5865
rect 11927 5865 12010 5882
rect 12068 5882 12268 5920
rect 12068 5865 12151 5882
rect 11927 5848 11943 5865
rect 11877 5832 11943 5848
rect 12135 5848 12151 5865
rect 12185 5865 12268 5882
rect 12326 5882 12526 5920
rect 12326 5865 12409 5882
rect 12185 5848 12201 5865
rect 12135 5832 12201 5848
rect 12393 5848 12409 5865
rect 12443 5865 12526 5882
rect 12443 5848 12459 5865
rect 12393 5832 12459 5848
rect 5254 5773 5320 5789
rect 5254 5756 5270 5773
rect 5187 5739 5270 5756
rect 5304 5756 5320 5773
rect 5512 5773 5578 5789
rect 5512 5756 5528 5773
rect 5304 5739 5387 5756
rect 5187 5701 5387 5739
rect 5445 5739 5528 5756
rect 5562 5756 5578 5773
rect 5770 5773 5836 5789
rect 5770 5756 5786 5773
rect 5562 5739 5645 5756
rect 5445 5701 5645 5739
rect 5703 5739 5786 5756
rect 5820 5756 5836 5773
rect 6028 5773 6094 5789
rect 6028 5756 6044 5773
rect 5820 5739 5903 5756
rect 5703 5701 5903 5739
rect 5961 5739 6044 5756
rect 6078 5756 6094 5773
rect 6286 5773 6352 5789
rect 6286 5756 6302 5773
rect 6078 5739 6161 5756
rect 5961 5701 6161 5739
rect 6219 5739 6302 5756
rect 6336 5756 6352 5773
rect 6544 5773 6610 5789
rect 6544 5756 6560 5773
rect 6336 5739 6419 5756
rect 6219 5701 6419 5739
rect 6477 5739 6560 5756
rect 6594 5756 6610 5773
rect 6802 5773 6868 5789
rect 6802 5756 6818 5773
rect 6594 5739 6677 5756
rect 6477 5701 6677 5739
rect 6735 5739 6818 5756
rect 6852 5756 6868 5773
rect 7060 5773 7126 5789
rect 7060 5756 7076 5773
rect 6852 5739 6935 5756
rect 6735 5701 6935 5739
rect 6993 5739 7076 5756
rect 7110 5756 7126 5773
rect 7924 5773 7990 5789
rect 7924 5756 7940 5773
rect 7110 5739 7193 5756
rect 6993 5701 7193 5739
rect 7857 5739 7940 5756
rect 7974 5756 7990 5773
rect 8182 5773 8248 5789
rect 8182 5756 8198 5773
rect 7974 5739 8057 5756
rect 7857 5701 8057 5739
rect 8115 5739 8198 5756
rect 8232 5756 8248 5773
rect 8440 5773 8506 5789
rect 8440 5756 8456 5773
rect 8232 5739 8315 5756
rect 8115 5701 8315 5739
rect 8373 5739 8456 5756
rect 8490 5756 8506 5773
rect 8698 5773 8764 5789
rect 8698 5756 8714 5773
rect 8490 5739 8573 5756
rect 8373 5701 8573 5739
rect 8631 5739 8714 5756
rect 8748 5756 8764 5773
rect 8956 5773 9022 5789
rect 8956 5756 8972 5773
rect 8748 5739 8831 5756
rect 8631 5701 8831 5739
rect 8889 5739 8972 5756
rect 9006 5756 9022 5773
rect 9214 5773 9280 5789
rect 9214 5756 9230 5773
rect 9006 5739 9089 5756
rect 8889 5701 9089 5739
rect 9147 5739 9230 5756
rect 9264 5756 9280 5773
rect 9472 5773 9538 5789
rect 9472 5756 9488 5773
rect 9264 5739 9347 5756
rect 9147 5701 9347 5739
rect 9405 5739 9488 5756
rect 9522 5756 9538 5773
rect 9730 5773 9796 5789
rect 9730 5756 9746 5773
rect 9522 5739 9605 5756
rect 9405 5701 9605 5739
rect 9663 5739 9746 5756
rect 9780 5756 9796 5773
rect 10587 5774 10653 5790
rect 10587 5757 10603 5774
rect 9780 5739 9863 5756
rect 9663 5701 9863 5739
rect 10520 5740 10603 5757
rect 10637 5757 10653 5774
rect 10845 5774 10911 5790
rect 10845 5757 10861 5774
rect 10637 5740 10720 5757
rect 10520 5702 10720 5740
rect 10778 5740 10861 5757
rect 10895 5757 10911 5774
rect 11103 5774 11169 5790
rect 11103 5757 11119 5774
rect 10895 5740 10978 5757
rect 10778 5702 10978 5740
rect 11036 5740 11119 5757
rect 11153 5757 11169 5774
rect 11361 5774 11427 5790
rect 11361 5757 11377 5774
rect 11153 5740 11236 5757
rect 11036 5702 11236 5740
rect 11294 5740 11377 5757
rect 11411 5757 11427 5774
rect 11619 5774 11685 5790
rect 11619 5757 11635 5774
rect 11411 5740 11494 5757
rect 11294 5702 11494 5740
rect 11552 5740 11635 5757
rect 11669 5757 11685 5774
rect 11877 5774 11943 5790
rect 11877 5757 11893 5774
rect 11669 5740 11752 5757
rect 11552 5702 11752 5740
rect 11810 5740 11893 5757
rect 11927 5757 11943 5774
rect 12135 5774 12201 5790
rect 12135 5757 12151 5774
rect 11927 5740 12010 5757
rect 11810 5702 12010 5740
rect 12068 5740 12151 5757
rect 12185 5757 12201 5774
rect 12393 5774 12459 5790
rect 12393 5757 12409 5774
rect 12185 5740 12268 5757
rect 12068 5702 12268 5740
rect 12326 5740 12409 5757
rect 12443 5757 12459 5774
rect 12443 5740 12526 5757
rect 12326 5702 12526 5740
rect 5187 5463 5387 5501
rect 5187 5446 5270 5463
rect 5254 5429 5270 5446
rect 5304 5446 5387 5463
rect 5445 5463 5645 5501
rect 5445 5446 5528 5463
rect 5304 5429 5320 5446
rect 5254 5413 5320 5429
rect 5512 5429 5528 5446
rect 5562 5446 5645 5463
rect 5703 5463 5903 5501
rect 5703 5446 5786 5463
rect 5562 5429 5578 5446
rect 5512 5413 5578 5429
rect 5770 5429 5786 5446
rect 5820 5446 5903 5463
rect 5961 5463 6161 5501
rect 5961 5446 6044 5463
rect 5820 5429 5836 5446
rect 5770 5413 5836 5429
rect 6028 5429 6044 5446
rect 6078 5446 6161 5463
rect 6219 5463 6419 5501
rect 6219 5446 6302 5463
rect 6078 5429 6094 5446
rect 6028 5413 6094 5429
rect 6286 5429 6302 5446
rect 6336 5446 6419 5463
rect 6477 5463 6677 5501
rect 6477 5446 6560 5463
rect 6336 5429 6352 5446
rect 6286 5413 6352 5429
rect 6544 5429 6560 5446
rect 6594 5446 6677 5463
rect 6735 5463 6935 5501
rect 6735 5446 6818 5463
rect 6594 5429 6610 5446
rect 6544 5413 6610 5429
rect 6802 5429 6818 5446
rect 6852 5446 6935 5463
rect 6993 5463 7193 5501
rect 6993 5446 7076 5463
rect 6852 5429 6868 5446
rect 6802 5413 6868 5429
rect 7060 5429 7076 5446
rect 7110 5446 7193 5463
rect 7857 5463 8057 5501
rect 7857 5446 7940 5463
rect 7110 5429 7126 5446
rect 7060 5413 7126 5429
rect 7924 5429 7940 5446
rect 7974 5446 8057 5463
rect 8115 5463 8315 5501
rect 8115 5446 8198 5463
rect 7974 5429 7990 5446
rect 7924 5413 7990 5429
rect 8182 5429 8198 5446
rect 8232 5446 8315 5463
rect 8373 5463 8573 5501
rect 8373 5446 8456 5463
rect 8232 5429 8248 5446
rect 8182 5413 8248 5429
rect 8440 5429 8456 5446
rect 8490 5446 8573 5463
rect 8631 5463 8831 5501
rect 8631 5446 8714 5463
rect 8490 5429 8506 5446
rect 8440 5413 8506 5429
rect 8698 5429 8714 5446
rect 8748 5446 8831 5463
rect 8889 5463 9089 5501
rect 8889 5446 8972 5463
rect 8748 5429 8764 5446
rect 8698 5413 8764 5429
rect 8956 5429 8972 5446
rect 9006 5446 9089 5463
rect 9147 5463 9347 5501
rect 9147 5446 9230 5463
rect 9006 5429 9022 5446
rect 8956 5413 9022 5429
rect 9214 5429 9230 5446
rect 9264 5446 9347 5463
rect 9405 5463 9605 5501
rect 9405 5446 9488 5463
rect 9264 5429 9280 5446
rect 9214 5413 9280 5429
rect 9472 5429 9488 5446
rect 9522 5446 9605 5463
rect 9663 5463 9863 5501
rect 9663 5446 9746 5463
rect 9522 5429 9538 5446
rect 9472 5413 9538 5429
rect 9730 5429 9746 5446
rect 9780 5446 9863 5463
rect 10520 5464 10720 5502
rect 10520 5447 10603 5464
rect 9780 5429 9796 5446
rect 9730 5413 9796 5429
rect 10587 5430 10603 5447
rect 10637 5447 10720 5464
rect 10778 5464 10978 5502
rect 10778 5447 10861 5464
rect 10637 5430 10653 5447
rect 10587 5414 10653 5430
rect 10845 5430 10861 5447
rect 10895 5447 10978 5464
rect 11036 5464 11236 5502
rect 11036 5447 11119 5464
rect 10895 5430 10911 5447
rect 10845 5414 10911 5430
rect 11103 5430 11119 5447
rect 11153 5447 11236 5464
rect 11294 5464 11494 5502
rect 11294 5447 11377 5464
rect 11153 5430 11169 5447
rect 11103 5414 11169 5430
rect 11361 5430 11377 5447
rect 11411 5447 11494 5464
rect 11552 5464 11752 5502
rect 11552 5447 11635 5464
rect 11411 5430 11427 5447
rect 11361 5414 11427 5430
rect 11619 5430 11635 5447
rect 11669 5447 11752 5464
rect 11810 5464 12010 5502
rect 11810 5447 11893 5464
rect 11669 5430 11685 5447
rect 11619 5414 11685 5430
rect 11877 5430 11893 5447
rect 11927 5447 12010 5464
rect 12068 5464 12268 5502
rect 12068 5447 12151 5464
rect 11927 5430 11943 5447
rect 11877 5414 11943 5430
rect 12135 5430 12151 5447
rect 12185 5447 12268 5464
rect 12326 5464 12526 5502
rect 12326 5447 12409 5464
rect 12185 5430 12201 5447
rect 12135 5414 12201 5430
rect 12393 5430 12409 5447
rect 12443 5447 12526 5464
rect 12443 5430 12459 5447
rect 12393 5414 12459 5430
rect 5254 5355 5320 5371
rect 5254 5338 5270 5355
rect 5187 5321 5270 5338
rect 5304 5338 5320 5355
rect 5512 5355 5578 5371
rect 5512 5338 5528 5355
rect 5304 5321 5387 5338
rect 5187 5283 5387 5321
rect 5445 5321 5528 5338
rect 5562 5338 5578 5355
rect 5770 5355 5836 5371
rect 5770 5338 5786 5355
rect 5562 5321 5645 5338
rect 5445 5283 5645 5321
rect 5703 5321 5786 5338
rect 5820 5338 5836 5355
rect 6028 5355 6094 5371
rect 6028 5338 6044 5355
rect 5820 5321 5903 5338
rect 5703 5283 5903 5321
rect 5961 5321 6044 5338
rect 6078 5338 6094 5355
rect 6286 5355 6352 5371
rect 6286 5338 6302 5355
rect 6078 5321 6161 5338
rect 5961 5283 6161 5321
rect 6219 5321 6302 5338
rect 6336 5338 6352 5355
rect 6544 5355 6610 5371
rect 6544 5338 6560 5355
rect 6336 5321 6419 5338
rect 6219 5283 6419 5321
rect 6477 5321 6560 5338
rect 6594 5338 6610 5355
rect 6802 5355 6868 5371
rect 6802 5338 6818 5355
rect 6594 5321 6677 5338
rect 6477 5283 6677 5321
rect 6735 5321 6818 5338
rect 6852 5338 6868 5355
rect 7060 5355 7126 5371
rect 7060 5338 7076 5355
rect 6852 5321 6935 5338
rect 6735 5283 6935 5321
rect 6993 5321 7076 5338
rect 7110 5338 7126 5355
rect 7924 5355 7990 5371
rect 7924 5338 7940 5355
rect 7110 5321 7193 5338
rect 6993 5283 7193 5321
rect 7857 5321 7940 5338
rect 7974 5338 7990 5355
rect 8182 5355 8248 5371
rect 8182 5338 8198 5355
rect 7974 5321 8057 5338
rect 7857 5283 8057 5321
rect 8115 5321 8198 5338
rect 8232 5338 8248 5355
rect 8440 5355 8506 5371
rect 8440 5338 8456 5355
rect 8232 5321 8315 5338
rect 8115 5283 8315 5321
rect 8373 5321 8456 5338
rect 8490 5338 8506 5355
rect 8698 5355 8764 5371
rect 8698 5338 8714 5355
rect 8490 5321 8573 5338
rect 8373 5283 8573 5321
rect 8631 5321 8714 5338
rect 8748 5338 8764 5355
rect 8956 5355 9022 5371
rect 8956 5338 8972 5355
rect 8748 5321 8831 5338
rect 8631 5283 8831 5321
rect 8889 5321 8972 5338
rect 9006 5338 9022 5355
rect 9214 5355 9280 5371
rect 9214 5338 9230 5355
rect 9006 5321 9089 5338
rect 8889 5283 9089 5321
rect 9147 5321 9230 5338
rect 9264 5338 9280 5355
rect 9472 5355 9538 5371
rect 9472 5338 9488 5355
rect 9264 5321 9347 5338
rect 9147 5283 9347 5321
rect 9405 5321 9488 5338
rect 9522 5338 9538 5355
rect 9730 5355 9796 5371
rect 9730 5338 9746 5355
rect 9522 5321 9605 5338
rect 9405 5283 9605 5321
rect 9663 5321 9746 5338
rect 9780 5338 9796 5355
rect 10587 5356 10653 5372
rect 10587 5339 10603 5356
rect 9780 5321 9863 5338
rect 9663 5283 9863 5321
rect 10520 5322 10603 5339
rect 10637 5339 10653 5356
rect 10845 5356 10911 5372
rect 10845 5339 10861 5356
rect 10637 5322 10720 5339
rect 10520 5284 10720 5322
rect 10778 5322 10861 5339
rect 10895 5339 10911 5356
rect 11103 5356 11169 5372
rect 11103 5339 11119 5356
rect 10895 5322 10978 5339
rect 10778 5284 10978 5322
rect 11036 5322 11119 5339
rect 11153 5339 11169 5356
rect 11361 5356 11427 5372
rect 11361 5339 11377 5356
rect 11153 5322 11236 5339
rect 11036 5284 11236 5322
rect 11294 5322 11377 5339
rect 11411 5339 11427 5356
rect 11619 5356 11685 5372
rect 11619 5339 11635 5356
rect 11411 5322 11494 5339
rect 11294 5284 11494 5322
rect 11552 5322 11635 5339
rect 11669 5339 11685 5356
rect 11877 5356 11943 5372
rect 11877 5339 11893 5356
rect 11669 5322 11752 5339
rect 11552 5284 11752 5322
rect 11810 5322 11893 5339
rect 11927 5339 11943 5356
rect 12135 5356 12201 5372
rect 12135 5339 12151 5356
rect 11927 5322 12010 5339
rect 11810 5284 12010 5322
rect 12068 5322 12151 5339
rect 12185 5339 12201 5356
rect 12393 5356 12459 5372
rect 12393 5339 12409 5356
rect 12185 5322 12268 5339
rect 12068 5284 12268 5322
rect 12326 5322 12409 5339
rect 12443 5339 12459 5356
rect 12443 5322 12526 5339
rect 12326 5284 12526 5322
rect 5187 5045 5387 5083
rect 5187 5028 5270 5045
rect 5254 5011 5270 5028
rect 5304 5028 5387 5045
rect 5445 5045 5645 5083
rect 5445 5028 5528 5045
rect 5304 5011 5320 5028
rect 5254 4995 5320 5011
rect 5512 5011 5528 5028
rect 5562 5028 5645 5045
rect 5703 5045 5903 5083
rect 5703 5028 5786 5045
rect 5562 5011 5578 5028
rect 5512 4995 5578 5011
rect 5770 5011 5786 5028
rect 5820 5028 5903 5045
rect 5961 5045 6161 5083
rect 5961 5028 6044 5045
rect 5820 5011 5836 5028
rect 5770 4995 5836 5011
rect 6028 5011 6044 5028
rect 6078 5028 6161 5045
rect 6219 5045 6419 5083
rect 6219 5028 6302 5045
rect 6078 5011 6094 5028
rect 6028 4995 6094 5011
rect 6286 5011 6302 5028
rect 6336 5028 6419 5045
rect 6477 5045 6677 5083
rect 6477 5028 6560 5045
rect 6336 5011 6352 5028
rect 6286 4995 6352 5011
rect 6544 5011 6560 5028
rect 6594 5028 6677 5045
rect 6735 5045 6935 5083
rect 6735 5028 6818 5045
rect 6594 5011 6610 5028
rect 6544 4995 6610 5011
rect 6802 5011 6818 5028
rect 6852 5028 6935 5045
rect 6993 5045 7193 5083
rect 6993 5028 7076 5045
rect 6852 5011 6868 5028
rect 6802 4995 6868 5011
rect 7060 5011 7076 5028
rect 7110 5028 7193 5045
rect 7857 5045 8057 5083
rect 7857 5028 7940 5045
rect 7110 5011 7126 5028
rect 7060 4995 7126 5011
rect 7924 5011 7940 5028
rect 7974 5028 8057 5045
rect 8115 5045 8315 5083
rect 8115 5028 8198 5045
rect 7974 5011 7990 5028
rect 7924 4995 7990 5011
rect 8182 5011 8198 5028
rect 8232 5028 8315 5045
rect 8373 5045 8573 5083
rect 8373 5028 8456 5045
rect 8232 5011 8248 5028
rect 8182 4995 8248 5011
rect 8440 5011 8456 5028
rect 8490 5028 8573 5045
rect 8631 5045 8831 5083
rect 8631 5028 8714 5045
rect 8490 5011 8506 5028
rect 8440 4995 8506 5011
rect 8698 5011 8714 5028
rect 8748 5028 8831 5045
rect 8889 5045 9089 5083
rect 8889 5028 8972 5045
rect 8748 5011 8764 5028
rect 8698 4995 8764 5011
rect 8956 5011 8972 5028
rect 9006 5028 9089 5045
rect 9147 5045 9347 5083
rect 9147 5028 9230 5045
rect 9006 5011 9022 5028
rect 8956 4995 9022 5011
rect 9214 5011 9230 5028
rect 9264 5028 9347 5045
rect 9405 5045 9605 5083
rect 9405 5028 9488 5045
rect 9264 5011 9280 5028
rect 9214 4995 9280 5011
rect 9472 5011 9488 5028
rect 9522 5028 9605 5045
rect 9663 5045 9863 5083
rect 9663 5028 9746 5045
rect 9522 5011 9538 5028
rect 9472 4995 9538 5011
rect 9730 5011 9746 5028
rect 9780 5028 9863 5045
rect 10520 5046 10720 5084
rect 10520 5029 10603 5046
rect 9780 5011 9796 5028
rect 9730 4995 9796 5011
rect 10587 5012 10603 5029
rect 10637 5029 10720 5046
rect 10778 5046 10978 5084
rect 10778 5029 10861 5046
rect 10637 5012 10653 5029
rect 10587 4996 10653 5012
rect 10845 5012 10861 5029
rect 10895 5029 10978 5046
rect 11036 5046 11236 5084
rect 11036 5029 11119 5046
rect 10895 5012 10911 5029
rect 10845 4996 10911 5012
rect 11103 5012 11119 5029
rect 11153 5029 11236 5046
rect 11294 5046 11494 5084
rect 11294 5029 11377 5046
rect 11153 5012 11169 5029
rect 11103 4996 11169 5012
rect 11361 5012 11377 5029
rect 11411 5029 11494 5046
rect 11552 5046 11752 5084
rect 11552 5029 11635 5046
rect 11411 5012 11427 5029
rect 11361 4996 11427 5012
rect 11619 5012 11635 5029
rect 11669 5029 11752 5046
rect 11810 5046 12010 5084
rect 11810 5029 11893 5046
rect 11669 5012 11685 5029
rect 11619 4996 11685 5012
rect 11877 5012 11893 5029
rect 11927 5029 12010 5046
rect 12068 5046 12268 5084
rect 12068 5029 12151 5046
rect 11927 5012 11943 5029
rect 11877 4996 11943 5012
rect 12135 5012 12151 5029
rect 12185 5029 12268 5046
rect 12326 5046 12526 5084
rect 12326 5029 12409 5046
rect 12185 5012 12201 5029
rect 12135 4996 12201 5012
rect 12393 5012 12409 5029
rect 12443 5029 12526 5046
rect 12443 5012 12459 5029
rect 12393 4996 12459 5012
rect 5254 4937 5320 4953
rect 5254 4920 5270 4937
rect 5187 4903 5270 4920
rect 5304 4920 5320 4937
rect 5512 4937 5578 4953
rect 5512 4920 5528 4937
rect 5304 4903 5387 4920
rect 5187 4865 5387 4903
rect 5445 4903 5528 4920
rect 5562 4920 5578 4937
rect 5770 4937 5836 4953
rect 5770 4920 5786 4937
rect 5562 4903 5645 4920
rect 5445 4865 5645 4903
rect 5703 4903 5786 4920
rect 5820 4920 5836 4937
rect 6028 4937 6094 4953
rect 6028 4920 6044 4937
rect 5820 4903 5903 4920
rect 5703 4865 5903 4903
rect 5961 4903 6044 4920
rect 6078 4920 6094 4937
rect 6286 4937 6352 4953
rect 6286 4920 6302 4937
rect 6078 4903 6161 4920
rect 5961 4865 6161 4903
rect 6219 4903 6302 4920
rect 6336 4920 6352 4937
rect 6544 4937 6610 4953
rect 6544 4920 6560 4937
rect 6336 4903 6419 4920
rect 6219 4865 6419 4903
rect 6477 4903 6560 4920
rect 6594 4920 6610 4937
rect 6802 4937 6868 4953
rect 6802 4920 6818 4937
rect 6594 4903 6677 4920
rect 6477 4865 6677 4903
rect 6735 4903 6818 4920
rect 6852 4920 6868 4937
rect 7060 4937 7126 4953
rect 7060 4920 7076 4937
rect 6852 4903 6935 4920
rect 6735 4865 6935 4903
rect 6993 4903 7076 4920
rect 7110 4920 7126 4937
rect 7924 4937 7990 4953
rect 7924 4920 7940 4937
rect 7110 4903 7193 4920
rect 6993 4865 7193 4903
rect 7857 4903 7940 4920
rect 7974 4920 7990 4937
rect 8182 4937 8248 4953
rect 8182 4920 8198 4937
rect 7974 4903 8057 4920
rect 7857 4865 8057 4903
rect 8115 4903 8198 4920
rect 8232 4920 8248 4937
rect 8440 4937 8506 4953
rect 8440 4920 8456 4937
rect 8232 4903 8315 4920
rect 8115 4865 8315 4903
rect 8373 4903 8456 4920
rect 8490 4920 8506 4937
rect 8698 4937 8764 4953
rect 8698 4920 8714 4937
rect 8490 4903 8573 4920
rect 8373 4865 8573 4903
rect 8631 4903 8714 4920
rect 8748 4920 8764 4937
rect 8956 4937 9022 4953
rect 8956 4920 8972 4937
rect 8748 4903 8831 4920
rect 8631 4865 8831 4903
rect 8889 4903 8972 4920
rect 9006 4920 9022 4937
rect 9214 4937 9280 4953
rect 9214 4920 9230 4937
rect 9006 4903 9089 4920
rect 8889 4865 9089 4903
rect 9147 4903 9230 4920
rect 9264 4920 9280 4937
rect 9472 4937 9538 4953
rect 9472 4920 9488 4937
rect 9264 4903 9347 4920
rect 9147 4865 9347 4903
rect 9405 4903 9488 4920
rect 9522 4920 9538 4937
rect 9730 4937 9796 4953
rect 9730 4920 9746 4937
rect 9522 4903 9605 4920
rect 9405 4865 9605 4903
rect 9663 4903 9746 4920
rect 9780 4920 9796 4937
rect 10587 4938 10653 4954
rect 10587 4921 10603 4938
rect 9780 4903 9863 4920
rect 9663 4865 9863 4903
rect 10520 4904 10603 4921
rect 10637 4921 10653 4938
rect 10845 4938 10911 4954
rect 10845 4921 10861 4938
rect 10637 4904 10720 4921
rect 10520 4866 10720 4904
rect 10778 4904 10861 4921
rect 10895 4921 10911 4938
rect 11103 4938 11169 4954
rect 11103 4921 11119 4938
rect 10895 4904 10978 4921
rect 10778 4866 10978 4904
rect 11036 4904 11119 4921
rect 11153 4921 11169 4938
rect 11361 4938 11427 4954
rect 11361 4921 11377 4938
rect 11153 4904 11236 4921
rect 11036 4866 11236 4904
rect 11294 4904 11377 4921
rect 11411 4921 11427 4938
rect 11619 4938 11685 4954
rect 11619 4921 11635 4938
rect 11411 4904 11494 4921
rect 11294 4866 11494 4904
rect 11552 4904 11635 4921
rect 11669 4921 11685 4938
rect 11877 4938 11943 4954
rect 11877 4921 11893 4938
rect 11669 4904 11752 4921
rect 11552 4866 11752 4904
rect 11810 4904 11893 4921
rect 11927 4921 11943 4938
rect 12135 4938 12201 4954
rect 12135 4921 12151 4938
rect 11927 4904 12010 4921
rect 11810 4866 12010 4904
rect 12068 4904 12151 4921
rect 12185 4921 12201 4938
rect 12393 4938 12459 4954
rect 12393 4921 12409 4938
rect 12185 4904 12268 4921
rect 12068 4866 12268 4904
rect 12326 4904 12409 4921
rect 12443 4921 12459 4938
rect 12443 4904 12526 4921
rect 12326 4866 12526 4904
rect 5187 4627 5387 4665
rect 5187 4610 5270 4627
rect 5254 4593 5270 4610
rect 5304 4610 5387 4627
rect 5445 4627 5645 4665
rect 5445 4610 5528 4627
rect 5304 4593 5320 4610
rect 5254 4577 5320 4593
rect 5512 4593 5528 4610
rect 5562 4610 5645 4627
rect 5703 4627 5903 4665
rect 5703 4610 5786 4627
rect 5562 4593 5578 4610
rect 5512 4577 5578 4593
rect 5770 4593 5786 4610
rect 5820 4610 5903 4627
rect 5961 4627 6161 4665
rect 5961 4610 6044 4627
rect 5820 4593 5836 4610
rect 5770 4577 5836 4593
rect 6028 4593 6044 4610
rect 6078 4610 6161 4627
rect 6219 4627 6419 4665
rect 6219 4610 6302 4627
rect 6078 4593 6094 4610
rect 6028 4577 6094 4593
rect 6286 4593 6302 4610
rect 6336 4610 6419 4627
rect 6477 4627 6677 4665
rect 6477 4610 6560 4627
rect 6336 4593 6352 4610
rect 6286 4577 6352 4593
rect 6544 4593 6560 4610
rect 6594 4610 6677 4627
rect 6735 4627 6935 4665
rect 6735 4610 6818 4627
rect 6594 4593 6610 4610
rect 6544 4577 6610 4593
rect 6802 4593 6818 4610
rect 6852 4610 6935 4627
rect 6993 4627 7193 4665
rect 6993 4610 7076 4627
rect 6852 4593 6868 4610
rect 6802 4577 6868 4593
rect 7060 4593 7076 4610
rect 7110 4610 7193 4627
rect 7857 4627 8057 4665
rect 7857 4610 7940 4627
rect 7110 4593 7126 4610
rect 7060 4577 7126 4593
rect 7924 4593 7940 4610
rect 7974 4610 8057 4627
rect 8115 4627 8315 4665
rect 8115 4610 8198 4627
rect 7974 4593 7990 4610
rect 7924 4577 7990 4593
rect 8182 4593 8198 4610
rect 8232 4610 8315 4627
rect 8373 4627 8573 4665
rect 8373 4610 8456 4627
rect 8232 4593 8248 4610
rect 8182 4577 8248 4593
rect 8440 4593 8456 4610
rect 8490 4610 8573 4627
rect 8631 4627 8831 4665
rect 8631 4610 8714 4627
rect 8490 4593 8506 4610
rect 8440 4577 8506 4593
rect 8698 4593 8714 4610
rect 8748 4610 8831 4627
rect 8889 4627 9089 4665
rect 8889 4610 8972 4627
rect 8748 4593 8764 4610
rect 8698 4577 8764 4593
rect 8956 4593 8972 4610
rect 9006 4610 9089 4627
rect 9147 4627 9347 4665
rect 9147 4610 9230 4627
rect 9006 4593 9022 4610
rect 8956 4577 9022 4593
rect 9214 4593 9230 4610
rect 9264 4610 9347 4627
rect 9405 4627 9605 4665
rect 9405 4610 9488 4627
rect 9264 4593 9280 4610
rect 9214 4577 9280 4593
rect 9472 4593 9488 4610
rect 9522 4610 9605 4627
rect 9663 4627 9863 4665
rect 9663 4610 9746 4627
rect 9522 4593 9538 4610
rect 9472 4577 9538 4593
rect 9730 4593 9746 4610
rect 9780 4610 9863 4627
rect 10520 4628 10720 4666
rect 10520 4611 10603 4628
rect 9780 4593 9796 4610
rect 9730 4577 9796 4593
rect 10587 4594 10603 4611
rect 10637 4611 10720 4628
rect 10778 4628 10978 4666
rect 10778 4611 10861 4628
rect 10637 4594 10653 4611
rect 10587 4578 10653 4594
rect 10845 4594 10861 4611
rect 10895 4611 10978 4628
rect 11036 4628 11236 4666
rect 11036 4611 11119 4628
rect 10895 4594 10911 4611
rect 10845 4578 10911 4594
rect 11103 4594 11119 4611
rect 11153 4611 11236 4628
rect 11294 4628 11494 4666
rect 11294 4611 11377 4628
rect 11153 4594 11169 4611
rect 11103 4578 11169 4594
rect 11361 4594 11377 4611
rect 11411 4611 11494 4628
rect 11552 4628 11752 4666
rect 11552 4611 11635 4628
rect 11411 4594 11427 4611
rect 11361 4578 11427 4594
rect 11619 4594 11635 4611
rect 11669 4611 11752 4628
rect 11810 4628 12010 4666
rect 11810 4611 11893 4628
rect 11669 4594 11685 4611
rect 11619 4578 11685 4594
rect 11877 4594 11893 4611
rect 11927 4611 12010 4628
rect 12068 4628 12268 4666
rect 12068 4611 12151 4628
rect 11927 4594 11943 4611
rect 11877 4578 11943 4594
rect 12135 4594 12151 4611
rect 12185 4611 12268 4628
rect 12326 4628 12526 4666
rect 12326 4611 12409 4628
rect 12185 4594 12201 4611
rect 12135 4578 12201 4594
rect 12393 4594 12409 4611
rect 12443 4611 12526 4628
rect 12443 4594 12459 4611
rect 12393 4578 12459 4594
rect 5254 4519 5320 4535
rect 5254 4502 5270 4519
rect 5187 4485 5270 4502
rect 5304 4502 5320 4519
rect 5512 4519 5578 4535
rect 5512 4502 5528 4519
rect 5304 4485 5387 4502
rect 5187 4447 5387 4485
rect 5445 4485 5528 4502
rect 5562 4502 5578 4519
rect 5770 4519 5836 4535
rect 5770 4502 5786 4519
rect 5562 4485 5645 4502
rect 5445 4447 5645 4485
rect 5703 4485 5786 4502
rect 5820 4502 5836 4519
rect 6028 4519 6094 4535
rect 6028 4502 6044 4519
rect 5820 4485 5903 4502
rect 5703 4447 5903 4485
rect 5961 4485 6044 4502
rect 6078 4502 6094 4519
rect 6286 4519 6352 4535
rect 6286 4502 6302 4519
rect 6078 4485 6161 4502
rect 5961 4447 6161 4485
rect 6219 4485 6302 4502
rect 6336 4502 6352 4519
rect 6544 4519 6610 4535
rect 6544 4502 6560 4519
rect 6336 4485 6419 4502
rect 6219 4447 6419 4485
rect 6477 4485 6560 4502
rect 6594 4502 6610 4519
rect 6802 4519 6868 4535
rect 6802 4502 6818 4519
rect 6594 4485 6677 4502
rect 6477 4447 6677 4485
rect 6735 4485 6818 4502
rect 6852 4502 6868 4519
rect 7060 4519 7126 4535
rect 7060 4502 7076 4519
rect 6852 4485 6935 4502
rect 6735 4447 6935 4485
rect 6993 4485 7076 4502
rect 7110 4502 7126 4519
rect 7924 4519 7990 4535
rect 7924 4502 7940 4519
rect 7110 4485 7193 4502
rect 6993 4447 7193 4485
rect 7857 4485 7940 4502
rect 7974 4502 7990 4519
rect 8182 4519 8248 4535
rect 8182 4502 8198 4519
rect 7974 4485 8057 4502
rect 7857 4447 8057 4485
rect 8115 4485 8198 4502
rect 8232 4502 8248 4519
rect 8440 4519 8506 4535
rect 8440 4502 8456 4519
rect 8232 4485 8315 4502
rect 8115 4447 8315 4485
rect 8373 4485 8456 4502
rect 8490 4502 8506 4519
rect 8698 4519 8764 4535
rect 8698 4502 8714 4519
rect 8490 4485 8573 4502
rect 8373 4447 8573 4485
rect 8631 4485 8714 4502
rect 8748 4502 8764 4519
rect 8956 4519 9022 4535
rect 8956 4502 8972 4519
rect 8748 4485 8831 4502
rect 8631 4447 8831 4485
rect 8889 4485 8972 4502
rect 9006 4502 9022 4519
rect 9214 4519 9280 4535
rect 9214 4502 9230 4519
rect 9006 4485 9089 4502
rect 8889 4447 9089 4485
rect 9147 4485 9230 4502
rect 9264 4502 9280 4519
rect 9472 4519 9538 4535
rect 9472 4502 9488 4519
rect 9264 4485 9347 4502
rect 9147 4447 9347 4485
rect 9405 4485 9488 4502
rect 9522 4502 9538 4519
rect 9730 4519 9796 4535
rect 9730 4502 9746 4519
rect 9522 4485 9605 4502
rect 9405 4447 9605 4485
rect 9663 4485 9746 4502
rect 9780 4502 9796 4519
rect 10587 4520 10653 4536
rect 10587 4503 10603 4520
rect 9780 4485 9863 4502
rect 9663 4447 9863 4485
rect 10520 4486 10603 4503
rect 10637 4503 10653 4520
rect 10845 4520 10911 4536
rect 10845 4503 10861 4520
rect 10637 4486 10720 4503
rect 10520 4448 10720 4486
rect 10778 4486 10861 4503
rect 10895 4503 10911 4520
rect 11103 4520 11169 4536
rect 11103 4503 11119 4520
rect 10895 4486 10978 4503
rect 10778 4448 10978 4486
rect 11036 4486 11119 4503
rect 11153 4503 11169 4520
rect 11361 4520 11427 4536
rect 11361 4503 11377 4520
rect 11153 4486 11236 4503
rect 11036 4448 11236 4486
rect 11294 4486 11377 4503
rect 11411 4503 11427 4520
rect 11619 4520 11685 4536
rect 11619 4503 11635 4520
rect 11411 4486 11494 4503
rect 11294 4448 11494 4486
rect 11552 4486 11635 4503
rect 11669 4503 11685 4520
rect 11877 4520 11943 4536
rect 11877 4503 11893 4520
rect 11669 4486 11752 4503
rect 11552 4448 11752 4486
rect 11810 4486 11893 4503
rect 11927 4503 11943 4520
rect 12135 4520 12201 4536
rect 12135 4503 12151 4520
rect 11927 4486 12010 4503
rect 11810 4448 12010 4486
rect 12068 4486 12151 4503
rect 12185 4503 12201 4520
rect 12393 4520 12459 4536
rect 12393 4503 12409 4520
rect 12185 4486 12268 4503
rect 12068 4448 12268 4486
rect 12326 4486 12409 4503
rect 12443 4503 12459 4520
rect 12443 4486 12526 4503
rect 12326 4448 12526 4486
rect 5187 4209 5387 4247
rect 5187 4192 5270 4209
rect 5254 4175 5270 4192
rect 5304 4192 5387 4209
rect 5445 4209 5645 4247
rect 5445 4192 5528 4209
rect 5304 4175 5320 4192
rect 5254 4159 5320 4175
rect 5512 4175 5528 4192
rect 5562 4192 5645 4209
rect 5703 4209 5903 4247
rect 5703 4192 5786 4209
rect 5562 4175 5578 4192
rect 5512 4159 5578 4175
rect 5770 4175 5786 4192
rect 5820 4192 5903 4209
rect 5961 4209 6161 4247
rect 5961 4192 6044 4209
rect 5820 4175 5836 4192
rect 5770 4159 5836 4175
rect 6028 4175 6044 4192
rect 6078 4192 6161 4209
rect 6219 4209 6419 4247
rect 6219 4192 6302 4209
rect 6078 4175 6094 4192
rect 6028 4159 6094 4175
rect 6286 4175 6302 4192
rect 6336 4192 6419 4209
rect 6477 4209 6677 4247
rect 6477 4192 6560 4209
rect 6336 4175 6352 4192
rect 6286 4159 6352 4175
rect 6544 4175 6560 4192
rect 6594 4192 6677 4209
rect 6735 4209 6935 4247
rect 6735 4192 6818 4209
rect 6594 4175 6610 4192
rect 6544 4159 6610 4175
rect 6802 4175 6818 4192
rect 6852 4192 6935 4209
rect 6993 4209 7193 4247
rect 6993 4192 7076 4209
rect 6852 4175 6868 4192
rect 6802 4159 6868 4175
rect 7060 4175 7076 4192
rect 7110 4192 7193 4209
rect 7857 4209 8057 4247
rect 7857 4192 7940 4209
rect 7110 4175 7126 4192
rect 7060 4159 7126 4175
rect 7924 4175 7940 4192
rect 7974 4192 8057 4209
rect 8115 4209 8315 4247
rect 8115 4192 8198 4209
rect 7974 4175 7990 4192
rect 7924 4159 7990 4175
rect 8182 4175 8198 4192
rect 8232 4192 8315 4209
rect 8373 4209 8573 4247
rect 8373 4192 8456 4209
rect 8232 4175 8248 4192
rect 8182 4159 8248 4175
rect 8440 4175 8456 4192
rect 8490 4192 8573 4209
rect 8631 4209 8831 4247
rect 8631 4192 8714 4209
rect 8490 4175 8506 4192
rect 8440 4159 8506 4175
rect 8698 4175 8714 4192
rect 8748 4192 8831 4209
rect 8889 4209 9089 4247
rect 8889 4192 8972 4209
rect 8748 4175 8764 4192
rect 8698 4159 8764 4175
rect 8956 4175 8972 4192
rect 9006 4192 9089 4209
rect 9147 4209 9347 4247
rect 9147 4192 9230 4209
rect 9006 4175 9022 4192
rect 8956 4159 9022 4175
rect 9214 4175 9230 4192
rect 9264 4192 9347 4209
rect 9405 4209 9605 4247
rect 9405 4192 9488 4209
rect 9264 4175 9280 4192
rect 9214 4159 9280 4175
rect 9472 4175 9488 4192
rect 9522 4192 9605 4209
rect 9663 4209 9863 4247
rect 9663 4192 9746 4209
rect 9522 4175 9538 4192
rect 9472 4159 9538 4175
rect 9730 4175 9746 4192
rect 9780 4192 9863 4209
rect 10520 4210 10720 4248
rect 10520 4193 10603 4210
rect 9780 4175 9796 4192
rect 9730 4159 9796 4175
rect 10587 4176 10603 4193
rect 10637 4193 10720 4210
rect 10778 4210 10978 4248
rect 10778 4193 10861 4210
rect 10637 4176 10653 4193
rect 10587 4160 10653 4176
rect 10845 4176 10861 4193
rect 10895 4193 10978 4210
rect 11036 4210 11236 4248
rect 11036 4193 11119 4210
rect 10895 4176 10911 4193
rect 10845 4160 10911 4176
rect 11103 4176 11119 4193
rect 11153 4193 11236 4210
rect 11294 4210 11494 4248
rect 11294 4193 11377 4210
rect 11153 4176 11169 4193
rect 11103 4160 11169 4176
rect 11361 4176 11377 4193
rect 11411 4193 11494 4210
rect 11552 4210 11752 4248
rect 11552 4193 11635 4210
rect 11411 4176 11427 4193
rect 11361 4160 11427 4176
rect 11619 4176 11635 4193
rect 11669 4193 11752 4210
rect 11810 4210 12010 4248
rect 11810 4193 11893 4210
rect 11669 4176 11685 4193
rect 11619 4160 11685 4176
rect 11877 4176 11893 4193
rect 11927 4193 12010 4210
rect 12068 4210 12268 4248
rect 12068 4193 12151 4210
rect 11927 4176 11943 4193
rect 11877 4160 11943 4176
rect 12135 4176 12151 4193
rect 12185 4193 12268 4210
rect 12326 4210 12526 4248
rect 12326 4193 12409 4210
rect 12185 4176 12201 4193
rect 12135 4160 12201 4176
rect 12393 4176 12409 4193
rect 12443 4193 12526 4210
rect 12443 4176 12459 4193
rect 12393 4160 12459 4176
rect 5254 4101 5320 4117
rect 5254 4084 5270 4101
rect 5187 4067 5270 4084
rect 5304 4084 5320 4101
rect 5512 4101 5578 4117
rect 5512 4084 5528 4101
rect 5304 4067 5387 4084
rect 5187 4029 5387 4067
rect 5445 4067 5528 4084
rect 5562 4084 5578 4101
rect 5770 4101 5836 4117
rect 5770 4084 5786 4101
rect 5562 4067 5645 4084
rect 5445 4029 5645 4067
rect 5703 4067 5786 4084
rect 5820 4084 5836 4101
rect 6028 4101 6094 4117
rect 6028 4084 6044 4101
rect 5820 4067 5903 4084
rect 5703 4029 5903 4067
rect 5961 4067 6044 4084
rect 6078 4084 6094 4101
rect 6286 4101 6352 4117
rect 6286 4084 6302 4101
rect 6078 4067 6161 4084
rect 5961 4029 6161 4067
rect 6219 4067 6302 4084
rect 6336 4084 6352 4101
rect 6544 4101 6610 4117
rect 6544 4084 6560 4101
rect 6336 4067 6419 4084
rect 6219 4029 6419 4067
rect 6477 4067 6560 4084
rect 6594 4084 6610 4101
rect 6802 4101 6868 4117
rect 6802 4084 6818 4101
rect 6594 4067 6677 4084
rect 6477 4029 6677 4067
rect 6735 4067 6818 4084
rect 6852 4084 6868 4101
rect 7060 4101 7126 4117
rect 7060 4084 7076 4101
rect 6852 4067 6935 4084
rect 6735 4029 6935 4067
rect 6993 4067 7076 4084
rect 7110 4084 7126 4101
rect 7924 4101 7990 4117
rect 7924 4084 7940 4101
rect 7110 4067 7193 4084
rect 6993 4029 7193 4067
rect 7857 4067 7940 4084
rect 7974 4084 7990 4101
rect 8182 4101 8248 4117
rect 8182 4084 8198 4101
rect 7974 4067 8057 4084
rect 7857 4029 8057 4067
rect 8115 4067 8198 4084
rect 8232 4084 8248 4101
rect 8440 4101 8506 4117
rect 8440 4084 8456 4101
rect 8232 4067 8315 4084
rect 8115 4029 8315 4067
rect 8373 4067 8456 4084
rect 8490 4084 8506 4101
rect 8698 4101 8764 4117
rect 8698 4084 8714 4101
rect 8490 4067 8573 4084
rect 8373 4029 8573 4067
rect 8631 4067 8714 4084
rect 8748 4084 8764 4101
rect 8956 4101 9022 4117
rect 8956 4084 8972 4101
rect 8748 4067 8831 4084
rect 8631 4029 8831 4067
rect 8889 4067 8972 4084
rect 9006 4084 9022 4101
rect 9214 4101 9280 4117
rect 9214 4084 9230 4101
rect 9006 4067 9089 4084
rect 8889 4029 9089 4067
rect 9147 4067 9230 4084
rect 9264 4084 9280 4101
rect 9472 4101 9538 4117
rect 9472 4084 9488 4101
rect 9264 4067 9347 4084
rect 9147 4029 9347 4067
rect 9405 4067 9488 4084
rect 9522 4084 9538 4101
rect 9730 4101 9796 4117
rect 9730 4084 9746 4101
rect 9522 4067 9605 4084
rect 9405 4029 9605 4067
rect 9663 4067 9746 4084
rect 9780 4084 9796 4101
rect 10587 4102 10653 4118
rect 10587 4085 10603 4102
rect 9780 4067 9863 4084
rect 9663 4029 9863 4067
rect 10520 4068 10603 4085
rect 10637 4085 10653 4102
rect 10845 4102 10911 4118
rect 10845 4085 10861 4102
rect 10637 4068 10720 4085
rect 10520 4030 10720 4068
rect 10778 4068 10861 4085
rect 10895 4085 10911 4102
rect 11103 4102 11169 4118
rect 11103 4085 11119 4102
rect 10895 4068 10978 4085
rect 10778 4030 10978 4068
rect 11036 4068 11119 4085
rect 11153 4085 11169 4102
rect 11361 4102 11427 4118
rect 11361 4085 11377 4102
rect 11153 4068 11236 4085
rect 11036 4030 11236 4068
rect 11294 4068 11377 4085
rect 11411 4085 11427 4102
rect 11619 4102 11685 4118
rect 11619 4085 11635 4102
rect 11411 4068 11494 4085
rect 11294 4030 11494 4068
rect 11552 4068 11635 4085
rect 11669 4085 11685 4102
rect 11877 4102 11943 4118
rect 11877 4085 11893 4102
rect 11669 4068 11752 4085
rect 11552 4030 11752 4068
rect 11810 4068 11893 4085
rect 11927 4085 11943 4102
rect 12135 4102 12201 4118
rect 12135 4085 12151 4102
rect 11927 4068 12010 4085
rect 11810 4030 12010 4068
rect 12068 4068 12151 4085
rect 12185 4085 12201 4102
rect 12393 4102 12459 4118
rect 12393 4085 12409 4102
rect 12185 4068 12268 4085
rect 12068 4030 12268 4068
rect 12326 4068 12409 4085
rect 12443 4085 12459 4102
rect 12443 4068 12526 4085
rect 12326 4030 12526 4068
rect 5187 3791 5387 3829
rect 5187 3774 5270 3791
rect 5254 3757 5270 3774
rect 5304 3774 5387 3791
rect 5445 3791 5645 3829
rect 5445 3774 5528 3791
rect 5304 3757 5320 3774
rect 5254 3741 5320 3757
rect 5512 3757 5528 3774
rect 5562 3774 5645 3791
rect 5703 3791 5903 3829
rect 5703 3774 5786 3791
rect 5562 3757 5578 3774
rect 5512 3741 5578 3757
rect 5770 3757 5786 3774
rect 5820 3774 5903 3791
rect 5961 3791 6161 3829
rect 5961 3774 6044 3791
rect 5820 3757 5836 3774
rect 5770 3741 5836 3757
rect 6028 3757 6044 3774
rect 6078 3774 6161 3791
rect 6219 3791 6419 3829
rect 6219 3774 6302 3791
rect 6078 3757 6094 3774
rect 6028 3741 6094 3757
rect 6286 3757 6302 3774
rect 6336 3774 6419 3791
rect 6477 3791 6677 3829
rect 6477 3774 6560 3791
rect 6336 3757 6352 3774
rect 6286 3741 6352 3757
rect 6544 3757 6560 3774
rect 6594 3774 6677 3791
rect 6735 3791 6935 3829
rect 6735 3774 6818 3791
rect 6594 3757 6610 3774
rect 6544 3741 6610 3757
rect 6802 3757 6818 3774
rect 6852 3774 6935 3791
rect 6993 3791 7193 3829
rect 6993 3774 7076 3791
rect 6852 3757 6868 3774
rect 6802 3741 6868 3757
rect 7060 3757 7076 3774
rect 7110 3774 7193 3791
rect 7857 3791 8057 3829
rect 7857 3774 7940 3791
rect 7110 3757 7126 3774
rect 7060 3741 7126 3757
rect 7924 3757 7940 3774
rect 7974 3774 8057 3791
rect 8115 3791 8315 3829
rect 8115 3774 8198 3791
rect 7974 3757 7990 3774
rect 7924 3741 7990 3757
rect 8182 3757 8198 3774
rect 8232 3774 8315 3791
rect 8373 3791 8573 3829
rect 8373 3774 8456 3791
rect 8232 3757 8248 3774
rect 8182 3741 8248 3757
rect 8440 3757 8456 3774
rect 8490 3774 8573 3791
rect 8631 3791 8831 3829
rect 8631 3774 8714 3791
rect 8490 3757 8506 3774
rect 8440 3741 8506 3757
rect 8698 3757 8714 3774
rect 8748 3774 8831 3791
rect 8889 3791 9089 3829
rect 8889 3774 8972 3791
rect 8748 3757 8764 3774
rect 8698 3741 8764 3757
rect 8956 3757 8972 3774
rect 9006 3774 9089 3791
rect 9147 3791 9347 3829
rect 9147 3774 9230 3791
rect 9006 3757 9022 3774
rect 8956 3741 9022 3757
rect 9214 3757 9230 3774
rect 9264 3774 9347 3791
rect 9405 3791 9605 3829
rect 9405 3774 9488 3791
rect 9264 3757 9280 3774
rect 9214 3741 9280 3757
rect 9472 3757 9488 3774
rect 9522 3774 9605 3791
rect 9663 3791 9863 3829
rect 9663 3774 9746 3791
rect 9522 3757 9538 3774
rect 9472 3741 9538 3757
rect 9730 3757 9746 3774
rect 9780 3774 9863 3791
rect 10520 3792 10720 3830
rect 10520 3775 10603 3792
rect 9780 3757 9796 3774
rect 9730 3741 9796 3757
rect 10587 3758 10603 3775
rect 10637 3775 10720 3792
rect 10778 3792 10978 3830
rect 10778 3775 10861 3792
rect 10637 3758 10653 3775
rect 10587 3742 10653 3758
rect 10845 3758 10861 3775
rect 10895 3775 10978 3792
rect 11036 3792 11236 3830
rect 11036 3775 11119 3792
rect 10895 3758 10911 3775
rect 10845 3742 10911 3758
rect 11103 3758 11119 3775
rect 11153 3775 11236 3792
rect 11294 3792 11494 3830
rect 11294 3775 11377 3792
rect 11153 3758 11169 3775
rect 11103 3742 11169 3758
rect 11361 3758 11377 3775
rect 11411 3775 11494 3792
rect 11552 3792 11752 3830
rect 11552 3775 11635 3792
rect 11411 3758 11427 3775
rect 11361 3742 11427 3758
rect 11619 3758 11635 3775
rect 11669 3775 11752 3792
rect 11810 3792 12010 3830
rect 11810 3775 11893 3792
rect 11669 3758 11685 3775
rect 11619 3742 11685 3758
rect 11877 3758 11893 3775
rect 11927 3775 12010 3792
rect 12068 3792 12268 3830
rect 12068 3775 12151 3792
rect 11927 3758 11943 3775
rect 11877 3742 11943 3758
rect 12135 3758 12151 3775
rect 12185 3775 12268 3792
rect 12326 3792 12526 3830
rect 12326 3775 12409 3792
rect 12185 3758 12201 3775
rect 12135 3742 12201 3758
rect 12393 3758 12409 3775
rect 12443 3775 12526 3792
rect 12443 3758 12459 3775
rect 12393 3742 12459 3758
rect 5134 3449 5200 3465
rect 5134 3432 5150 3449
rect 5067 3415 5150 3432
rect 5184 3432 5200 3449
rect 5674 3449 5740 3465
rect 5674 3432 5690 3449
rect 5184 3415 5267 3432
rect 5067 3377 5267 3415
rect 5607 3415 5690 3432
rect 5724 3432 5740 3449
rect 6154 3449 6220 3465
rect 6154 3432 6170 3449
rect 5724 3415 5807 3432
rect 5607 3377 5807 3415
rect 6087 3415 6170 3432
rect 6204 3432 6220 3449
rect 6657 3451 6723 3467
rect 6657 3434 6673 3451
rect 6204 3415 6287 3432
rect 6087 3377 6287 3415
rect 6590 3417 6673 3434
rect 6707 3434 6723 3451
rect 7167 3461 7233 3477
rect 7167 3444 7183 3461
rect 6707 3417 6790 3434
rect 6590 3379 6790 3417
rect 7100 3427 7183 3444
rect 7217 3444 7233 3461
rect 7804 3449 7870 3465
rect 7217 3427 7300 3444
rect 7804 3432 7820 3449
rect 7100 3389 7300 3427
rect 7737 3415 7820 3432
rect 7854 3432 7870 3449
rect 8344 3449 8410 3465
rect 8344 3432 8360 3449
rect 7854 3415 7937 3432
rect 7737 3377 7937 3415
rect 8277 3415 8360 3432
rect 8394 3432 8410 3449
rect 8824 3449 8890 3465
rect 8824 3432 8840 3449
rect 8394 3415 8477 3432
rect 8277 3377 8477 3415
rect 8757 3415 8840 3432
rect 8874 3432 8890 3449
rect 9327 3451 9393 3467
rect 9327 3434 9343 3451
rect 8874 3415 8957 3432
rect 8757 3377 8957 3415
rect 9260 3417 9343 3434
rect 9377 3434 9393 3451
rect 9837 3461 9903 3477
rect 9837 3444 9853 3461
rect 9377 3417 9460 3434
rect 9260 3379 9460 3417
rect 9770 3427 9853 3444
rect 9887 3444 9903 3461
rect 10467 3450 10533 3466
rect 9887 3427 9970 3444
rect 10467 3433 10483 3450
rect 9770 3389 9970 3427
rect 10400 3416 10483 3433
rect 10517 3433 10533 3450
rect 11007 3450 11073 3466
rect 11007 3433 11023 3450
rect 10517 3416 10600 3433
rect 5067 3139 5267 3177
rect 5067 3122 5150 3139
rect 5134 3105 5150 3122
rect 5184 3122 5267 3139
rect 5607 3139 5807 3177
rect 5607 3122 5690 3139
rect 5184 3105 5200 3122
rect 5134 3089 5200 3105
rect 5674 3105 5690 3122
rect 5724 3122 5807 3139
rect 6087 3139 6287 3177
rect 6087 3122 6170 3139
rect 5724 3105 5740 3122
rect 5674 3089 5740 3105
rect 6154 3105 6170 3122
rect 6204 3122 6287 3139
rect 6590 3141 6790 3179
rect 6590 3124 6673 3141
rect 6204 3105 6220 3122
rect 6154 3089 6220 3105
rect 6657 3107 6673 3124
rect 6707 3124 6790 3141
rect 7100 3151 7300 3189
rect 10400 3378 10600 3416
rect 10940 3416 11023 3433
rect 11057 3433 11073 3450
rect 11487 3450 11553 3466
rect 11487 3433 11503 3450
rect 11057 3416 11140 3433
rect 10940 3378 11140 3416
rect 11420 3416 11503 3433
rect 11537 3433 11553 3450
rect 11990 3452 12056 3468
rect 11990 3435 12006 3452
rect 11537 3416 11620 3433
rect 11420 3378 11620 3416
rect 11923 3418 12006 3435
rect 12040 3435 12056 3452
rect 12500 3462 12566 3478
rect 12500 3445 12516 3462
rect 12040 3418 12123 3435
rect 11923 3380 12123 3418
rect 12433 3428 12516 3445
rect 12550 3445 12566 3462
rect 12550 3428 12633 3445
rect 12433 3390 12633 3428
rect 7100 3134 7183 3151
rect 6707 3107 6723 3124
rect 6657 3091 6723 3107
rect 7167 3117 7183 3134
rect 7217 3134 7300 3151
rect 7737 3139 7937 3177
rect 7217 3117 7233 3134
rect 7737 3122 7820 3139
rect 7167 3101 7233 3117
rect 7804 3105 7820 3122
rect 7854 3122 7937 3139
rect 8277 3139 8477 3177
rect 8277 3122 8360 3139
rect 7854 3105 7870 3122
rect 7804 3089 7870 3105
rect 8344 3105 8360 3122
rect 8394 3122 8477 3139
rect 8757 3139 8957 3177
rect 8757 3122 8840 3139
rect 8394 3105 8410 3122
rect 8344 3089 8410 3105
rect 8824 3105 8840 3122
rect 8874 3122 8957 3139
rect 9260 3141 9460 3179
rect 9260 3124 9343 3141
rect 8874 3105 8890 3122
rect 8824 3089 8890 3105
rect 9327 3107 9343 3124
rect 9377 3124 9460 3141
rect 9770 3151 9970 3189
rect 9770 3134 9853 3151
rect 9377 3107 9393 3124
rect 9327 3091 9393 3107
rect 9837 3117 9853 3134
rect 9887 3134 9970 3151
rect 10400 3140 10600 3178
rect 9887 3117 9903 3134
rect 10400 3123 10483 3140
rect 9837 3101 9903 3117
rect 10467 3106 10483 3123
rect 10517 3123 10600 3140
rect 10940 3140 11140 3178
rect 10940 3123 11023 3140
rect 10517 3106 10533 3123
rect 10467 3090 10533 3106
rect 11007 3106 11023 3123
rect 11057 3123 11140 3140
rect 11420 3140 11620 3178
rect 11420 3123 11503 3140
rect 11057 3106 11073 3123
rect 11007 3090 11073 3106
rect 11487 3106 11503 3123
rect 11537 3123 11620 3140
rect 11923 3142 12123 3180
rect 11923 3125 12006 3142
rect 11537 3106 11553 3123
rect 11487 3090 11553 3106
rect 11990 3108 12006 3125
rect 12040 3125 12123 3142
rect 12433 3152 12633 3190
rect 12433 3135 12516 3152
rect 12040 3108 12056 3125
rect 11990 3092 12056 3108
rect 12500 3118 12516 3135
rect 12550 3135 12633 3152
rect 12550 3118 12566 3135
rect 12500 3102 12566 3118
rect 5412 1930 5528 1958
rect 5412 1892 5436 1930
rect 5502 1892 5528 1930
rect 6064 1923 6250 1939
rect 6064 1906 6080 1923
rect 5412 1842 5528 1892
rect 5757 1889 6080 1906
rect 6234 1906 6250 1923
rect 6798 1929 6914 1957
rect 6234 1889 6557 1906
rect 5757 1842 6557 1889
rect 6798 1891 6822 1929
rect 6888 1891 6914 1929
rect 6798 1841 6914 1891
rect 7168 1929 7284 1957
rect 7168 1891 7192 1929
rect 7258 1891 7284 1929
rect 7168 1841 7284 1891
rect 7590 1929 7706 1957
rect 7590 1891 7614 1929
rect 7680 1891 7706 1929
rect 7590 1841 7706 1891
rect 8012 1929 8128 1957
rect 8012 1891 8036 1929
rect 8102 1891 8128 1929
rect 8741 1923 8927 1939
rect 8741 1906 8757 1923
rect 8012 1841 8128 1891
rect 8434 1889 8757 1906
rect 8911 1906 8927 1923
rect 9512 1933 9628 1961
rect 8911 1889 9234 1906
rect 8434 1842 9234 1889
rect 9512 1895 9536 1933
rect 9602 1895 9628 1933
rect 9512 1845 9628 1895
rect 9882 1933 9998 1961
rect 9882 1895 9906 1933
rect 9972 1895 9998 1933
rect 9882 1845 9998 1895
rect 10304 1933 10420 1961
rect 10304 1895 10328 1933
rect 10394 1895 10420 1933
rect 10304 1845 10420 1895
rect 10726 1933 10842 1961
rect 10726 1895 10750 1933
rect 10816 1895 10842 1933
rect 11405 1924 11591 1940
rect 11405 1907 11421 1924
rect 10726 1845 10842 1895
rect 11098 1890 11421 1907
rect 11575 1907 11591 1924
rect 12110 1930 12226 1958
rect 11575 1890 11898 1907
rect 5412 1668 5528 1732
rect 5757 1685 6557 1732
rect 11098 1843 11898 1890
rect 12110 1892 12134 1930
rect 12200 1892 12226 1930
rect 5757 1668 6080 1685
rect 6064 1651 6080 1668
rect 6234 1668 6557 1685
rect 6234 1651 6250 1668
rect 6798 1667 6914 1731
rect 7168 1667 7284 1731
rect 7590 1667 7706 1731
rect 8012 1667 8128 1731
rect 8434 1685 9234 1732
rect 8434 1668 8757 1685
rect 6064 1635 6250 1651
rect 8741 1651 8757 1668
rect 8911 1668 9234 1685
rect 9512 1671 9628 1735
rect 9882 1671 9998 1735
rect 10304 1671 10420 1735
rect 10726 1671 10842 1735
rect 12110 1842 12226 1892
rect 11098 1686 11898 1733
rect 11098 1669 11421 1686
rect 8911 1651 8927 1668
rect 8741 1635 8927 1651
rect 11405 1652 11421 1669
rect 11575 1669 11898 1686
rect 11575 1652 11591 1669
rect 12110 1668 12226 1732
rect 11405 1636 11591 1652
rect 5254 892 5320 908
rect 5254 875 5270 892
rect 5187 858 5270 875
rect 5304 875 5320 892
rect 5512 892 5578 908
rect 5512 875 5528 892
rect 5304 858 5387 875
rect 5187 820 5387 858
rect 5445 858 5528 875
rect 5562 875 5578 892
rect 5770 892 5836 908
rect 5770 875 5786 892
rect 5562 858 5645 875
rect 5445 820 5645 858
rect 5703 858 5786 875
rect 5820 875 5836 892
rect 6028 892 6094 908
rect 6028 875 6044 892
rect 5820 858 5903 875
rect 5703 820 5903 858
rect 5961 858 6044 875
rect 6078 875 6094 892
rect 6286 892 6352 908
rect 6286 875 6302 892
rect 6078 858 6161 875
rect 5961 820 6161 858
rect 6219 858 6302 875
rect 6336 875 6352 892
rect 6544 892 6610 908
rect 6544 875 6560 892
rect 6336 858 6419 875
rect 6219 820 6419 858
rect 6477 858 6560 875
rect 6594 875 6610 892
rect 6802 892 6868 908
rect 6802 875 6818 892
rect 6594 858 6677 875
rect 6477 820 6677 858
rect 6735 858 6818 875
rect 6852 875 6868 892
rect 7060 892 7126 908
rect 7060 875 7076 892
rect 6852 858 6935 875
rect 6735 820 6935 858
rect 6993 858 7076 875
rect 7110 875 7126 892
rect 7924 892 7990 908
rect 7924 875 7940 892
rect 7110 858 7193 875
rect 6993 820 7193 858
rect 7857 858 7940 875
rect 7974 875 7990 892
rect 8182 892 8248 908
rect 8182 875 8198 892
rect 7974 858 8057 875
rect 7857 820 8057 858
rect 8115 858 8198 875
rect 8232 875 8248 892
rect 8440 892 8506 908
rect 8440 875 8456 892
rect 8232 858 8315 875
rect 8115 820 8315 858
rect 8373 858 8456 875
rect 8490 875 8506 892
rect 8698 892 8764 908
rect 8698 875 8714 892
rect 8490 858 8573 875
rect 8373 820 8573 858
rect 8631 858 8714 875
rect 8748 875 8764 892
rect 8956 892 9022 908
rect 8956 875 8972 892
rect 8748 858 8831 875
rect 8631 820 8831 858
rect 8889 858 8972 875
rect 9006 875 9022 892
rect 9214 892 9280 908
rect 9214 875 9230 892
rect 9006 858 9089 875
rect 8889 820 9089 858
rect 9147 858 9230 875
rect 9264 875 9280 892
rect 9472 892 9538 908
rect 9472 875 9488 892
rect 9264 858 9347 875
rect 9147 820 9347 858
rect 9405 858 9488 875
rect 9522 875 9538 892
rect 9730 892 9796 908
rect 9730 875 9746 892
rect 9522 858 9605 875
rect 9405 820 9605 858
rect 9663 858 9746 875
rect 9780 875 9796 892
rect 10587 893 10653 909
rect 10587 876 10603 893
rect 9780 858 9863 875
rect 9663 820 9863 858
rect 10520 859 10603 876
rect 10637 876 10653 893
rect 10845 893 10911 909
rect 10845 876 10861 893
rect 10637 859 10720 876
rect 10520 821 10720 859
rect 10778 859 10861 876
rect 10895 876 10911 893
rect 11103 893 11169 909
rect 11103 876 11119 893
rect 10895 859 10978 876
rect 10778 821 10978 859
rect 11036 859 11119 876
rect 11153 876 11169 893
rect 11361 893 11427 909
rect 11361 876 11377 893
rect 11153 859 11236 876
rect 11036 821 11236 859
rect 11294 859 11377 876
rect 11411 876 11427 893
rect 11619 893 11685 909
rect 11619 876 11635 893
rect 11411 859 11494 876
rect 11294 821 11494 859
rect 11552 859 11635 876
rect 11669 876 11685 893
rect 11877 893 11943 909
rect 11877 876 11893 893
rect 11669 859 11752 876
rect 11552 821 11752 859
rect 11810 859 11893 876
rect 11927 876 11943 893
rect 12135 893 12201 909
rect 12135 876 12151 893
rect 11927 859 12010 876
rect 11810 821 12010 859
rect 12068 859 12151 876
rect 12185 876 12201 893
rect 12393 893 12459 909
rect 12393 876 12409 893
rect 12185 859 12268 876
rect 12068 821 12268 859
rect 12326 859 12409 876
rect 12443 876 12459 893
rect 12443 859 12526 876
rect 12326 821 12526 859
rect 5187 582 5387 620
rect 5187 565 5270 582
rect 5254 548 5270 565
rect 5304 565 5387 582
rect 5445 582 5645 620
rect 5445 565 5528 582
rect 5304 548 5320 565
rect 5254 532 5320 548
rect 5512 548 5528 565
rect 5562 565 5645 582
rect 5703 582 5903 620
rect 5703 565 5786 582
rect 5562 548 5578 565
rect 5512 532 5578 548
rect 5770 548 5786 565
rect 5820 565 5903 582
rect 5961 582 6161 620
rect 5961 565 6044 582
rect 5820 548 5836 565
rect 5770 532 5836 548
rect 6028 548 6044 565
rect 6078 565 6161 582
rect 6219 582 6419 620
rect 6219 565 6302 582
rect 6078 548 6094 565
rect 6028 532 6094 548
rect 6286 548 6302 565
rect 6336 565 6419 582
rect 6477 582 6677 620
rect 6477 565 6560 582
rect 6336 548 6352 565
rect 6286 532 6352 548
rect 6544 548 6560 565
rect 6594 565 6677 582
rect 6735 582 6935 620
rect 6735 565 6818 582
rect 6594 548 6610 565
rect 6544 532 6610 548
rect 6802 548 6818 565
rect 6852 565 6935 582
rect 6993 582 7193 620
rect 6993 565 7076 582
rect 6852 548 6868 565
rect 6802 532 6868 548
rect 7060 548 7076 565
rect 7110 565 7193 582
rect 7857 582 8057 620
rect 7857 565 7940 582
rect 7110 548 7126 565
rect 7060 532 7126 548
rect 7924 548 7940 565
rect 7974 565 8057 582
rect 8115 582 8315 620
rect 8115 565 8198 582
rect 7974 548 7990 565
rect 7924 532 7990 548
rect 8182 548 8198 565
rect 8232 565 8315 582
rect 8373 582 8573 620
rect 8373 565 8456 582
rect 8232 548 8248 565
rect 8182 532 8248 548
rect 8440 548 8456 565
rect 8490 565 8573 582
rect 8631 582 8831 620
rect 8631 565 8714 582
rect 8490 548 8506 565
rect 8440 532 8506 548
rect 8698 548 8714 565
rect 8748 565 8831 582
rect 8889 582 9089 620
rect 8889 565 8972 582
rect 8748 548 8764 565
rect 8698 532 8764 548
rect 8956 548 8972 565
rect 9006 565 9089 582
rect 9147 582 9347 620
rect 9147 565 9230 582
rect 9006 548 9022 565
rect 8956 532 9022 548
rect 9214 548 9230 565
rect 9264 565 9347 582
rect 9405 582 9605 620
rect 9405 565 9488 582
rect 9264 548 9280 565
rect 9214 532 9280 548
rect 9472 548 9488 565
rect 9522 565 9605 582
rect 9663 582 9863 620
rect 9663 565 9746 582
rect 9522 548 9538 565
rect 9472 532 9538 548
rect 9730 548 9746 565
rect 9780 565 9863 582
rect 10520 583 10720 621
rect 10520 566 10603 583
rect 9780 548 9796 565
rect 9730 532 9796 548
rect 10587 549 10603 566
rect 10637 566 10720 583
rect 10778 583 10978 621
rect 10778 566 10861 583
rect 10637 549 10653 566
rect 10587 533 10653 549
rect 10845 549 10861 566
rect 10895 566 10978 583
rect 11036 583 11236 621
rect 11036 566 11119 583
rect 10895 549 10911 566
rect 10845 533 10911 549
rect 11103 549 11119 566
rect 11153 566 11236 583
rect 11294 583 11494 621
rect 11294 566 11377 583
rect 11153 549 11169 566
rect 11103 533 11169 549
rect 11361 549 11377 566
rect 11411 566 11494 583
rect 11552 583 11752 621
rect 11552 566 11635 583
rect 11411 549 11427 566
rect 11361 533 11427 549
rect 11619 549 11635 566
rect 11669 566 11752 583
rect 11810 583 12010 621
rect 11810 566 11893 583
rect 11669 549 11685 566
rect 11619 533 11685 549
rect 11877 549 11893 566
rect 11927 566 12010 583
rect 12068 583 12268 621
rect 12068 566 12151 583
rect 11927 549 11943 566
rect 11877 533 11943 549
rect 12135 549 12151 566
rect 12185 566 12268 583
rect 12326 583 12526 621
rect 12326 566 12409 583
rect 12185 549 12201 566
rect 12135 533 12201 549
rect 12393 549 12409 566
rect 12443 566 12526 583
rect 12443 549 12459 566
rect 12393 533 12459 549
rect 5254 474 5320 490
rect 5254 457 5270 474
rect 5187 440 5270 457
rect 5304 457 5320 474
rect 5512 474 5578 490
rect 5512 457 5528 474
rect 5304 440 5387 457
rect 5187 402 5387 440
rect 5445 440 5528 457
rect 5562 457 5578 474
rect 5770 474 5836 490
rect 5770 457 5786 474
rect 5562 440 5645 457
rect 5445 402 5645 440
rect 5703 440 5786 457
rect 5820 457 5836 474
rect 6028 474 6094 490
rect 6028 457 6044 474
rect 5820 440 5903 457
rect 5703 402 5903 440
rect 5961 440 6044 457
rect 6078 457 6094 474
rect 6286 474 6352 490
rect 6286 457 6302 474
rect 6078 440 6161 457
rect 5961 402 6161 440
rect 6219 440 6302 457
rect 6336 457 6352 474
rect 6544 474 6610 490
rect 6544 457 6560 474
rect 6336 440 6419 457
rect 6219 402 6419 440
rect 6477 440 6560 457
rect 6594 457 6610 474
rect 6802 474 6868 490
rect 6802 457 6818 474
rect 6594 440 6677 457
rect 6477 402 6677 440
rect 6735 440 6818 457
rect 6852 457 6868 474
rect 7060 474 7126 490
rect 7060 457 7076 474
rect 6852 440 6935 457
rect 6735 402 6935 440
rect 6993 440 7076 457
rect 7110 457 7126 474
rect 7924 474 7990 490
rect 7924 457 7940 474
rect 7110 440 7193 457
rect 6993 402 7193 440
rect 7857 440 7940 457
rect 7974 457 7990 474
rect 8182 474 8248 490
rect 8182 457 8198 474
rect 7974 440 8057 457
rect 7857 402 8057 440
rect 8115 440 8198 457
rect 8232 457 8248 474
rect 8440 474 8506 490
rect 8440 457 8456 474
rect 8232 440 8315 457
rect 8115 402 8315 440
rect 8373 440 8456 457
rect 8490 457 8506 474
rect 8698 474 8764 490
rect 8698 457 8714 474
rect 8490 440 8573 457
rect 8373 402 8573 440
rect 8631 440 8714 457
rect 8748 457 8764 474
rect 8956 474 9022 490
rect 8956 457 8972 474
rect 8748 440 8831 457
rect 8631 402 8831 440
rect 8889 440 8972 457
rect 9006 457 9022 474
rect 9214 474 9280 490
rect 9214 457 9230 474
rect 9006 440 9089 457
rect 8889 402 9089 440
rect 9147 440 9230 457
rect 9264 457 9280 474
rect 9472 474 9538 490
rect 9472 457 9488 474
rect 9264 440 9347 457
rect 9147 402 9347 440
rect 9405 440 9488 457
rect 9522 457 9538 474
rect 9730 474 9796 490
rect 9730 457 9746 474
rect 9522 440 9605 457
rect 9405 402 9605 440
rect 9663 440 9746 457
rect 9780 457 9796 474
rect 10587 475 10653 491
rect 10587 458 10603 475
rect 9780 440 9863 457
rect 9663 402 9863 440
rect 10520 441 10603 458
rect 10637 458 10653 475
rect 10845 475 10911 491
rect 10845 458 10861 475
rect 10637 441 10720 458
rect 10520 403 10720 441
rect 10778 441 10861 458
rect 10895 458 10911 475
rect 11103 475 11169 491
rect 11103 458 11119 475
rect 10895 441 10978 458
rect 10778 403 10978 441
rect 11036 441 11119 458
rect 11153 458 11169 475
rect 11361 475 11427 491
rect 11361 458 11377 475
rect 11153 441 11236 458
rect 11036 403 11236 441
rect 11294 441 11377 458
rect 11411 458 11427 475
rect 11619 475 11685 491
rect 11619 458 11635 475
rect 11411 441 11494 458
rect 11294 403 11494 441
rect 11552 441 11635 458
rect 11669 458 11685 475
rect 11877 475 11943 491
rect 11877 458 11893 475
rect 11669 441 11752 458
rect 11552 403 11752 441
rect 11810 441 11893 458
rect 11927 458 11943 475
rect 12135 475 12201 491
rect 12135 458 12151 475
rect 11927 441 12010 458
rect 11810 403 12010 441
rect 12068 441 12151 458
rect 12185 458 12201 475
rect 12393 475 12459 491
rect 12393 458 12409 475
rect 12185 441 12268 458
rect 12068 403 12268 441
rect 12326 441 12409 458
rect 12443 458 12459 475
rect 12443 441 12526 458
rect 12326 403 12526 441
rect 5187 164 5387 202
rect 5187 147 5270 164
rect 5254 130 5270 147
rect 5304 147 5387 164
rect 5445 164 5645 202
rect 5445 147 5528 164
rect 5304 130 5320 147
rect 5254 114 5320 130
rect 5512 130 5528 147
rect 5562 147 5645 164
rect 5703 164 5903 202
rect 5703 147 5786 164
rect 5562 130 5578 147
rect 5512 114 5578 130
rect 5770 130 5786 147
rect 5820 147 5903 164
rect 5961 164 6161 202
rect 5961 147 6044 164
rect 5820 130 5836 147
rect 5770 114 5836 130
rect 6028 130 6044 147
rect 6078 147 6161 164
rect 6219 164 6419 202
rect 6219 147 6302 164
rect 6078 130 6094 147
rect 6028 114 6094 130
rect 6286 130 6302 147
rect 6336 147 6419 164
rect 6477 164 6677 202
rect 6477 147 6560 164
rect 6336 130 6352 147
rect 6286 114 6352 130
rect 6544 130 6560 147
rect 6594 147 6677 164
rect 6735 164 6935 202
rect 6735 147 6818 164
rect 6594 130 6610 147
rect 6544 114 6610 130
rect 6802 130 6818 147
rect 6852 147 6935 164
rect 6993 164 7193 202
rect 6993 147 7076 164
rect 6852 130 6868 147
rect 6802 114 6868 130
rect 7060 130 7076 147
rect 7110 147 7193 164
rect 7857 164 8057 202
rect 7857 147 7940 164
rect 7110 130 7126 147
rect 7060 114 7126 130
rect 7924 130 7940 147
rect 7974 147 8057 164
rect 8115 164 8315 202
rect 8115 147 8198 164
rect 7974 130 7990 147
rect 7924 114 7990 130
rect 8182 130 8198 147
rect 8232 147 8315 164
rect 8373 164 8573 202
rect 8373 147 8456 164
rect 8232 130 8248 147
rect 8182 114 8248 130
rect 8440 130 8456 147
rect 8490 147 8573 164
rect 8631 164 8831 202
rect 8631 147 8714 164
rect 8490 130 8506 147
rect 8440 114 8506 130
rect 8698 130 8714 147
rect 8748 147 8831 164
rect 8889 164 9089 202
rect 8889 147 8972 164
rect 8748 130 8764 147
rect 8698 114 8764 130
rect 8956 130 8972 147
rect 9006 147 9089 164
rect 9147 164 9347 202
rect 9147 147 9230 164
rect 9006 130 9022 147
rect 8956 114 9022 130
rect 9214 130 9230 147
rect 9264 147 9347 164
rect 9405 164 9605 202
rect 9405 147 9488 164
rect 9264 130 9280 147
rect 9214 114 9280 130
rect 9472 130 9488 147
rect 9522 147 9605 164
rect 9663 164 9863 202
rect 9663 147 9746 164
rect 9522 130 9538 147
rect 9472 114 9538 130
rect 9730 130 9746 147
rect 9780 147 9863 164
rect 10520 165 10720 203
rect 10520 148 10603 165
rect 9780 130 9796 147
rect 9730 114 9796 130
rect 10587 131 10603 148
rect 10637 148 10720 165
rect 10778 165 10978 203
rect 10778 148 10861 165
rect 10637 131 10653 148
rect 10587 115 10653 131
rect 10845 131 10861 148
rect 10895 148 10978 165
rect 11036 165 11236 203
rect 11036 148 11119 165
rect 10895 131 10911 148
rect 10845 115 10911 131
rect 11103 131 11119 148
rect 11153 148 11236 165
rect 11294 165 11494 203
rect 11294 148 11377 165
rect 11153 131 11169 148
rect 11103 115 11169 131
rect 11361 131 11377 148
rect 11411 148 11494 165
rect 11552 165 11752 203
rect 11552 148 11635 165
rect 11411 131 11427 148
rect 11361 115 11427 131
rect 11619 131 11635 148
rect 11669 148 11752 165
rect 11810 165 12010 203
rect 11810 148 11893 165
rect 11669 131 11685 148
rect 11619 115 11685 131
rect 11877 131 11893 148
rect 11927 148 12010 165
rect 12068 165 12268 203
rect 12068 148 12151 165
rect 11927 131 11943 148
rect 11877 115 11943 131
rect 12135 131 12151 148
rect 12185 148 12268 165
rect 12326 165 12526 203
rect 12326 148 12409 165
rect 12185 131 12201 148
rect 12135 115 12201 131
rect 12393 131 12409 148
rect 12443 148 12526 165
rect 12443 131 12459 148
rect 12393 115 12459 131
rect 5254 56 5320 72
rect 5254 39 5270 56
rect 5187 22 5270 39
rect 5304 39 5320 56
rect 5512 56 5578 72
rect 5512 39 5528 56
rect 5304 22 5387 39
rect 5187 -16 5387 22
rect 5445 22 5528 39
rect 5562 39 5578 56
rect 5770 56 5836 72
rect 5770 39 5786 56
rect 5562 22 5645 39
rect 5445 -16 5645 22
rect 5703 22 5786 39
rect 5820 39 5836 56
rect 6028 56 6094 72
rect 6028 39 6044 56
rect 5820 22 5903 39
rect 5703 -16 5903 22
rect 5961 22 6044 39
rect 6078 39 6094 56
rect 6286 56 6352 72
rect 6286 39 6302 56
rect 6078 22 6161 39
rect 5961 -16 6161 22
rect 6219 22 6302 39
rect 6336 39 6352 56
rect 6544 56 6610 72
rect 6544 39 6560 56
rect 6336 22 6419 39
rect 6219 -16 6419 22
rect 6477 22 6560 39
rect 6594 39 6610 56
rect 6802 56 6868 72
rect 6802 39 6818 56
rect 6594 22 6677 39
rect 6477 -16 6677 22
rect 6735 22 6818 39
rect 6852 39 6868 56
rect 7060 56 7126 72
rect 7060 39 7076 56
rect 6852 22 6935 39
rect 6735 -16 6935 22
rect 6993 22 7076 39
rect 7110 39 7126 56
rect 7924 56 7990 72
rect 7924 39 7940 56
rect 7110 22 7193 39
rect 6993 -16 7193 22
rect 7857 22 7940 39
rect 7974 39 7990 56
rect 8182 56 8248 72
rect 8182 39 8198 56
rect 7974 22 8057 39
rect 7857 -16 8057 22
rect 8115 22 8198 39
rect 8232 39 8248 56
rect 8440 56 8506 72
rect 8440 39 8456 56
rect 8232 22 8315 39
rect 8115 -16 8315 22
rect 8373 22 8456 39
rect 8490 39 8506 56
rect 8698 56 8764 72
rect 8698 39 8714 56
rect 8490 22 8573 39
rect 8373 -16 8573 22
rect 8631 22 8714 39
rect 8748 39 8764 56
rect 8956 56 9022 72
rect 8956 39 8972 56
rect 8748 22 8831 39
rect 8631 -16 8831 22
rect 8889 22 8972 39
rect 9006 39 9022 56
rect 9214 56 9280 72
rect 9214 39 9230 56
rect 9006 22 9089 39
rect 8889 -16 9089 22
rect 9147 22 9230 39
rect 9264 39 9280 56
rect 9472 56 9538 72
rect 9472 39 9488 56
rect 9264 22 9347 39
rect 9147 -16 9347 22
rect 9405 22 9488 39
rect 9522 39 9538 56
rect 9730 56 9796 72
rect 9730 39 9746 56
rect 9522 22 9605 39
rect 9405 -16 9605 22
rect 9663 22 9746 39
rect 9780 39 9796 56
rect 10587 57 10653 73
rect 10587 40 10603 57
rect 9780 22 9863 39
rect 9663 -16 9863 22
rect 10520 23 10603 40
rect 10637 40 10653 57
rect 10845 57 10911 73
rect 10845 40 10861 57
rect 10637 23 10720 40
rect 10520 -15 10720 23
rect 10778 23 10861 40
rect 10895 40 10911 57
rect 11103 57 11169 73
rect 11103 40 11119 57
rect 10895 23 10978 40
rect 10778 -15 10978 23
rect 11036 23 11119 40
rect 11153 40 11169 57
rect 11361 57 11427 73
rect 11361 40 11377 57
rect 11153 23 11236 40
rect 11036 -15 11236 23
rect 11294 23 11377 40
rect 11411 40 11427 57
rect 11619 57 11685 73
rect 11619 40 11635 57
rect 11411 23 11494 40
rect 11294 -15 11494 23
rect 11552 23 11635 40
rect 11669 40 11685 57
rect 11877 57 11943 73
rect 11877 40 11893 57
rect 11669 23 11752 40
rect 11552 -15 11752 23
rect 11810 23 11893 40
rect 11927 40 11943 57
rect 12135 57 12201 73
rect 12135 40 12151 57
rect 11927 23 12010 40
rect 11810 -15 12010 23
rect 12068 23 12151 40
rect 12185 40 12201 57
rect 12393 57 12459 73
rect 12393 40 12409 57
rect 12185 23 12268 40
rect 12068 -15 12268 23
rect 12326 23 12409 40
rect 12443 40 12459 57
rect 12443 23 12526 40
rect 12326 -15 12526 23
rect 5187 -254 5387 -216
rect 5187 -271 5270 -254
rect 5254 -288 5270 -271
rect 5304 -271 5387 -254
rect 5445 -254 5645 -216
rect 5445 -271 5528 -254
rect 5304 -288 5320 -271
rect 5254 -304 5320 -288
rect 5512 -288 5528 -271
rect 5562 -271 5645 -254
rect 5703 -254 5903 -216
rect 5703 -271 5786 -254
rect 5562 -288 5578 -271
rect 5512 -304 5578 -288
rect 5770 -288 5786 -271
rect 5820 -271 5903 -254
rect 5961 -254 6161 -216
rect 5961 -271 6044 -254
rect 5820 -288 5836 -271
rect 5770 -304 5836 -288
rect 6028 -288 6044 -271
rect 6078 -271 6161 -254
rect 6219 -254 6419 -216
rect 6219 -271 6302 -254
rect 6078 -288 6094 -271
rect 6028 -304 6094 -288
rect 6286 -288 6302 -271
rect 6336 -271 6419 -254
rect 6477 -254 6677 -216
rect 6477 -271 6560 -254
rect 6336 -288 6352 -271
rect 6286 -304 6352 -288
rect 6544 -288 6560 -271
rect 6594 -271 6677 -254
rect 6735 -254 6935 -216
rect 6735 -271 6818 -254
rect 6594 -288 6610 -271
rect 6544 -304 6610 -288
rect 6802 -288 6818 -271
rect 6852 -271 6935 -254
rect 6993 -254 7193 -216
rect 6993 -271 7076 -254
rect 6852 -288 6868 -271
rect 6802 -304 6868 -288
rect 7060 -288 7076 -271
rect 7110 -271 7193 -254
rect 7857 -254 8057 -216
rect 7857 -271 7940 -254
rect 7110 -288 7126 -271
rect 7060 -304 7126 -288
rect 7924 -288 7940 -271
rect 7974 -271 8057 -254
rect 8115 -254 8315 -216
rect 8115 -271 8198 -254
rect 7974 -288 7990 -271
rect 7924 -304 7990 -288
rect 8182 -288 8198 -271
rect 8232 -271 8315 -254
rect 8373 -254 8573 -216
rect 8373 -271 8456 -254
rect 8232 -288 8248 -271
rect 8182 -304 8248 -288
rect 8440 -288 8456 -271
rect 8490 -271 8573 -254
rect 8631 -254 8831 -216
rect 8631 -271 8714 -254
rect 8490 -288 8506 -271
rect 8440 -304 8506 -288
rect 8698 -288 8714 -271
rect 8748 -271 8831 -254
rect 8889 -254 9089 -216
rect 8889 -271 8972 -254
rect 8748 -288 8764 -271
rect 8698 -304 8764 -288
rect 8956 -288 8972 -271
rect 9006 -271 9089 -254
rect 9147 -254 9347 -216
rect 9147 -271 9230 -254
rect 9006 -288 9022 -271
rect 8956 -304 9022 -288
rect 9214 -288 9230 -271
rect 9264 -271 9347 -254
rect 9405 -254 9605 -216
rect 9405 -271 9488 -254
rect 9264 -288 9280 -271
rect 9214 -304 9280 -288
rect 9472 -288 9488 -271
rect 9522 -271 9605 -254
rect 9663 -254 9863 -216
rect 9663 -271 9746 -254
rect 9522 -288 9538 -271
rect 9472 -304 9538 -288
rect 9730 -288 9746 -271
rect 9780 -271 9863 -254
rect 10520 -253 10720 -215
rect 10520 -270 10603 -253
rect 9780 -288 9796 -271
rect 9730 -304 9796 -288
rect 10587 -287 10603 -270
rect 10637 -270 10720 -253
rect 10778 -253 10978 -215
rect 10778 -270 10861 -253
rect 10637 -287 10653 -270
rect 10587 -303 10653 -287
rect 10845 -287 10861 -270
rect 10895 -270 10978 -253
rect 11036 -253 11236 -215
rect 11036 -270 11119 -253
rect 10895 -287 10911 -270
rect 10845 -303 10911 -287
rect 11103 -287 11119 -270
rect 11153 -270 11236 -253
rect 11294 -253 11494 -215
rect 11294 -270 11377 -253
rect 11153 -287 11169 -270
rect 11103 -303 11169 -287
rect 11361 -287 11377 -270
rect 11411 -270 11494 -253
rect 11552 -253 11752 -215
rect 11552 -270 11635 -253
rect 11411 -287 11427 -270
rect 11361 -303 11427 -287
rect 11619 -287 11635 -270
rect 11669 -270 11752 -253
rect 11810 -253 12010 -215
rect 11810 -270 11893 -253
rect 11669 -287 11685 -270
rect 11619 -303 11685 -287
rect 11877 -287 11893 -270
rect 11927 -270 12010 -253
rect 12068 -253 12268 -215
rect 12068 -270 12151 -253
rect 11927 -287 11943 -270
rect 11877 -303 11943 -287
rect 12135 -287 12151 -270
rect 12185 -270 12268 -253
rect 12326 -253 12526 -215
rect 12326 -270 12409 -253
rect 12185 -287 12201 -270
rect 12135 -303 12201 -287
rect 12393 -287 12409 -270
rect 12443 -270 12526 -253
rect 12443 -287 12459 -270
rect 12393 -303 12459 -287
rect 5254 -362 5320 -346
rect 5254 -379 5270 -362
rect 5187 -396 5270 -379
rect 5304 -379 5320 -362
rect 5512 -362 5578 -346
rect 5512 -379 5528 -362
rect 5304 -396 5387 -379
rect 5187 -434 5387 -396
rect 5445 -396 5528 -379
rect 5562 -379 5578 -362
rect 5770 -362 5836 -346
rect 5770 -379 5786 -362
rect 5562 -396 5645 -379
rect 5445 -434 5645 -396
rect 5703 -396 5786 -379
rect 5820 -379 5836 -362
rect 6028 -362 6094 -346
rect 6028 -379 6044 -362
rect 5820 -396 5903 -379
rect 5703 -434 5903 -396
rect 5961 -396 6044 -379
rect 6078 -379 6094 -362
rect 6286 -362 6352 -346
rect 6286 -379 6302 -362
rect 6078 -396 6161 -379
rect 5961 -434 6161 -396
rect 6219 -396 6302 -379
rect 6336 -379 6352 -362
rect 6544 -362 6610 -346
rect 6544 -379 6560 -362
rect 6336 -396 6419 -379
rect 6219 -434 6419 -396
rect 6477 -396 6560 -379
rect 6594 -379 6610 -362
rect 6802 -362 6868 -346
rect 6802 -379 6818 -362
rect 6594 -396 6677 -379
rect 6477 -434 6677 -396
rect 6735 -396 6818 -379
rect 6852 -379 6868 -362
rect 7060 -362 7126 -346
rect 7060 -379 7076 -362
rect 6852 -396 6935 -379
rect 6735 -434 6935 -396
rect 6993 -396 7076 -379
rect 7110 -379 7126 -362
rect 7924 -362 7990 -346
rect 7924 -379 7940 -362
rect 7110 -396 7193 -379
rect 6993 -434 7193 -396
rect 7857 -396 7940 -379
rect 7974 -379 7990 -362
rect 8182 -362 8248 -346
rect 8182 -379 8198 -362
rect 7974 -396 8057 -379
rect 7857 -434 8057 -396
rect 8115 -396 8198 -379
rect 8232 -379 8248 -362
rect 8440 -362 8506 -346
rect 8440 -379 8456 -362
rect 8232 -396 8315 -379
rect 8115 -434 8315 -396
rect 8373 -396 8456 -379
rect 8490 -379 8506 -362
rect 8698 -362 8764 -346
rect 8698 -379 8714 -362
rect 8490 -396 8573 -379
rect 8373 -434 8573 -396
rect 8631 -396 8714 -379
rect 8748 -379 8764 -362
rect 8956 -362 9022 -346
rect 8956 -379 8972 -362
rect 8748 -396 8831 -379
rect 8631 -434 8831 -396
rect 8889 -396 8972 -379
rect 9006 -379 9022 -362
rect 9214 -362 9280 -346
rect 9214 -379 9230 -362
rect 9006 -396 9089 -379
rect 8889 -434 9089 -396
rect 9147 -396 9230 -379
rect 9264 -379 9280 -362
rect 9472 -362 9538 -346
rect 9472 -379 9488 -362
rect 9264 -396 9347 -379
rect 9147 -434 9347 -396
rect 9405 -396 9488 -379
rect 9522 -379 9538 -362
rect 9730 -362 9796 -346
rect 9730 -379 9746 -362
rect 9522 -396 9605 -379
rect 9405 -434 9605 -396
rect 9663 -396 9746 -379
rect 9780 -379 9796 -362
rect 10587 -361 10653 -345
rect 10587 -378 10603 -361
rect 9780 -396 9863 -379
rect 9663 -434 9863 -396
rect 10520 -395 10603 -378
rect 10637 -378 10653 -361
rect 10845 -361 10911 -345
rect 10845 -378 10861 -361
rect 10637 -395 10720 -378
rect 10520 -433 10720 -395
rect 10778 -395 10861 -378
rect 10895 -378 10911 -361
rect 11103 -361 11169 -345
rect 11103 -378 11119 -361
rect 10895 -395 10978 -378
rect 10778 -433 10978 -395
rect 11036 -395 11119 -378
rect 11153 -378 11169 -361
rect 11361 -361 11427 -345
rect 11361 -378 11377 -361
rect 11153 -395 11236 -378
rect 11036 -433 11236 -395
rect 11294 -395 11377 -378
rect 11411 -378 11427 -361
rect 11619 -361 11685 -345
rect 11619 -378 11635 -361
rect 11411 -395 11494 -378
rect 11294 -433 11494 -395
rect 11552 -395 11635 -378
rect 11669 -378 11685 -361
rect 11877 -361 11943 -345
rect 11877 -378 11893 -361
rect 11669 -395 11752 -378
rect 11552 -433 11752 -395
rect 11810 -395 11893 -378
rect 11927 -378 11943 -361
rect 12135 -361 12201 -345
rect 12135 -378 12151 -361
rect 11927 -395 12010 -378
rect 11810 -433 12010 -395
rect 12068 -395 12151 -378
rect 12185 -378 12201 -361
rect 12393 -361 12459 -345
rect 12393 -378 12409 -361
rect 12185 -395 12268 -378
rect 12068 -433 12268 -395
rect 12326 -395 12409 -378
rect 12443 -378 12459 -361
rect 12443 -395 12526 -378
rect 12326 -433 12526 -395
rect 5187 -672 5387 -634
rect 5187 -689 5270 -672
rect 5254 -706 5270 -689
rect 5304 -689 5387 -672
rect 5445 -672 5645 -634
rect 5445 -689 5528 -672
rect 5304 -706 5320 -689
rect 5254 -722 5320 -706
rect 5512 -706 5528 -689
rect 5562 -689 5645 -672
rect 5703 -672 5903 -634
rect 5703 -689 5786 -672
rect 5562 -706 5578 -689
rect 5512 -722 5578 -706
rect 5770 -706 5786 -689
rect 5820 -689 5903 -672
rect 5961 -672 6161 -634
rect 5961 -689 6044 -672
rect 5820 -706 5836 -689
rect 5770 -722 5836 -706
rect 6028 -706 6044 -689
rect 6078 -689 6161 -672
rect 6219 -672 6419 -634
rect 6219 -689 6302 -672
rect 6078 -706 6094 -689
rect 6028 -722 6094 -706
rect 6286 -706 6302 -689
rect 6336 -689 6419 -672
rect 6477 -672 6677 -634
rect 6477 -689 6560 -672
rect 6336 -706 6352 -689
rect 6286 -722 6352 -706
rect 6544 -706 6560 -689
rect 6594 -689 6677 -672
rect 6735 -672 6935 -634
rect 6735 -689 6818 -672
rect 6594 -706 6610 -689
rect 6544 -722 6610 -706
rect 6802 -706 6818 -689
rect 6852 -689 6935 -672
rect 6993 -672 7193 -634
rect 6993 -689 7076 -672
rect 6852 -706 6868 -689
rect 6802 -722 6868 -706
rect 7060 -706 7076 -689
rect 7110 -689 7193 -672
rect 7857 -672 8057 -634
rect 7857 -689 7940 -672
rect 7110 -706 7126 -689
rect 7060 -722 7126 -706
rect 7924 -706 7940 -689
rect 7974 -689 8057 -672
rect 8115 -672 8315 -634
rect 8115 -689 8198 -672
rect 7974 -706 7990 -689
rect 7924 -722 7990 -706
rect 8182 -706 8198 -689
rect 8232 -689 8315 -672
rect 8373 -672 8573 -634
rect 8373 -689 8456 -672
rect 8232 -706 8248 -689
rect 8182 -722 8248 -706
rect 8440 -706 8456 -689
rect 8490 -689 8573 -672
rect 8631 -672 8831 -634
rect 8631 -689 8714 -672
rect 8490 -706 8506 -689
rect 8440 -722 8506 -706
rect 8698 -706 8714 -689
rect 8748 -689 8831 -672
rect 8889 -672 9089 -634
rect 8889 -689 8972 -672
rect 8748 -706 8764 -689
rect 8698 -722 8764 -706
rect 8956 -706 8972 -689
rect 9006 -689 9089 -672
rect 9147 -672 9347 -634
rect 9147 -689 9230 -672
rect 9006 -706 9022 -689
rect 8956 -722 9022 -706
rect 9214 -706 9230 -689
rect 9264 -689 9347 -672
rect 9405 -672 9605 -634
rect 9405 -689 9488 -672
rect 9264 -706 9280 -689
rect 9214 -722 9280 -706
rect 9472 -706 9488 -689
rect 9522 -689 9605 -672
rect 9663 -672 9863 -634
rect 9663 -689 9746 -672
rect 9522 -706 9538 -689
rect 9472 -722 9538 -706
rect 9730 -706 9746 -689
rect 9780 -689 9863 -672
rect 10520 -671 10720 -633
rect 10520 -688 10603 -671
rect 9780 -706 9796 -689
rect 9730 -722 9796 -706
rect 10587 -705 10603 -688
rect 10637 -688 10720 -671
rect 10778 -671 10978 -633
rect 10778 -688 10861 -671
rect 10637 -705 10653 -688
rect 10587 -721 10653 -705
rect 10845 -705 10861 -688
rect 10895 -688 10978 -671
rect 11036 -671 11236 -633
rect 11036 -688 11119 -671
rect 10895 -705 10911 -688
rect 10845 -721 10911 -705
rect 11103 -705 11119 -688
rect 11153 -688 11236 -671
rect 11294 -671 11494 -633
rect 11294 -688 11377 -671
rect 11153 -705 11169 -688
rect 11103 -721 11169 -705
rect 11361 -705 11377 -688
rect 11411 -688 11494 -671
rect 11552 -671 11752 -633
rect 11552 -688 11635 -671
rect 11411 -705 11427 -688
rect 11361 -721 11427 -705
rect 11619 -705 11635 -688
rect 11669 -688 11752 -671
rect 11810 -671 12010 -633
rect 11810 -688 11893 -671
rect 11669 -705 11685 -688
rect 11619 -721 11685 -705
rect 11877 -705 11893 -688
rect 11927 -688 12010 -671
rect 12068 -671 12268 -633
rect 12068 -688 12151 -671
rect 11927 -705 11943 -688
rect 11877 -721 11943 -705
rect 12135 -705 12151 -688
rect 12185 -688 12268 -671
rect 12326 -671 12526 -633
rect 12326 -688 12409 -671
rect 12185 -705 12201 -688
rect 12135 -721 12201 -705
rect 12393 -705 12409 -688
rect 12443 -688 12526 -671
rect 12443 -705 12459 -688
rect 12393 -721 12459 -705
rect 5254 -780 5320 -764
rect 5254 -797 5270 -780
rect 5187 -814 5270 -797
rect 5304 -797 5320 -780
rect 5512 -780 5578 -764
rect 5512 -797 5528 -780
rect 5304 -814 5387 -797
rect 5187 -852 5387 -814
rect 5445 -814 5528 -797
rect 5562 -797 5578 -780
rect 5770 -780 5836 -764
rect 5770 -797 5786 -780
rect 5562 -814 5645 -797
rect 5445 -852 5645 -814
rect 5703 -814 5786 -797
rect 5820 -797 5836 -780
rect 6028 -780 6094 -764
rect 6028 -797 6044 -780
rect 5820 -814 5903 -797
rect 5703 -852 5903 -814
rect 5961 -814 6044 -797
rect 6078 -797 6094 -780
rect 6286 -780 6352 -764
rect 6286 -797 6302 -780
rect 6078 -814 6161 -797
rect 5961 -852 6161 -814
rect 6219 -814 6302 -797
rect 6336 -797 6352 -780
rect 6544 -780 6610 -764
rect 6544 -797 6560 -780
rect 6336 -814 6419 -797
rect 6219 -852 6419 -814
rect 6477 -814 6560 -797
rect 6594 -797 6610 -780
rect 6802 -780 6868 -764
rect 6802 -797 6818 -780
rect 6594 -814 6677 -797
rect 6477 -852 6677 -814
rect 6735 -814 6818 -797
rect 6852 -797 6868 -780
rect 7060 -780 7126 -764
rect 7060 -797 7076 -780
rect 6852 -814 6935 -797
rect 6735 -852 6935 -814
rect 6993 -814 7076 -797
rect 7110 -797 7126 -780
rect 7924 -780 7990 -764
rect 7924 -797 7940 -780
rect 7110 -814 7193 -797
rect 6993 -852 7193 -814
rect 7857 -814 7940 -797
rect 7974 -797 7990 -780
rect 8182 -780 8248 -764
rect 8182 -797 8198 -780
rect 7974 -814 8057 -797
rect 7857 -852 8057 -814
rect 8115 -814 8198 -797
rect 8232 -797 8248 -780
rect 8440 -780 8506 -764
rect 8440 -797 8456 -780
rect 8232 -814 8315 -797
rect 8115 -852 8315 -814
rect 8373 -814 8456 -797
rect 8490 -797 8506 -780
rect 8698 -780 8764 -764
rect 8698 -797 8714 -780
rect 8490 -814 8573 -797
rect 8373 -852 8573 -814
rect 8631 -814 8714 -797
rect 8748 -797 8764 -780
rect 8956 -780 9022 -764
rect 8956 -797 8972 -780
rect 8748 -814 8831 -797
rect 8631 -852 8831 -814
rect 8889 -814 8972 -797
rect 9006 -797 9022 -780
rect 9214 -780 9280 -764
rect 9214 -797 9230 -780
rect 9006 -814 9089 -797
rect 8889 -852 9089 -814
rect 9147 -814 9230 -797
rect 9264 -797 9280 -780
rect 9472 -780 9538 -764
rect 9472 -797 9488 -780
rect 9264 -814 9347 -797
rect 9147 -852 9347 -814
rect 9405 -814 9488 -797
rect 9522 -797 9538 -780
rect 9730 -780 9796 -764
rect 9730 -797 9746 -780
rect 9522 -814 9605 -797
rect 9405 -852 9605 -814
rect 9663 -814 9746 -797
rect 9780 -797 9796 -780
rect 10587 -779 10653 -763
rect 10587 -796 10603 -779
rect 9780 -814 9863 -797
rect 9663 -852 9863 -814
rect 10520 -813 10603 -796
rect 10637 -796 10653 -779
rect 10845 -779 10911 -763
rect 10845 -796 10861 -779
rect 10637 -813 10720 -796
rect 10520 -851 10720 -813
rect 10778 -813 10861 -796
rect 10895 -796 10911 -779
rect 11103 -779 11169 -763
rect 11103 -796 11119 -779
rect 10895 -813 10978 -796
rect 10778 -851 10978 -813
rect 11036 -813 11119 -796
rect 11153 -796 11169 -779
rect 11361 -779 11427 -763
rect 11361 -796 11377 -779
rect 11153 -813 11236 -796
rect 11036 -851 11236 -813
rect 11294 -813 11377 -796
rect 11411 -796 11427 -779
rect 11619 -779 11685 -763
rect 11619 -796 11635 -779
rect 11411 -813 11494 -796
rect 11294 -851 11494 -813
rect 11552 -813 11635 -796
rect 11669 -796 11685 -779
rect 11877 -779 11943 -763
rect 11877 -796 11893 -779
rect 11669 -813 11752 -796
rect 11552 -851 11752 -813
rect 11810 -813 11893 -796
rect 11927 -796 11943 -779
rect 12135 -779 12201 -763
rect 12135 -796 12151 -779
rect 11927 -813 12010 -796
rect 11810 -851 12010 -813
rect 12068 -813 12151 -796
rect 12185 -796 12201 -779
rect 12393 -779 12459 -763
rect 12393 -796 12409 -779
rect 12185 -813 12268 -796
rect 12068 -851 12268 -813
rect 12326 -813 12409 -796
rect 12443 -796 12459 -779
rect 12443 -813 12526 -796
rect 12326 -851 12526 -813
rect 5187 -1090 5387 -1052
rect 5187 -1107 5270 -1090
rect 5254 -1124 5270 -1107
rect 5304 -1107 5387 -1090
rect 5445 -1090 5645 -1052
rect 5445 -1107 5528 -1090
rect 5304 -1124 5320 -1107
rect 5254 -1140 5320 -1124
rect 5512 -1124 5528 -1107
rect 5562 -1107 5645 -1090
rect 5703 -1090 5903 -1052
rect 5703 -1107 5786 -1090
rect 5562 -1124 5578 -1107
rect 5512 -1140 5578 -1124
rect 5770 -1124 5786 -1107
rect 5820 -1107 5903 -1090
rect 5961 -1090 6161 -1052
rect 5961 -1107 6044 -1090
rect 5820 -1124 5836 -1107
rect 5770 -1140 5836 -1124
rect 6028 -1124 6044 -1107
rect 6078 -1107 6161 -1090
rect 6219 -1090 6419 -1052
rect 6219 -1107 6302 -1090
rect 6078 -1124 6094 -1107
rect 6028 -1140 6094 -1124
rect 6286 -1124 6302 -1107
rect 6336 -1107 6419 -1090
rect 6477 -1090 6677 -1052
rect 6477 -1107 6560 -1090
rect 6336 -1124 6352 -1107
rect 6286 -1140 6352 -1124
rect 6544 -1124 6560 -1107
rect 6594 -1107 6677 -1090
rect 6735 -1090 6935 -1052
rect 6735 -1107 6818 -1090
rect 6594 -1124 6610 -1107
rect 6544 -1140 6610 -1124
rect 6802 -1124 6818 -1107
rect 6852 -1107 6935 -1090
rect 6993 -1090 7193 -1052
rect 6993 -1107 7076 -1090
rect 6852 -1124 6868 -1107
rect 6802 -1140 6868 -1124
rect 7060 -1124 7076 -1107
rect 7110 -1107 7193 -1090
rect 7857 -1090 8057 -1052
rect 7857 -1107 7940 -1090
rect 7110 -1124 7126 -1107
rect 7060 -1140 7126 -1124
rect 7924 -1124 7940 -1107
rect 7974 -1107 8057 -1090
rect 8115 -1090 8315 -1052
rect 8115 -1107 8198 -1090
rect 7974 -1124 7990 -1107
rect 7924 -1140 7990 -1124
rect 8182 -1124 8198 -1107
rect 8232 -1107 8315 -1090
rect 8373 -1090 8573 -1052
rect 8373 -1107 8456 -1090
rect 8232 -1124 8248 -1107
rect 8182 -1140 8248 -1124
rect 8440 -1124 8456 -1107
rect 8490 -1107 8573 -1090
rect 8631 -1090 8831 -1052
rect 8631 -1107 8714 -1090
rect 8490 -1124 8506 -1107
rect 8440 -1140 8506 -1124
rect 8698 -1124 8714 -1107
rect 8748 -1107 8831 -1090
rect 8889 -1090 9089 -1052
rect 8889 -1107 8972 -1090
rect 8748 -1124 8764 -1107
rect 8698 -1140 8764 -1124
rect 8956 -1124 8972 -1107
rect 9006 -1107 9089 -1090
rect 9147 -1090 9347 -1052
rect 9147 -1107 9230 -1090
rect 9006 -1124 9022 -1107
rect 8956 -1140 9022 -1124
rect 9214 -1124 9230 -1107
rect 9264 -1107 9347 -1090
rect 9405 -1090 9605 -1052
rect 9405 -1107 9488 -1090
rect 9264 -1124 9280 -1107
rect 9214 -1140 9280 -1124
rect 9472 -1124 9488 -1107
rect 9522 -1107 9605 -1090
rect 9663 -1090 9863 -1052
rect 9663 -1107 9746 -1090
rect 9522 -1124 9538 -1107
rect 9472 -1140 9538 -1124
rect 9730 -1124 9746 -1107
rect 9780 -1107 9863 -1090
rect 10520 -1089 10720 -1051
rect 10520 -1106 10603 -1089
rect 9780 -1124 9796 -1107
rect 9730 -1140 9796 -1124
rect 10587 -1123 10603 -1106
rect 10637 -1106 10720 -1089
rect 10778 -1089 10978 -1051
rect 10778 -1106 10861 -1089
rect 10637 -1123 10653 -1106
rect 10587 -1139 10653 -1123
rect 10845 -1123 10861 -1106
rect 10895 -1106 10978 -1089
rect 11036 -1089 11236 -1051
rect 11036 -1106 11119 -1089
rect 10895 -1123 10911 -1106
rect 10845 -1139 10911 -1123
rect 11103 -1123 11119 -1106
rect 11153 -1106 11236 -1089
rect 11294 -1089 11494 -1051
rect 11294 -1106 11377 -1089
rect 11153 -1123 11169 -1106
rect 11103 -1139 11169 -1123
rect 11361 -1123 11377 -1106
rect 11411 -1106 11494 -1089
rect 11552 -1089 11752 -1051
rect 11552 -1106 11635 -1089
rect 11411 -1123 11427 -1106
rect 11361 -1139 11427 -1123
rect 11619 -1123 11635 -1106
rect 11669 -1106 11752 -1089
rect 11810 -1089 12010 -1051
rect 11810 -1106 11893 -1089
rect 11669 -1123 11685 -1106
rect 11619 -1139 11685 -1123
rect 11877 -1123 11893 -1106
rect 11927 -1106 12010 -1089
rect 12068 -1089 12268 -1051
rect 12068 -1106 12151 -1089
rect 11927 -1123 11943 -1106
rect 11877 -1139 11943 -1123
rect 12135 -1123 12151 -1106
rect 12185 -1106 12268 -1089
rect 12326 -1089 12526 -1051
rect 12326 -1106 12409 -1089
rect 12185 -1123 12201 -1106
rect 12135 -1139 12201 -1123
rect 12393 -1123 12409 -1106
rect 12443 -1106 12526 -1089
rect 12443 -1123 12459 -1106
rect 12393 -1139 12459 -1123
rect 5254 -1198 5320 -1182
rect 5254 -1215 5270 -1198
rect 5187 -1232 5270 -1215
rect 5304 -1215 5320 -1198
rect 5512 -1198 5578 -1182
rect 5512 -1215 5528 -1198
rect 5304 -1232 5387 -1215
rect 5187 -1270 5387 -1232
rect 5445 -1232 5528 -1215
rect 5562 -1215 5578 -1198
rect 5770 -1198 5836 -1182
rect 5770 -1215 5786 -1198
rect 5562 -1232 5645 -1215
rect 5445 -1270 5645 -1232
rect 5703 -1232 5786 -1215
rect 5820 -1215 5836 -1198
rect 6028 -1198 6094 -1182
rect 6028 -1215 6044 -1198
rect 5820 -1232 5903 -1215
rect 5703 -1270 5903 -1232
rect 5961 -1232 6044 -1215
rect 6078 -1215 6094 -1198
rect 6286 -1198 6352 -1182
rect 6286 -1215 6302 -1198
rect 6078 -1232 6161 -1215
rect 5961 -1270 6161 -1232
rect 6219 -1232 6302 -1215
rect 6336 -1215 6352 -1198
rect 6544 -1198 6610 -1182
rect 6544 -1215 6560 -1198
rect 6336 -1232 6419 -1215
rect 6219 -1270 6419 -1232
rect 6477 -1232 6560 -1215
rect 6594 -1215 6610 -1198
rect 6802 -1198 6868 -1182
rect 6802 -1215 6818 -1198
rect 6594 -1232 6677 -1215
rect 6477 -1270 6677 -1232
rect 6735 -1232 6818 -1215
rect 6852 -1215 6868 -1198
rect 7060 -1198 7126 -1182
rect 7060 -1215 7076 -1198
rect 6852 -1232 6935 -1215
rect 6735 -1270 6935 -1232
rect 6993 -1232 7076 -1215
rect 7110 -1215 7126 -1198
rect 7924 -1198 7990 -1182
rect 7924 -1215 7940 -1198
rect 7110 -1232 7193 -1215
rect 6993 -1270 7193 -1232
rect 7857 -1232 7940 -1215
rect 7974 -1215 7990 -1198
rect 8182 -1198 8248 -1182
rect 8182 -1215 8198 -1198
rect 7974 -1232 8057 -1215
rect 7857 -1270 8057 -1232
rect 8115 -1232 8198 -1215
rect 8232 -1215 8248 -1198
rect 8440 -1198 8506 -1182
rect 8440 -1215 8456 -1198
rect 8232 -1232 8315 -1215
rect 8115 -1270 8315 -1232
rect 8373 -1232 8456 -1215
rect 8490 -1215 8506 -1198
rect 8698 -1198 8764 -1182
rect 8698 -1215 8714 -1198
rect 8490 -1232 8573 -1215
rect 8373 -1270 8573 -1232
rect 8631 -1232 8714 -1215
rect 8748 -1215 8764 -1198
rect 8956 -1198 9022 -1182
rect 8956 -1215 8972 -1198
rect 8748 -1232 8831 -1215
rect 8631 -1270 8831 -1232
rect 8889 -1232 8972 -1215
rect 9006 -1215 9022 -1198
rect 9214 -1198 9280 -1182
rect 9214 -1215 9230 -1198
rect 9006 -1232 9089 -1215
rect 8889 -1270 9089 -1232
rect 9147 -1232 9230 -1215
rect 9264 -1215 9280 -1198
rect 9472 -1198 9538 -1182
rect 9472 -1215 9488 -1198
rect 9264 -1232 9347 -1215
rect 9147 -1270 9347 -1232
rect 9405 -1232 9488 -1215
rect 9522 -1215 9538 -1198
rect 9730 -1198 9796 -1182
rect 9730 -1215 9746 -1198
rect 9522 -1232 9605 -1215
rect 9405 -1270 9605 -1232
rect 9663 -1232 9746 -1215
rect 9780 -1215 9796 -1198
rect 10587 -1197 10653 -1181
rect 10587 -1214 10603 -1197
rect 9780 -1232 9863 -1215
rect 9663 -1270 9863 -1232
rect 10520 -1231 10603 -1214
rect 10637 -1214 10653 -1197
rect 10845 -1197 10911 -1181
rect 10845 -1214 10861 -1197
rect 10637 -1231 10720 -1214
rect 10520 -1269 10720 -1231
rect 10778 -1231 10861 -1214
rect 10895 -1214 10911 -1197
rect 11103 -1197 11169 -1181
rect 11103 -1214 11119 -1197
rect 10895 -1231 10978 -1214
rect 10778 -1269 10978 -1231
rect 11036 -1231 11119 -1214
rect 11153 -1214 11169 -1197
rect 11361 -1197 11427 -1181
rect 11361 -1214 11377 -1197
rect 11153 -1231 11236 -1214
rect 11036 -1269 11236 -1231
rect 11294 -1231 11377 -1214
rect 11411 -1214 11427 -1197
rect 11619 -1197 11685 -1181
rect 11619 -1214 11635 -1197
rect 11411 -1231 11494 -1214
rect 11294 -1269 11494 -1231
rect 11552 -1231 11635 -1214
rect 11669 -1214 11685 -1197
rect 11877 -1197 11943 -1181
rect 11877 -1214 11893 -1197
rect 11669 -1231 11752 -1214
rect 11552 -1269 11752 -1231
rect 11810 -1231 11893 -1214
rect 11927 -1214 11943 -1197
rect 12135 -1197 12201 -1181
rect 12135 -1214 12151 -1197
rect 11927 -1231 12010 -1214
rect 11810 -1269 12010 -1231
rect 12068 -1231 12151 -1214
rect 12185 -1214 12201 -1197
rect 12393 -1197 12459 -1181
rect 12393 -1214 12409 -1197
rect 12185 -1231 12268 -1214
rect 12068 -1269 12268 -1231
rect 12326 -1231 12409 -1214
rect 12443 -1214 12459 -1197
rect 12443 -1231 12526 -1214
rect 12326 -1269 12526 -1231
rect 5187 -1508 5387 -1470
rect 5187 -1525 5270 -1508
rect 5254 -1542 5270 -1525
rect 5304 -1525 5387 -1508
rect 5445 -1508 5645 -1470
rect 5445 -1525 5528 -1508
rect 5304 -1542 5320 -1525
rect 5254 -1558 5320 -1542
rect 5512 -1542 5528 -1525
rect 5562 -1525 5645 -1508
rect 5703 -1508 5903 -1470
rect 5703 -1525 5786 -1508
rect 5562 -1542 5578 -1525
rect 5512 -1558 5578 -1542
rect 5770 -1542 5786 -1525
rect 5820 -1525 5903 -1508
rect 5961 -1508 6161 -1470
rect 5961 -1525 6044 -1508
rect 5820 -1542 5836 -1525
rect 5770 -1558 5836 -1542
rect 6028 -1542 6044 -1525
rect 6078 -1525 6161 -1508
rect 6219 -1508 6419 -1470
rect 6219 -1525 6302 -1508
rect 6078 -1542 6094 -1525
rect 6028 -1558 6094 -1542
rect 6286 -1542 6302 -1525
rect 6336 -1525 6419 -1508
rect 6477 -1508 6677 -1470
rect 6477 -1525 6560 -1508
rect 6336 -1542 6352 -1525
rect 6286 -1558 6352 -1542
rect 6544 -1542 6560 -1525
rect 6594 -1525 6677 -1508
rect 6735 -1508 6935 -1470
rect 6735 -1525 6818 -1508
rect 6594 -1542 6610 -1525
rect 6544 -1558 6610 -1542
rect 6802 -1542 6818 -1525
rect 6852 -1525 6935 -1508
rect 6993 -1508 7193 -1470
rect 6993 -1525 7076 -1508
rect 6852 -1542 6868 -1525
rect 6802 -1558 6868 -1542
rect 7060 -1542 7076 -1525
rect 7110 -1525 7193 -1508
rect 7857 -1508 8057 -1470
rect 7857 -1525 7940 -1508
rect 7110 -1542 7126 -1525
rect 7060 -1558 7126 -1542
rect 7924 -1542 7940 -1525
rect 7974 -1525 8057 -1508
rect 8115 -1508 8315 -1470
rect 8115 -1525 8198 -1508
rect 7974 -1542 7990 -1525
rect 7924 -1558 7990 -1542
rect 8182 -1542 8198 -1525
rect 8232 -1525 8315 -1508
rect 8373 -1508 8573 -1470
rect 8373 -1525 8456 -1508
rect 8232 -1542 8248 -1525
rect 8182 -1558 8248 -1542
rect 8440 -1542 8456 -1525
rect 8490 -1525 8573 -1508
rect 8631 -1508 8831 -1470
rect 8631 -1525 8714 -1508
rect 8490 -1542 8506 -1525
rect 8440 -1558 8506 -1542
rect 8698 -1542 8714 -1525
rect 8748 -1525 8831 -1508
rect 8889 -1508 9089 -1470
rect 8889 -1525 8972 -1508
rect 8748 -1542 8764 -1525
rect 8698 -1558 8764 -1542
rect 8956 -1542 8972 -1525
rect 9006 -1525 9089 -1508
rect 9147 -1508 9347 -1470
rect 9147 -1525 9230 -1508
rect 9006 -1542 9022 -1525
rect 8956 -1558 9022 -1542
rect 9214 -1542 9230 -1525
rect 9264 -1525 9347 -1508
rect 9405 -1508 9605 -1470
rect 9405 -1525 9488 -1508
rect 9264 -1542 9280 -1525
rect 9214 -1558 9280 -1542
rect 9472 -1542 9488 -1525
rect 9522 -1525 9605 -1508
rect 9663 -1508 9863 -1470
rect 9663 -1525 9746 -1508
rect 9522 -1542 9538 -1525
rect 9472 -1558 9538 -1542
rect 9730 -1542 9746 -1525
rect 9780 -1525 9863 -1508
rect 10520 -1507 10720 -1469
rect 10520 -1524 10603 -1507
rect 9780 -1542 9796 -1525
rect 9730 -1558 9796 -1542
rect 10587 -1541 10603 -1524
rect 10637 -1524 10720 -1507
rect 10778 -1507 10978 -1469
rect 10778 -1524 10861 -1507
rect 10637 -1541 10653 -1524
rect 10587 -1557 10653 -1541
rect 10845 -1541 10861 -1524
rect 10895 -1524 10978 -1507
rect 11036 -1507 11236 -1469
rect 11036 -1524 11119 -1507
rect 10895 -1541 10911 -1524
rect 10845 -1557 10911 -1541
rect 11103 -1541 11119 -1524
rect 11153 -1524 11236 -1507
rect 11294 -1507 11494 -1469
rect 11294 -1524 11377 -1507
rect 11153 -1541 11169 -1524
rect 11103 -1557 11169 -1541
rect 11361 -1541 11377 -1524
rect 11411 -1524 11494 -1507
rect 11552 -1507 11752 -1469
rect 11552 -1524 11635 -1507
rect 11411 -1541 11427 -1524
rect 11361 -1557 11427 -1541
rect 11619 -1541 11635 -1524
rect 11669 -1524 11752 -1507
rect 11810 -1507 12010 -1469
rect 11810 -1524 11893 -1507
rect 11669 -1541 11685 -1524
rect 11619 -1557 11685 -1541
rect 11877 -1541 11893 -1524
rect 11927 -1524 12010 -1507
rect 12068 -1507 12268 -1469
rect 12068 -1524 12151 -1507
rect 11927 -1541 11943 -1524
rect 11877 -1557 11943 -1541
rect 12135 -1541 12151 -1524
rect 12185 -1524 12268 -1507
rect 12326 -1507 12526 -1469
rect 12326 -1524 12409 -1507
rect 12185 -1541 12201 -1524
rect 12135 -1557 12201 -1541
rect 12393 -1541 12409 -1524
rect 12443 -1524 12526 -1507
rect 12443 -1541 12459 -1524
rect 12393 -1557 12459 -1541
rect 5254 -1616 5320 -1600
rect 5254 -1633 5270 -1616
rect 5187 -1650 5270 -1633
rect 5304 -1633 5320 -1616
rect 5512 -1616 5578 -1600
rect 5512 -1633 5528 -1616
rect 5304 -1650 5387 -1633
rect 5187 -1688 5387 -1650
rect 5445 -1650 5528 -1633
rect 5562 -1633 5578 -1616
rect 5770 -1616 5836 -1600
rect 5770 -1633 5786 -1616
rect 5562 -1650 5645 -1633
rect 5445 -1688 5645 -1650
rect 5703 -1650 5786 -1633
rect 5820 -1633 5836 -1616
rect 6028 -1616 6094 -1600
rect 6028 -1633 6044 -1616
rect 5820 -1650 5903 -1633
rect 5703 -1688 5903 -1650
rect 5961 -1650 6044 -1633
rect 6078 -1633 6094 -1616
rect 6286 -1616 6352 -1600
rect 6286 -1633 6302 -1616
rect 6078 -1650 6161 -1633
rect 5961 -1688 6161 -1650
rect 6219 -1650 6302 -1633
rect 6336 -1633 6352 -1616
rect 6544 -1616 6610 -1600
rect 6544 -1633 6560 -1616
rect 6336 -1650 6419 -1633
rect 6219 -1688 6419 -1650
rect 6477 -1650 6560 -1633
rect 6594 -1633 6610 -1616
rect 6802 -1616 6868 -1600
rect 6802 -1633 6818 -1616
rect 6594 -1650 6677 -1633
rect 6477 -1688 6677 -1650
rect 6735 -1650 6818 -1633
rect 6852 -1633 6868 -1616
rect 7060 -1616 7126 -1600
rect 7060 -1633 7076 -1616
rect 6852 -1650 6935 -1633
rect 6735 -1688 6935 -1650
rect 6993 -1650 7076 -1633
rect 7110 -1633 7126 -1616
rect 7924 -1616 7990 -1600
rect 7924 -1633 7940 -1616
rect 7110 -1650 7193 -1633
rect 6993 -1688 7193 -1650
rect 7857 -1650 7940 -1633
rect 7974 -1633 7990 -1616
rect 8182 -1616 8248 -1600
rect 8182 -1633 8198 -1616
rect 7974 -1650 8057 -1633
rect 7857 -1688 8057 -1650
rect 8115 -1650 8198 -1633
rect 8232 -1633 8248 -1616
rect 8440 -1616 8506 -1600
rect 8440 -1633 8456 -1616
rect 8232 -1650 8315 -1633
rect 8115 -1688 8315 -1650
rect 8373 -1650 8456 -1633
rect 8490 -1633 8506 -1616
rect 8698 -1616 8764 -1600
rect 8698 -1633 8714 -1616
rect 8490 -1650 8573 -1633
rect 8373 -1688 8573 -1650
rect 8631 -1650 8714 -1633
rect 8748 -1633 8764 -1616
rect 8956 -1616 9022 -1600
rect 8956 -1633 8972 -1616
rect 8748 -1650 8831 -1633
rect 8631 -1688 8831 -1650
rect 8889 -1650 8972 -1633
rect 9006 -1633 9022 -1616
rect 9214 -1616 9280 -1600
rect 9214 -1633 9230 -1616
rect 9006 -1650 9089 -1633
rect 8889 -1688 9089 -1650
rect 9147 -1650 9230 -1633
rect 9264 -1633 9280 -1616
rect 9472 -1616 9538 -1600
rect 9472 -1633 9488 -1616
rect 9264 -1650 9347 -1633
rect 9147 -1688 9347 -1650
rect 9405 -1650 9488 -1633
rect 9522 -1633 9538 -1616
rect 9730 -1616 9796 -1600
rect 9730 -1633 9746 -1616
rect 9522 -1650 9605 -1633
rect 9405 -1688 9605 -1650
rect 9663 -1650 9746 -1633
rect 9780 -1633 9796 -1616
rect 10587 -1615 10653 -1599
rect 10587 -1632 10603 -1615
rect 9780 -1650 9863 -1633
rect 9663 -1688 9863 -1650
rect 10520 -1649 10603 -1632
rect 10637 -1632 10653 -1615
rect 10845 -1615 10911 -1599
rect 10845 -1632 10861 -1615
rect 10637 -1649 10720 -1632
rect 10520 -1687 10720 -1649
rect 10778 -1649 10861 -1632
rect 10895 -1632 10911 -1615
rect 11103 -1615 11169 -1599
rect 11103 -1632 11119 -1615
rect 10895 -1649 10978 -1632
rect 10778 -1687 10978 -1649
rect 11036 -1649 11119 -1632
rect 11153 -1632 11169 -1615
rect 11361 -1615 11427 -1599
rect 11361 -1632 11377 -1615
rect 11153 -1649 11236 -1632
rect 11036 -1687 11236 -1649
rect 11294 -1649 11377 -1632
rect 11411 -1632 11427 -1615
rect 11619 -1615 11685 -1599
rect 11619 -1632 11635 -1615
rect 11411 -1649 11494 -1632
rect 11294 -1687 11494 -1649
rect 11552 -1649 11635 -1632
rect 11669 -1632 11685 -1615
rect 11877 -1615 11943 -1599
rect 11877 -1632 11893 -1615
rect 11669 -1649 11752 -1632
rect 11552 -1687 11752 -1649
rect 11810 -1649 11893 -1632
rect 11927 -1632 11943 -1615
rect 12135 -1615 12201 -1599
rect 12135 -1632 12151 -1615
rect 11927 -1649 12010 -1632
rect 11810 -1687 12010 -1649
rect 12068 -1649 12151 -1632
rect 12185 -1632 12201 -1615
rect 12393 -1615 12459 -1599
rect 12393 -1632 12409 -1615
rect 12185 -1649 12268 -1632
rect 12068 -1687 12268 -1649
rect 12326 -1649 12409 -1632
rect 12443 -1632 12459 -1615
rect 12443 -1649 12526 -1632
rect 12326 -1687 12526 -1649
rect 5187 -1926 5387 -1888
rect 5187 -1943 5270 -1926
rect 5254 -1960 5270 -1943
rect 5304 -1943 5387 -1926
rect 5445 -1926 5645 -1888
rect 5445 -1943 5528 -1926
rect 5304 -1960 5320 -1943
rect 5254 -1976 5320 -1960
rect 5512 -1960 5528 -1943
rect 5562 -1943 5645 -1926
rect 5703 -1926 5903 -1888
rect 5703 -1943 5786 -1926
rect 5562 -1960 5578 -1943
rect 5512 -1976 5578 -1960
rect 5770 -1960 5786 -1943
rect 5820 -1943 5903 -1926
rect 5961 -1926 6161 -1888
rect 5961 -1943 6044 -1926
rect 5820 -1960 5836 -1943
rect 5770 -1976 5836 -1960
rect 6028 -1960 6044 -1943
rect 6078 -1943 6161 -1926
rect 6219 -1926 6419 -1888
rect 6219 -1943 6302 -1926
rect 6078 -1960 6094 -1943
rect 6028 -1976 6094 -1960
rect 6286 -1960 6302 -1943
rect 6336 -1943 6419 -1926
rect 6477 -1926 6677 -1888
rect 6477 -1943 6560 -1926
rect 6336 -1960 6352 -1943
rect 6286 -1976 6352 -1960
rect 6544 -1960 6560 -1943
rect 6594 -1943 6677 -1926
rect 6735 -1926 6935 -1888
rect 6735 -1943 6818 -1926
rect 6594 -1960 6610 -1943
rect 6544 -1976 6610 -1960
rect 6802 -1960 6818 -1943
rect 6852 -1943 6935 -1926
rect 6993 -1926 7193 -1888
rect 6993 -1943 7076 -1926
rect 6852 -1960 6868 -1943
rect 6802 -1976 6868 -1960
rect 7060 -1960 7076 -1943
rect 7110 -1943 7193 -1926
rect 7857 -1926 8057 -1888
rect 7857 -1943 7940 -1926
rect 7110 -1960 7126 -1943
rect 7060 -1976 7126 -1960
rect 7924 -1960 7940 -1943
rect 7974 -1943 8057 -1926
rect 8115 -1926 8315 -1888
rect 8115 -1943 8198 -1926
rect 7974 -1960 7990 -1943
rect 7924 -1976 7990 -1960
rect 8182 -1960 8198 -1943
rect 8232 -1943 8315 -1926
rect 8373 -1926 8573 -1888
rect 8373 -1943 8456 -1926
rect 8232 -1960 8248 -1943
rect 8182 -1976 8248 -1960
rect 8440 -1960 8456 -1943
rect 8490 -1943 8573 -1926
rect 8631 -1926 8831 -1888
rect 8631 -1943 8714 -1926
rect 8490 -1960 8506 -1943
rect 8440 -1976 8506 -1960
rect 8698 -1960 8714 -1943
rect 8748 -1943 8831 -1926
rect 8889 -1926 9089 -1888
rect 8889 -1943 8972 -1926
rect 8748 -1960 8764 -1943
rect 8698 -1976 8764 -1960
rect 8956 -1960 8972 -1943
rect 9006 -1943 9089 -1926
rect 9147 -1926 9347 -1888
rect 9147 -1943 9230 -1926
rect 9006 -1960 9022 -1943
rect 8956 -1976 9022 -1960
rect 9214 -1960 9230 -1943
rect 9264 -1943 9347 -1926
rect 9405 -1926 9605 -1888
rect 9405 -1943 9488 -1926
rect 9264 -1960 9280 -1943
rect 9214 -1976 9280 -1960
rect 9472 -1960 9488 -1943
rect 9522 -1943 9605 -1926
rect 9663 -1926 9863 -1888
rect 9663 -1943 9746 -1926
rect 9522 -1960 9538 -1943
rect 9472 -1976 9538 -1960
rect 9730 -1960 9746 -1943
rect 9780 -1943 9863 -1926
rect 10520 -1925 10720 -1887
rect 10520 -1942 10603 -1925
rect 9780 -1960 9796 -1943
rect 9730 -1976 9796 -1960
rect 10587 -1959 10603 -1942
rect 10637 -1942 10720 -1925
rect 10778 -1925 10978 -1887
rect 10778 -1942 10861 -1925
rect 10637 -1959 10653 -1942
rect 10587 -1975 10653 -1959
rect 10845 -1959 10861 -1942
rect 10895 -1942 10978 -1925
rect 11036 -1925 11236 -1887
rect 11036 -1942 11119 -1925
rect 10895 -1959 10911 -1942
rect 10845 -1975 10911 -1959
rect 11103 -1959 11119 -1942
rect 11153 -1942 11236 -1925
rect 11294 -1925 11494 -1887
rect 11294 -1942 11377 -1925
rect 11153 -1959 11169 -1942
rect 11103 -1975 11169 -1959
rect 11361 -1959 11377 -1942
rect 11411 -1942 11494 -1925
rect 11552 -1925 11752 -1887
rect 11552 -1942 11635 -1925
rect 11411 -1959 11427 -1942
rect 11361 -1975 11427 -1959
rect 11619 -1959 11635 -1942
rect 11669 -1942 11752 -1925
rect 11810 -1925 12010 -1887
rect 11810 -1942 11893 -1925
rect 11669 -1959 11685 -1942
rect 11619 -1975 11685 -1959
rect 11877 -1959 11893 -1942
rect 11927 -1942 12010 -1925
rect 12068 -1925 12268 -1887
rect 12068 -1942 12151 -1925
rect 11927 -1959 11943 -1942
rect 11877 -1975 11943 -1959
rect 12135 -1959 12151 -1942
rect 12185 -1942 12268 -1925
rect 12326 -1925 12526 -1887
rect 12326 -1942 12409 -1925
rect 12185 -1959 12201 -1942
rect 12135 -1975 12201 -1959
rect 12393 -1959 12409 -1942
rect 12443 -1942 12526 -1925
rect 12443 -1959 12459 -1942
rect 12393 -1975 12459 -1959
rect 5134 -2268 5200 -2252
rect 5134 -2285 5150 -2268
rect 5067 -2302 5150 -2285
rect 5184 -2285 5200 -2268
rect 5674 -2268 5740 -2252
rect 5674 -2285 5690 -2268
rect 5184 -2302 5267 -2285
rect 5067 -2340 5267 -2302
rect 5607 -2302 5690 -2285
rect 5724 -2285 5740 -2268
rect 6154 -2268 6220 -2252
rect 6154 -2285 6170 -2268
rect 5724 -2302 5807 -2285
rect 5607 -2340 5807 -2302
rect 6087 -2302 6170 -2285
rect 6204 -2285 6220 -2268
rect 6657 -2266 6723 -2250
rect 6657 -2283 6673 -2266
rect 6204 -2302 6287 -2285
rect 6087 -2340 6287 -2302
rect 6590 -2300 6673 -2283
rect 6707 -2283 6723 -2266
rect 7167 -2256 7233 -2240
rect 7167 -2273 7183 -2256
rect 6707 -2300 6790 -2283
rect 6590 -2338 6790 -2300
rect 7100 -2290 7183 -2273
rect 7217 -2273 7233 -2256
rect 7804 -2268 7870 -2252
rect 7217 -2290 7300 -2273
rect 7804 -2285 7820 -2268
rect 7100 -2328 7300 -2290
rect 7737 -2302 7820 -2285
rect 7854 -2285 7870 -2268
rect 8344 -2268 8410 -2252
rect 8344 -2285 8360 -2268
rect 7854 -2302 7937 -2285
rect 7737 -2340 7937 -2302
rect 8277 -2302 8360 -2285
rect 8394 -2285 8410 -2268
rect 8824 -2268 8890 -2252
rect 8824 -2285 8840 -2268
rect 8394 -2302 8477 -2285
rect 8277 -2340 8477 -2302
rect 8757 -2302 8840 -2285
rect 8874 -2285 8890 -2268
rect 9327 -2266 9393 -2250
rect 9327 -2283 9343 -2266
rect 8874 -2302 8957 -2285
rect 8757 -2340 8957 -2302
rect 9260 -2300 9343 -2283
rect 9377 -2283 9393 -2266
rect 9837 -2256 9903 -2240
rect 9837 -2273 9853 -2256
rect 9377 -2300 9460 -2283
rect 9260 -2338 9460 -2300
rect 9770 -2290 9853 -2273
rect 9887 -2273 9903 -2256
rect 10467 -2267 10533 -2251
rect 9887 -2290 9970 -2273
rect 10467 -2284 10483 -2267
rect 9770 -2328 9970 -2290
rect 10400 -2301 10483 -2284
rect 10517 -2284 10533 -2267
rect 11007 -2267 11073 -2251
rect 11007 -2284 11023 -2267
rect 10517 -2301 10600 -2284
rect 5067 -2578 5267 -2540
rect 5067 -2595 5150 -2578
rect 5134 -2612 5150 -2595
rect 5184 -2595 5267 -2578
rect 5607 -2578 5807 -2540
rect 5607 -2595 5690 -2578
rect 5184 -2612 5200 -2595
rect 5134 -2628 5200 -2612
rect 5674 -2612 5690 -2595
rect 5724 -2595 5807 -2578
rect 6087 -2578 6287 -2540
rect 6087 -2595 6170 -2578
rect 5724 -2612 5740 -2595
rect 5674 -2628 5740 -2612
rect 6154 -2612 6170 -2595
rect 6204 -2595 6287 -2578
rect 6590 -2576 6790 -2538
rect 6590 -2593 6673 -2576
rect 6204 -2612 6220 -2595
rect 6154 -2628 6220 -2612
rect 6657 -2610 6673 -2593
rect 6707 -2593 6790 -2576
rect 7100 -2566 7300 -2528
rect 10400 -2339 10600 -2301
rect 10940 -2301 11023 -2284
rect 11057 -2284 11073 -2267
rect 11487 -2267 11553 -2251
rect 11487 -2284 11503 -2267
rect 11057 -2301 11140 -2284
rect 10940 -2339 11140 -2301
rect 11420 -2301 11503 -2284
rect 11537 -2284 11553 -2267
rect 11990 -2265 12056 -2249
rect 11990 -2282 12006 -2265
rect 11537 -2301 11620 -2284
rect 11420 -2339 11620 -2301
rect 11923 -2299 12006 -2282
rect 12040 -2282 12056 -2265
rect 12500 -2255 12566 -2239
rect 12500 -2272 12516 -2255
rect 12040 -2299 12123 -2282
rect 11923 -2337 12123 -2299
rect 12433 -2289 12516 -2272
rect 12550 -2272 12566 -2255
rect 12550 -2289 12633 -2272
rect 12433 -2327 12633 -2289
rect 7100 -2583 7183 -2566
rect 6707 -2610 6723 -2593
rect 6657 -2626 6723 -2610
rect 7167 -2600 7183 -2583
rect 7217 -2583 7300 -2566
rect 7737 -2578 7937 -2540
rect 7217 -2600 7233 -2583
rect 7737 -2595 7820 -2578
rect 7167 -2616 7233 -2600
rect 7804 -2612 7820 -2595
rect 7854 -2595 7937 -2578
rect 8277 -2578 8477 -2540
rect 8277 -2595 8360 -2578
rect 7854 -2612 7870 -2595
rect 7804 -2628 7870 -2612
rect 8344 -2612 8360 -2595
rect 8394 -2595 8477 -2578
rect 8757 -2578 8957 -2540
rect 8757 -2595 8840 -2578
rect 8394 -2612 8410 -2595
rect 8344 -2628 8410 -2612
rect 8824 -2612 8840 -2595
rect 8874 -2595 8957 -2578
rect 9260 -2576 9460 -2538
rect 9260 -2593 9343 -2576
rect 8874 -2612 8890 -2595
rect 8824 -2628 8890 -2612
rect 9327 -2610 9343 -2593
rect 9377 -2593 9460 -2576
rect 9770 -2566 9970 -2528
rect 9770 -2583 9853 -2566
rect 9377 -2610 9393 -2593
rect 9327 -2626 9393 -2610
rect 9837 -2600 9853 -2583
rect 9887 -2583 9970 -2566
rect 10400 -2577 10600 -2539
rect 9887 -2600 9903 -2583
rect 10400 -2594 10483 -2577
rect 9837 -2616 9903 -2600
rect 10467 -2611 10483 -2594
rect 10517 -2594 10600 -2577
rect 10940 -2577 11140 -2539
rect 10940 -2594 11023 -2577
rect 10517 -2611 10533 -2594
rect 10467 -2627 10533 -2611
rect 11007 -2611 11023 -2594
rect 11057 -2594 11140 -2577
rect 11420 -2577 11620 -2539
rect 11420 -2594 11503 -2577
rect 11057 -2611 11073 -2594
rect 11007 -2627 11073 -2611
rect 11487 -2611 11503 -2594
rect 11537 -2594 11620 -2577
rect 11923 -2575 12123 -2537
rect 11923 -2592 12006 -2575
rect 11537 -2611 11553 -2594
rect 11487 -2627 11553 -2611
rect 11990 -2609 12006 -2592
rect 12040 -2592 12123 -2575
rect 12433 -2565 12633 -2527
rect 12433 -2582 12516 -2565
rect 12040 -2609 12056 -2592
rect 11990 -2625 12056 -2609
rect 12500 -2599 12516 -2582
rect 12550 -2582 12633 -2565
rect 12550 -2599 12566 -2582
rect 12500 -2615 12566 -2599
rect 12710 -3368 12776 -3352
rect 12710 -3402 12726 -3368
rect 12760 -3402 12776 -3368
rect 12710 -3418 12776 -3402
rect 12728 -3449 12758 -3418
rect 5457 -3994 5573 -3966
rect 5457 -4032 5481 -3994
rect 5547 -4032 5573 -3994
rect 6072 -4002 6258 -3986
rect 6072 -4019 6088 -4002
rect 5457 -4082 5573 -4032
rect 5765 -4036 6088 -4019
rect 6242 -4019 6258 -4002
rect 6798 -3996 6914 -3968
rect 6242 -4036 6565 -4019
rect 5765 -4083 6565 -4036
rect 6798 -4034 6822 -3996
rect 6888 -4034 6914 -3996
rect 5457 -4256 5573 -4192
rect 6798 -4084 6914 -4034
rect 7168 -3996 7284 -3968
rect 7168 -4034 7192 -3996
rect 7258 -4034 7284 -3996
rect 7168 -4084 7284 -4034
rect 7590 -3996 7706 -3968
rect 7590 -4034 7614 -3996
rect 7680 -4034 7706 -3996
rect 7590 -4084 7706 -4034
rect 8012 -3996 8128 -3968
rect 8012 -4034 8036 -3996
rect 8102 -4034 8128 -3996
rect 8742 -4002 8928 -3986
rect 8742 -4019 8758 -4002
rect 8012 -4084 8128 -4034
rect 8435 -4036 8758 -4019
rect 8912 -4019 8928 -4002
rect 9499 -3996 9615 -3968
rect 8912 -4036 9235 -4019
rect 8435 -4083 9235 -4036
rect 9499 -4034 9523 -3996
rect 9589 -4034 9615 -3996
rect 5765 -4240 6565 -4193
rect 9499 -4084 9615 -4034
rect 9869 -3996 9985 -3968
rect 9869 -4034 9893 -3996
rect 9959 -4034 9985 -3996
rect 9869 -4084 9985 -4034
rect 10291 -3996 10407 -3968
rect 10291 -4034 10315 -3996
rect 10381 -4034 10407 -3996
rect 10291 -4084 10407 -4034
rect 10713 -3996 10829 -3968
rect 10713 -4034 10737 -3996
rect 10803 -4034 10829 -3996
rect 11405 -4001 11591 -3985
rect 11405 -4018 11421 -4001
rect 10713 -4084 10829 -4034
rect 11098 -4035 11421 -4018
rect 11575 -4018 11591 -4001
rect 11575 -4035 11898 -4018
rect 11098 -4082 11898 -4035
rect 5765 -4257 6088 -4240
rect 6072 -4274 6088 -4257
rect 6242 -4257 6565 -4240
rect 6242 -4274 6258 -4257
rect 6798 -4258 6914 -4194
rect 7168 -4258 7284 -4194
rect 7590 -4258 7706 -4194
rect 8012 -4258 8128 -4194
rect 8435 -4240 9235 -4193
rect 8435 -4257 8758 -4240
rect 6072 -4290 6258 -4274
rect 8742 -4274 8758 -4257
rect 8912 -4257 9235 -4240
rect 8912 -4274 8928 -4257
rect 9499 -4258 9615 -4194
rect 9869 -4258 9985 -4194
rect 10291 -4258 10407 -4194
rect 10713 -4258 10829 -4194
rect 11098 -4239 11898 -4192
rect 11098 -4256 11421 -4239
rect 8742 -4290 8928 -4274
rect 11405 -4273 11421 -4256
rect 11575 -4256 11898 -4239
rect 11575 -4273 11591 -4256
rect 11405 -4289 11591 -4273
rect 13100 -3370 13166 -3354
rect 13100 -3404 13116 -3370
rect 13150 -3404 13166 -3370
rect 13100 -3420 13166 -3404
rect 13118 -3451 13148 -3420
rect 12728 -3816 12758 -3785
rect 12710 -3832 12776 -3816
rect 12710 -3866 12726 -3832
rect 12760 -3866 12776 -3832
rect 12710 -3882 12776 -3866
rect 13118 -3818 13148 -3787
rect 13100 -3834 13166 -3818
rect 13100 -3868 13116 -3834
rect 13150 -3868 13166 -3834
rect 13100 -3884 13166 -3868
rect 12714 -4164 12780 -4148
rect 12714 -4198 12730 -4164
rect 12764 -4198 12780 -4164
rect 12714 -4214 12780 -4198
rect 12732 -4236 12762 -4214
rect 13104 -4164 13170 -4148
rect 13104 -4198 13120 -4164
rect 13154 -4198 13170 -4164
rect 13104 -4214 13170 -4198
rect 13122 -4236 13152 -4214
rect 12732 -4342 12762 -4320
rect 12714 -4358 12780 -4342
rect 12714 -4392 12730 -4358
rect 12764 -4392 12780 -4358
rect 12714 -4408 12780 -4392
rect 13122 -4342 13152 -4320
rect 13104 -4358 13170 -4342
rect 13104 -4392 13120 -4358
rect 13154 -4392 13170 -4358
rect 13104 -4408 13170 -4392
rect 5254 -5012 5320 -4996
rect 5254 -5029 5270 -5012
rect 5187 -5046 5270 -5029
rect 5304 -5029 5320 -5012
rect 5512 -5012 5578 -4996
rect 5512 -5029 5528 -5012
rect 5304 -5046 5387 -5029
rect 5187 -5084 5387 -5046
rect 5445 -5046 5528 -5029
rect 5562 -5029 5578 -5012
rect 5770 -5012 5836 -4996
rect 5770 -5029 5786 -5012
rect 5562 -5046 5645 -5029
rect 5445 -5084 5645 -5046
rect 5703 -5046 5786 -5029
rect 5820 -5029 5836 -5012
rect 6028 -5012 6094 -4996
rect 6028 -5029 6044 -5012
rect 5820 -5046 5903 -5029
rect 5703 -5084 5903 -5046
rect 5961 -5046 6044 -5029
rect 6078 -5029 6094 -5012
rect 6286 -5012 6352 -4996
rect 6286 -5029 6302 -5012
rect 6078 -5046 6161 -5029
rect 5961 -5084 6161 -5046
rect 6219 -5046 6302 -5029
rect 6336 -5029 6352 -5012
rect 6544 -5012 6610 -4996
rect 6544 -5029 6560 -5012
rect 6336 -5046 6419 -5029
rect 6219 -5084 6419 -5046
rect 6477 -5046 6560 -5029
rect 6594 -5029 6610 -5012
rect 6802 -5012 6868 -4996
rect 6802 -5029 6818 -5012
rect 6594 -5046 6677 -5029
rect 6477 -5084 6677 -5046
rect 6735 -5046 6818 -5029
rect 6852 -5029 6868 -5012
rect 7060 -5012 7126 -4996
rect 7060 -5029 7076 -5012
rect 6852 -5046 6935 -5029
rect 6735 -5084 6935 -5046
rect 6993 -5046 7076 -5029
rect 7110 -5029 7126 -5012
rect 7924 -5012 7990 -4996
rect 7924 -5029 7940 -5012
rect 7110 -5046 7193 -5029
rect 6993 -5084 7193 -5046
rect 7857 -5046 7940 -5029
rect 7974 -5029 7990 -5012
rect 8182 -5012 8248 -4996
rect 8182 -5029 8198 -5012
rect 7974 -5046 8057 -5029
rect 7857 -5084 8057 -5046
rect 8115 -5046 8198 -5029
rect 8232 -5029 8248 -5012
rect 8440 -5012 8506 -4996
rect 8440 -5029 8456 -5012
rect 8232 -5046 8315 -5029
rect 8115 -5084 8315 -5046
rect 8373 -5046 8456 -5029
rect 8490 -5029 8506 -5012
rect 8698 -5012 8764 -4996
rect 8698 -5029 8714 -5012
rect 8490 -5046 8573 -5029
rect 8373 -5084 8573 -5046
rect 8631 -5046 8714 -5029
rect 8748 -5029 8764 -5012
rect 8956 -5012 9022 -4996
rect 8956 -5029 8972 -5012
rect 8748 -5046 8831 -5029
rect 8631 -5084 8831 -5046
rect 8889 -5046 8972 -5029
rect 9006 -5029 9022 -5012
rect 9214 -5012 9280 -4996
rect 9214 -5029 9230 -5012
rect 9006 -5046 9089 -5029
rect 8889 -5084 9089 -5046
rect 9147 -5046 9230 -5029
rect 9264 -5029 9280 -5012
rect 9472 -5012 9538 -4996
rect 9472 -5029 9488 -5012
rect 9264 -5046 9347 -5029
rect 9147 -5084 9347 -5046
rect 9405 -5046 9488 -5029
rect 9522 -5029 9538 -5012
rect 9730 -5012 9796 -4996
rect 9730 -5029 9746 -5012
rect 9522 -5046 9605 -5029
rect 9405 -5084 9605 -5046
rect 9663 -5046 9746 -5029
rect 9780 -5029 9796 -5012
rect 10587 -5011 10653 -4995
rect 10587 -5028 10603 -5011
rect 9780 -5046 9863 -5029
rect 9663 -5084 9863 -5046
rect 10520 -5045 10603 -5028
rect 10637 -5028 10653 -5011
rect 10845 -5011 10911 -4995
rect 10845 -5028 10861 -5011
rect 10637 -5045 10720 -5028
rect 10520 -5083 10720 -5045
rect 10778 -5045 10861 -5028
rect 10895 -5028 10911 -5011
rect 11103 -5011 11169 -4995
rect 11103 -5028 11119 -5011
rect 10895 -5045 10978 -5028
rect 10778 -5083 10978 -5045
rect 11036 -5045 11119 -5028
rect 11153 -5028 11169 -5011
rect 11361 -5011 11427 -4995
rect 11361 -5028 11377 -5011
rect 11153 -5045 11236 -5028
rect 11036 -5083 11236 -5045
rect 11294 -5045 11377 -5028
rect 11411 -5028 11427 -5011
rect 11619 -5011 11685 -4995
rect 11619 -5028 11635 -5011
rect 11411 -5045 11494 -5028
rect 11294 -5083 11494 -5045
rect 11552 -5045 11635 -5028
rect 11669 -5028 11685 -5011
rect 11877 -5011 11943 -4995
rect 11877 -5028 11893 -5011
rect 11669 -5045 11752 -5028
rect 11552 -5083 11752 -5045
rect 11810 -5045 11893 -5028
rect 11927 -5028 11943 -5011
rect 12135 -5011 12201 -4995
rect 12135 -5028 12151 -5011
rect 11927 -5045 12010 -5028
rect 11810 -5083 12010 -5045
rect 12068 -5045 12151 -5028
rect 12185 -5028 12201 -5011
rect 12393 -5011 12459 -4995
rect 12393 -5028 12409 -5011
rect 12185 -5045 12268 -5028
rect 12068 -5083 12268 -5045
rect 12326 -5045 12409 -5028
rect 12443 -5028 12459 -5011
rect 12443 -5045 12526 -5028
rect 12326 -5083 12526 -5045
rect 5187 -5322 5387 -5284
rect 5187 -5339 5270 -5322
rect 5254 -5356 5270 -5339
rect 5304 -5339 5387 -5322
rect 5445 -5322 5645 -5284
rect 5445 -5339 5528 -5322
rect 5304 -5356 5320 -5339
rect 5254 -5372 5320 -5356
rect 5512 -5356 5528 -5339
rect 5562 -5339 5645 -5322
rect 5703 -5322 5903 -5284
rect 5703 -5339 5786 -5322
rect 5562 -5356 5578 -5339
rect 5512 -5372 5578 -5356
rect 5770 -5356 5786 -5339
rect 5820 -5339 5903 -5322
rect 5961 -5322 6161 -5284
rect 5961 -5339 6044 -5322
rect 5820 -5356 5836 -5339
rect 5770 -5372 5836 -5356
rect 6028 -5356 6044 -5339
rect 6078 -5339 6161 -5322
rect 6219 -5322 6419 -5284
rect 6219 -5339 6302 -5322
rect 6078 -5356 6094 -5339
rect 6028 -5372 6094 -5356
rect 6286 -5356 6302 -5339
rect 6336 -5339 6419 -5322
rect 6477 -5322 6677 -5284
rect 6477 -5339 6560 -5322
rect 6336 -5356 6352 -5339
rect 6286 -5372 6352 -5356
rect 6544 -5356 6560 -5339
rect 6594 -5339 6677 -5322
rect 6735 -5322 6935 -5284
rect 6735 -5339 6818 -5322
rect 6594 -5356 6610 -5339
rect 6544 -5372 6610 -5356
rect 6802 -5356 6818 -5339
rect 6852 -5339 6935 -5322
rect 6993 -5322 7193 -5284
rect 6993 -5339 7076 -5322
rect 6852 -5356 6868 -5339
rect 6802 -5372 6868 -5356
rect 7060 -5356 7076 -5339
rect 7110 -5339 7193 -5322
rect 7857 -5322 8057 -5284
rect 7857 -5339 7940 -5322
rect 7110 -5356 7126 -5339
rect 7060 -5372 7126 -5356
rect 7924 -5356 7940 -5339
rect 7974 -5339 8057 -5322
rect 8115 -5322 8315 -5284
rect 8115 -5339 8198 -5322
rect 7974 -5356 7990 -5339
rect 7924 -5372 7990 -5356
rect 8182 -5356 8198 -5339
rect 8232 -5339 8315 -5322
rect 8373 -5322 8573 -5284
rect 8373 -5339 8456 -5322
rect 8232 -5356 8248 -5339
rect 8182 -5372 8248 -5356
rect 8440 -5356 8456 -5339
rect 8490 -5339 8573 -5322
rect 8631 -5322 8831 -5284
rect 8631 -5339 8714 -5322
rect 8490 -5356 8506 -5339
rect 8440 -5372 8506 -5356
rect 8698 -5356 8714 -5339
rect 8748 -5339 8831 -5322
rect 8889 -5322 9089 -5284
rect 8889 -5339 8972 -5322
rect 8748 -5356 8764 -5339
rect 8698 -5372 8764 -5356
rect 8956 -5356 8972 -5339
rect 9006 -5339 9089 -5322
rect 9147 -5322 9347 -5284
rect 9147 -5339 9230 -5322
rect 9006 -5356 9022 -5339
rect 8956 -5372 9022 -5356
rect 9214 -5356 9230 -5339
rect 9264 -5339 9347 -5322
rect 9405 -5322 9605 -5284
rect 9405 -5339 9488 -5322
rect 9264 -5356 9280 -5339
rect 9214 -5372 9280 -5356
rect 9472 -5356 9488 -5339
rect 9522 -5339 9605 -5322
rect 9663 -5322 9863 -5284
rect 9663 -5339 9746 -5322
rect 9522 -5356 9538 -5339
rect 9472 -5372 9538 -5356
rect 9730 -5356 9746 -5339
rect 9780 -5339 9863 -5322
rect 10520 -5321 10720 -5283
rect 10520 -5338 10603 -5321
rect 9780 -5356 9796 -5339
rect 9730 -5372 9796 -5356
rect 10587 -5355 10603 -5338
rect 10637 -5338 10720 -5321
rect 10778 -5321 10978 -5283
rect 10778 -5338 10861 -5321
rect 10637 -5355 10653 -5338
rect 10587 -5371 10653 -5355
rect 10845 -5355 10861 -5338
rect 10895 -5338 10978 -5321
rect 11036 -5321 11236 -5283
rect 11036 -5338 11119 -5321
rect 10895 -5355 10911 -5338
rect 10845 -5371 10911 -5355
rect 11103 -5355 11119 -5338
rect 11153 -5338 11236 -5321
rect 11294 -5321 11494 -5283
rect 11294 -5338 11377 -5321
rect 11153 -5355 11169 -5338
rect 11103 -5371 11169 -5355
rect 11361 -5355 11377 -5338
rect 11411 -5338 11494 -5321
rect 11552 -5321 11752 -5283
rect 11552 -5338 11635 -5321
rect 11411 -5355 11427 -5338
rect 11361 -5371 11427 -5355
rect 11619 -5355 11635 -5338
rect 11669 -5338 11752 -5321
rect 11810 -5321 12010 -5283
rect 11810 -5338 11893 -5321
rect 11669 -5355 11685 -5338
rect 11619 -5371 11685 -5355
rect 11877 -5355 11893 -5338
rect 11927 -5338 12010 -5321
rect 12068 -5321 12268 -5283
rect 12068 -5338 12151 -5321
rect 11927 -5355 11943 -5338
rect 11877 -5371 11943 -5355
rect 12135 -5355 12151 -5338
rect 12185 -5338 12268 -5321
rect 12326 -5321 12526 -5283
rect 12326 -5338 12409 -5321
rect 12185 -5355 12201 -5338
rect 12135 -5371 12201 -5355
rect 12393 -5355 12409 -5338
rect 12443 -5338 12526 -5321
rect 12443 -5355 12459 -5338
rect 12393 -5371 12459 -5355
rect 5254 -5430 5320 -5414
rect 5254 -5447 5270 -5430
rect 5187 -5464 5270 -5447
rect 5304 -5447 5320 -5430
rect 5512 -5430 5578 -5414
rect 5512 -5447 5528 -5430
rect 5304 -5464 5387 -5447
rect 5187 -5502 5387 -5464
rect 5445 -5464 5528 -5447
rect 5562 -5447 5578 -5430
rect 5770 -5430 5836 -5414
rect 5770 -5447 5786 -5430
rect 5562 -5464 5645 -5447
rect 5445 -5502 5645 -5464
rect 5703 -5464 5786 -5447
rect 5820 -5447 5836 -5430
rect 6028 -5430 6094 -5414
rect 6028 -5447 6044 -5430
rect 5820 -5464 5903 -5447
rect 5703 -5502 5903 -5464
rect 5961 -5464 6044 -5447
rect 6078 -5447 6094 -5430
rect 6286 -5430 6352 -5414
rect 6286 -5447 6302 -5430
rect 6078 -5464 6161 -5447
rect 5961 -5502 6161 -5464
rect 6219 -5464 6302 -5447
rect 6336 -5447 6352 -5430
rect 6544 -5430 6610 -5414
rect 6544 -5447 6560 -5430
rect 6336 -5464 6419 -5447
rect 6219 -5502 6419 -5464
rect 6477 -5464 6560 -5447
rect 6594 -5447 6610 -5430
rect 6802 -5430 6868 -5414
rect 6802 -5447 6818 -5430
rect 6594 -5464 6677 -5447
rect 6477 -5502 6677 -5464
rect 6735 -5464 6818 -5447
rect 6852 -5447 6868 -5430
rect 7060 -5430 7126 -5414
rect 7060 -5447 7076 -5430
rect 6852 -5464 6935 -5447
rect 6735 -5502 6935 -5464
rect 6993 -5464 7076 -5447
rect 7110 -5447 7126 -5430
rect 7924 -5430 7990 -5414
rect 7924 -5447 7940 -5430
rect 7110 -5464 7193 -5447
rect 6993 -5502 7193 -5464
rect 7857 -5464 7940 -5447
rect 7974 -5447 7990 -5430
rect 8182 -5430 8248 -5414
rect 8182 -5447 8198 -5430
rect 7974 -5464 8057 -5447
rect 7857 -5502 8057 -5464
rect 8115 -5464 8198 -5447
rect 8232 -5447 8248 -5430
rect 8440 -5430 8506 -5414
rect 8440 -5447 8456 -5430
rect 8232 -5464 8315 -5447
rect 8115 -5502 8315 -5464
rect 8373 -5464 8456 -5447
rect 8490 -5447 8506 -5430
rect 8698 -5430 8764 -5414
rect 8698 -5447 8714 -5430
rect 8490 -5464 8573 -5447
rect 8373 -5502 8573 -5464
rect 8631 -5464 8714 -5447
rect 8748 -5447 8764 -5430
rect 8956 -5430 9022 -5414
rect 8956 -5447 8972 -5430
rect 8748 -5464 8831 -5447
rect 8631 -5502 8831 -5464
rect 8889 -5464 8972 -5447
rect 9006 -5447 9022 -5430
rect 9214 -5430 9280 -5414
rect 9214 -5447 9230 -5430
rect 9006 -5464 9089 -5447
rect 8889 -5502 9089 -5464
rect 9147 -5464 9230 -5447
rect 9264 -5447 9280 -5430
rect 9472 -5430 9538 -5414
rect 9472 -5447 9488 -5430
rect 9264 -5464 9347 -5447
rect 9147 -5502 9347 -5464
rect 9405 -5464 9488 -5447
rect 9522 -5447 9538 -5430
rect 9730 -5430 9796 -5414
rect 9730 -5447 9746 -5430
rect 9522 -5464 9605 -5447
rect 9405 -5502 9605 -5464
rect 9663 -5464 9746 -5447
rect 9780 -5447 9796 -5430
rect 10587 -5429 10653 -5413
rect 10587 -5446 10603 -5429
rect 9780 -5464 9863 -5447
rect 9663 -5502 9863 -5464
rect 10520 -5463 10603 -5446
rect 10637 -5446 10653 -5429
rect 10845 -5429 10911 -5413
rect 10845 -5446 10861 -5429
rect 10637 -5463 10720 -5446
rect 10520 -5501 10720 -5463
rect 10778 -5463 10861 -5446
rect 10895 -5446 10911 -5429
rect 11103 -5429 11169 -5413
rect 11103 -5446 11119 -5429
rect 10895 -5463 10978 -5446
rect 10778 -5501 10978 -5463
rect 11036 -5463 11119 -5446
rect 11153 -5446 11169 -5429
rect 11361 -5429 11427 -5413
rect 11361 -5446 11377 -5429
rect 11153 -5463 11236 -5446
rect 11036 -5501 11236 -5463
rect 11294 -5463 11377 -5446
rect 11411 -5446 11427 -5429
rect 11619 -5429 11685 -5413
rect 11619 -5446 11635 -5429
rect 11411 -5463 11494 -5446
rect 11294 -5501 11494 -5463
rect 11552 -5463 11635 -5446
rect 11669 -5446 11685 -5429
rect 11877 -5429 11943 -5413
rect 11877 -5446 11893 -5429
rect 11669 -5463 11752 -5446
rect 11552 -5501 11752 -5463
rect 11810 -5463 11893 -5446
rect 11927 -5446 11943 -5429
rect 12135 -5429 12201 -5413
rect 12135 -5446 12151 -5429
rect 11927 -5463 12010 -5446
rect 11810 -5501 12010 -5463
rect 12068 -5463 12151 -5446
rect 12185 -5446 12201 -5429
rect 12393 -5429 12459 -5413
rect 12393 -5446 12409 -5429
rect 12185 -5463 12268 -5446
rect 12068 -5501 12268 -5463
rect 12326 -5463 12409 -5446
rect 12443 -5446 12459 -5429
rect 12443 -5463 12526 -5446
rect 12326 -5501 12526 -5463
rect 5187 -5740 5387 -5702
rect 5187 -5757 5270 -5740
rect 5254 -5774 5270 -5757
rect 5304 -5757 5387 -5740
rect 5445 -5740 5645 -5702
rect 5445 -5757 5528 -5740
rect 5304 -5774 5320 -5757
rect 5254 -5790 5320 -5774
rect 5512 -5774 5528 -5757
rect 5562 -5757 5645 -5740
rect 5703 -5740 5903 -5702
rect 5703 -5757 5786 -5740
rect 5562 -5774 5578 -5757
rect 5512 -5790 5578 -5774
rect 5770 -5774 5786 -5757
rect 5820 -5757 5903 -5740
rect 5961 -5740 6161 -5702
rect 5961 -5757 6044 -5740
rect 5820 -5774 5836 -5757
rect 5770 -5790 5836 -5774
rect 6028 -5774 6044 -5757
rect 6078 -5757 6161 -5740
rect 6219 -5740 6419 -5702
rect 6219 -5757 6302 -5740
rect 6078 -5774 6094 -5757
rect 6028 -5790 6094 -5774
rect 6286 -5774 6302 -5757
rect 6336 -5757 6419 -5740
rect 6477 -5740 6677 -5702
rect 6477 -5757 6560 -5740
rect 6336 -5774 6352 -5757
rect 6286 -5790 6352 -5774
rect 6544 -5774 6560 -5757
rect 6594 -5757 6677 -5740
rect 6735 -5740 6935 -5702
rect 6735 -5757 6818 -5740
rect 6594 -5774 6610 -5757
rect 6544 -5790 6610 -5774
rect 6802 -5774 6818 -5757
rect 6852 -5757 6935 -5740
rect 6993 -5740 7193 -5702
rect 6993 -5757 7076 -5740
rect 6852 -5774 6868 -5757
rect 6802 -5790 6868 -5774
rect 7060 -5774 7076 -5757
rect 7110 -5757 7193 -5740
rect 7857 -5740 8057 -5702
rect 7857 -5757 7940 -5740
rect 7110 -5774 7126 -5757
rect 7060 -5790 7126 -5774
rect 7924 -5774 7940 -5757
rect 7974 -5757 8057 -5740
rect 8115 -5740 8315 -5702
rect 8115 -5757 8198 -5740
rect 7974 -5774 7990 -5757
rect 7924 -5790 7990 -5774
rect 8182 -5774 8198 -5757
rect 8232 -5757 8315 -5740
rect 8373 -5740 8573 -5702
rect 8373 -5757 8456 -5740
rect 8232 -5774 8248 -5757
rect 8182 -5790 8248 -5774
rect 8440 -5774 8456 -5757
rect 8490 -5757 8573 -5740
rect 8631 -5740 8831 -5702
rect 8631 -5757 8714 -5740
rect 8490 -5774 8506 -5757
rect 8440 -5790 8506 -5774
rect 8698 -5774 8714 -5757
rect 8748 -5757 8831 -5740
rect 8889 -5740 9089 -5702
rect 8889 -5757 8972 -5740
rect 8748 -5774 8764 -5757
rect 8698 -5790 8764 -5774
rect 8956 -5774 8972 -5757
rect 9006 -5757 9089 -5740
rect 9147 -5740 9347 -5702
rect 9147 -5757 9230 -5740
rect 9006 -5774 9022 -5757
rect 8956 -5790 9022 -5774
rect 9214 -5774 9230 -5757
rect 9264 -5757 9347 -5740
rect 9405 -5740 9605 -5702
rect 9405 -5757 9488 -5740
rect 9264 -5774 9280 -5757
rect 9214 -5790 9280 -5774
rect 9472 -5774 9488 -5757
rect 9522 -5757 9605 -5740
rect 9663 -5740 9863 -5702
rect 9663 -5757 9746 -5740
rect 9522 -5774 9538 -5757
rect 9472 -5790 9538 -5774
rect 9730 -5774 9746 -5757
rect 9780 -5757 9863 -5740
rect 10520 -5739 10720 -5701
rect 10520 -5756 10603 -5739
rect 9780 -5774 9796 -5757
rect 9730 -5790 9796 -5774
rect 10587 -5773 10603 -5756
rect 10637 -5756 10720 -5739
rect 10778 -5739 10978 -5701
rect 10778 -5756 10861 -5739
rect 10637 -5773 10653 -5756
rect 10587 -5789 10653 -5773
rect 10845 -5773 10861 -5756
rect 10895 -5756 10978 -5739
rect 11036 -5739 11236 -5701
rect 11036 -5756 11119 -5739
rect 10895 -5773 10911 -5756
rect 10845 -5789 10911 -5773
rect 11103 -5773 11119 -5756
rect 11153 -5756 11236 -5739
rect 11294 -5739 11494 -5701
rect 11294 -5756 11377 -5739
rect 11153 -5773 11169 -5756
rect 11103 -5789 11169 -5773
rect 11361 -5773 11377 -5756
rect 11411 -5756 11494 -5739
rect 11552 -5739 11752 -5701
rect 11552 -5756 11635 -5739
rect 11411 -5773 11427 -5756
rect 11361 -5789 11427 -5773
rect 11619 -5773 11635 -5756
rect 11669 -5756 11752 -5739
rect 11810 -5739 12010 -5701
rect 11810 -5756 11893 -5739
rect 11669 -5773 11685 -5756
rect 11619 -5789 11685 -5773
rect 11877 -5773 11893 -5756
rect 11927 -5756 12010 -5739
rect 12068 -5739 12268 -5701
rect 12068 -5756 12151 -5739
rect 11927 -5773 11943 -5756
rect 11877 -5789 11943 -5773
rect 12135 -5773 12151 -5756
rect 12185 -5756 12268 -5739
rect 12326 -5739 12526 -5701
rect 12326 -5756 12409 -5739
rect 12185 -5773 12201 -5756
rect 12135 -5789 12201 -5773
rect 12393 -5773 12409 -5756
rect 12443 -5756 12526 -5739
rect 12443 -5773 12459 -5756
rect 12393 -5789 12459 -5773
rect 5254 -5848 5320 -5832
rect 5254 -5865 5270 -5848
rect 5187 -5882 5270 -5865
rect 5304 -5865 5320 -5848
rect 5512 -5848 5578 -5832
rect 5512 -5865 5528 -5848
rect 5304 -5882 5387 -5865
rect 5187 -5920 5387 -5882
rect 5445 -5882 5528 -5865
rect 5562 -5865 5578 -5848
rect 5770 -5848 5836 -5832
rect 5770 -5865 5786 -5848
rect 5562 -5882 5645 -5865
rect 5445 -5920 5645 -5882
rect 5703 -5882 5786 -5865
rect 5820 -5865 5836 -5848
rect 6028 -5848 6094 -5832
rect 6028 -5865 6044 -5848
rect 5820 -5882 5903 -5865
rect 5703 -5920 5903 -5882
rect 5961 -5882 6044 -5865
rect 6078 -5865 6094 -5848
rect 6286 -5848 6352 -5832
rect 6286 -5865 6302 -5848
rect 6078 -5882 6161 -5865
rect 5961 -5920 6161 -5882
rect 6219 -5882 6302 -5865
rect 6336 -5865 6352 -5848
rect 6544 -5848 6610 -5832
rect 6544 -5865 6560 -5848
rect 6336 -5882 6419 -5865
rect 6219 -5920 6419 -5882
rect 6477 -5882 6560 -5865
rect 6594 -5865 6610 -5848
rect 6802 -5848 6868 -5832
rect 6802 -5865 6818 -5848
rect 6594 -5882 6677 -5865
rect 6477 -5920 6677 -5882
rect 6735 -5882 6818 -5865
rect 6852 -5865 6868 -5848
rect 7060 -5848 7126 -5832
rect 7060 -5865 7076 -5848
rect 6852 -5882 6935 -5865
rect 6735 -5920 6935 -5882
rect 6993 -5882 7076 -5865
rect 7110 -5865 7126 -5848
rect 7924 -5848 7990 -5832
rect 7924 -5865 7940 -5848
rect 7110 -5882 7193 -5865
rect 6993 -5920 7193 -5882
rect 7857 -5882 7940 -5865
rect 7974 -5865 7990 -5848
rect 8182 -5848 8248 -5832
rect 8182 -5865 8198 -5848
rect 7974 -5882 8057 -5865
rect 7857 -5920 8057 -5882
rect 8115 -5882 8198 -5865
rect 8232 -5865 8248 -5848
rect 8440 -5848 8506 -5832
rect 8440 -5865 8456 -5848
rect 8232 -5882 8315 -5865
rect 8115 -5920 8315 -5882
rect 8373 -5882 8456 -5865
rect 8490 -5865 8506 -5848
rect 8698 -5848 8764 -5832
rect 8698 -5865 8714 -5848
rect 8490 -5882 8573 -5865
rect 8373 -5920 8573 -5882
rect 8631 -5882 8714 -5865
rect 8748 -5865 8764 -5848
rect 8956 -5848 9022 -5832
rect 8956 -5865 8972 -5848
rect 8748 -5882 8831 -5865
rect 8631 -5920 8831 -5882
rect 8889 -5882 8972 -5865
rect 9006 -5865 9022 -5848
rect 9214 -5848 9280 -5832
rect 9214 -5865 9230 -5848
rect 9006 -5882 9089 -5865
rect 8889 -5920 9089 -5882
rect 9147 -5882 9230 -5865
rect 9264 -5865 9280 -5848
rect 9472 -5848 9538 -5832
rect 9472 -5865 9488 -5848
rect 9264 -5882 9347 -5865
rect 9147 -5920 9347 -5882
rect 9405 -5882 9488 -5865
rect 9522 -5865 9538 -5848
rect 9730 -5848 9796 -5832
rect 9730 -5865 9746 -5848
rect 9522 -5882 9605 -5865
rect 9405 -5920 9605 -5882
rect 9663 -5882 9746 -5865
rect 9780 -5865 9796 -5848
rect 10587 -5847 10653 -5831
rect 10587 -5864 10603 -5847
rect 9780 -5882 9863 -5865
rect 9663 -5920 9863 -5882
rect 10520 -5881 10603 -5864
rect 10637 -5864 10653 -5847
rect 10845 -5847 10911 -5831
rect 10845 -5864 10861 -5847
rect 10637 -5881 10720 -5864
rect 10520 -5919 10720 -5881
rect 10778 -5881 10861 -5864
rect 10895 -5864 10911 -5847
rect 11103 -5847 11169 -5831
rect 11103 -5864 11119 -5847
rect 10895 -5881 10978 -5864
rect 10778 -5919 10978 -5881
rect 11036 -5881 11119 -5864
rect 11153 -5864 11169 -5847
rect 11361 -5847 11427 -5831
rect 11361 -5864 11377 -5847
rect 11153 -5881 11236 -5864
rect 11036 -5919 11236 -5881
rect 11294 -5881 11377 -5864
rect 11411 -5864 11427 -5847
rect 11619 -5847 11685 -5831
rect 11619 -5864 11635 -5847
rect 11411 -5881 11494 -5864
rect 11294 -5919 11494 -5881
rect 11552 -5881 11635 -5864
rect 11669 -5864 11685 -5847
rect 11877 -5847 11943 -5831
rect 11877 -5864 11893 -5847
rect 11669 -5881 11752 -5864
rect 11552 -5919 11752 -5881
rect 11810 -5881 11893 -5864
rect 11927 -5864 11943 -5847
rect 12135 -5847 12201 -5831
rect 12135 -5864 12151 -5847
rect 11927 -5881 12010 -5864
rect 11810 -5919 12010 -5881
rect 12068 -5881 12151 -5864
rect 12185 -5864 12201 -5847
rect 12393 -5847 12459 -5831
rect 12393 -5864 12409 -5847
rect 12185 -5881 12268 -5864
rect 12068 -5919 12268 -5881
rect 12326 -5881 12409 -5864
rect 12443 -5864 12459 -5847
rect 12443 -5881 12526 -5864
rect 12326 -5919 12526 -5881
rect 5187 -6158 5387 -6120
rect 5187 -6175 5270 -6158
rect 5254 -6192 5270 -6175
rect 5304 -6175 5387 -6158
rect 5445 -6158 5645 -6120
rect 5445 -6175 5528 -6158
rect 5304 -6192 5320 -6175
rect 5254 -6208 5320 -6192
rect 5512 -6192 5528 -6175
rect 5562 -6175 5645 -6158
rect 5703 -6158 5903 -6120
rect 5703 -6175 5786 -6158
rect 5562 -6192 5578 -6175
rect 5512 -6208 5578 -6192
rect 5770 -6192 5786 -6175
rect 5820 -6175 5903 -6158
rect 5961 -6158 6161 -6120
rect 5961 -6175 6044 -6158
rect 5820 -6192 5836 -6175
rect 5770 -6208 5836 -6192
rect 6028 -6192 6044 -6175
rect 6078 -6175 6161 -6158
rect 6219 -6158 6419 -6120
rect 6219 -6175 6302 -6158
rect 6078 -6192 6094 -6175
rect 6028 -6208 6094 -6192
rect 6286 -6192 6302 -6175
rect 6336 -6175 6419 -6158
rect 6477 -6158 6677 -6120
rect 6477 -6175 6560 -6158
rect 6336 -6192 6352 -6175
rect 6286 -6208 6352 -6192
rect 6544 -6192 6560 -6175
rect 6594 -6175 6677 -6158
rect 6735 -6158 6935 -6120
rect 6735 -6175 6818 -6158
rect 6594 -6192 6610 -6175
rect 6544 -6208 6610 -6192
rect 6802 -6192 6818 -6175
rect 6852 -6175 6935 -6158
rect 6993 -6158 7193 -6120
rect 6993 -6175 7076 -6158
rect 6852 -6192 6868 -6175
rect 6802 -6208 6868 -6192
rect 7060 -6192 7076 -6175
rect 7110 -6175 7193 -6158
rect 7857 -6158 8057 -6120
rect 7857 -6175 7940 -6158
rect 7110 -6192 7126 -6175
rect 7060 -6208 7126 -6192
rect 7924 -6192 7940 -6175
rect 7974 -6175 8057 -6158
rect 8115 -6158 8315 -6120
rect 8115 -6175 8198 -6158
rect 7974 -6192 7990 -6175
rect 7924 -6208 7990 -6192
rect 8182 -6192 8198 -6175
rect 8232 -6175 8315 -6158
rect 8373 -6158 8573 -6120
rect 8373 -6175 8456 -6158
rect 8232 -6192 8248 -6175
rect 8182 -6208 8248 -6192
rect 8440 -6192 8456 -6175
rect 8490 -6175 8573 -6158
rect 8631 -6158 8831 -6120
rect 8631 -6175 8714 -6158
rect 8490 -6192 8506 -6175
rect 8440 -6208 8506 -6192
rect 8698 -6192 8714 -6175
rect 8748 -6175 8831 -6158
rect 8889 -6158 9089 -6120
rect 8889 -6175 8972 -6158
rect 8748 -6192 8764 -6175
rect 8698 -6208 8764 -6192
rect 8956 -6192 8972 -6175
rect 9006 -6175 9089 -6158
rect 9147 -6158 9347 -6120
rect 9147 -6175 9230 -6158
rect 9006 -6192 9022 -6175
rect 8956 -6208 9022 -6192
rect 9214 -6192 9230 -6175
rect 9264 -6175 9347 -6158
rect 9405 -6158 9605 -6120
rect 9405 -6175 9488 -6158
rect 9264 -6192 9280 -6175
rect 9214 -6208 9280 -6192
rect 9472 -6192 9488 -6175
rect 9522 -6175 9605 -6158
rect 9663 -6158 9863 -6120
rect 9663 -6175 9746 -6158
rect 9522 -6192 9538 -6175
rect 9472 -6208 9538 -6192
rect 9730 -6192 9746 -6175
rect 9780 -6175 9863 -6158
rect 10520 -6157 10720 -6119
rect 10520 -6174 10603 -6157
rect 9780 -6192 9796 -6175
rect 9730 -6208 9796 -6192
rect 10587 -6191 10603 -6174
rect 10637 -6174 10720 -6157
rect 10778 -6157 10978 -6119
rect 10778 -6174 10861 -6157
rect 10637 -6191 10653 -6174
rect 10587 -6207 10653 -6191
rect 10845 -6191 10861 -6174
rect 10895 -6174 10978 -6157
rect 11036 -6157 11236 -6119
rect 11036 -6174 11119 -6157
rect 10895 -6191 10911 -6174
rect 10845 -6207 10911 -6191
rect 11103 -6191 11119 -6174
rect 11153 -6174 11236 -6157
rect 11294 -6157 11494 -6119
rect 11294 -6174 11377 -6157
rect 11153 -6191 11169 -6174
rect 11103 -6207 11169 -6191
rect 11361 -6191 11377 -6174
rect 11411 -6174 11494 -6157
rect 11552 -6157 11752 -6119
rect 11552 -6174 11635 -6157
rect 11411 -6191 11427 -6174
rect 11361 -6207 11427 -6191
rect 11619 -6191 11635 -6174
rect 11669 -6174 11752 -6157
rect 11810 -6157 12010 -6119
rect 11810 -6174 11893 -6157
rect 11669 -6191 11685 -6174
rect 11619 -6207 11685 -6191
rect 11877 -6191 11893 -6174
rect 11927 -6174 12010 -6157
rect 12068 -6157 12268 -6119
rect 12068 -6174 12151 -6157
rect 11927 -6191 11943 -6174
rect 11877 -6207 11943 -6191
rect 12135 -6191 12151 -6174
rect 12185 -6174 12268 -6157
rect 12326 -6157 12526 -6119
rect 12326 -6174 12409 -6157
rect 12185 -6191 12201 -6174
rect 12135 -6207 12201 -6191
rect 12393 -6191 12409 -6174
rect 12443 -6174 12526 -6157
rect 12443 -6191 12459 -6174
rect 12393 -6207 12459 -6191
rect 5254 -6266 5320 -6250
rect 5254 -6283 5270 -6266
rect 5187 -6300 5270 -6283
rect 5304 -6283 5320 -6266
rect 5512 -6266 5578 -6250
rect 5512 -6283 5528 -6266
rect 5304 -6300 5387 -6283
rect 5187 -6338 5387 -6300
rect 5445 -6300 5528 -6283
rect 5562 -6283 5578 -6266
rect 5770 -6266 5836 -6250
rect 5770 -6283 5786 -6266
rect 5562 -6300 5645 -6283
rect 5445 -6338 5645 -6300
rect 5703 -6300 5786 -6283
rect 5820 -6283 5836 -6266
rect 6028 -6266 6094 -6250
rect 6028 -6283 6044 -6266
rect 5820 -6300 5903 -6283
rect 5703 -6338 5903 -6300
rect 5961 -6300 6044 -6283
rect 6078 -6283 6094 -6266
rect 6286 -6266 6352 -6250
rect 6286 -6283 6302 -6266
rect 6078 -6300 6161 -6283
rect 5961 -6338 6161 -6300
rect 6219 -6300 6302 -6283
rect 6336 -6283 6352 -6266
rect 6544 -6266 6610 -6250
rect 6544 -6283 6560 -6266
rect 6336 -6300 6419 -6283
rect 6219 -6338 6419 -6300
rect 6477 -6300 6560 -6283
rect 6594 -6283 6610 -6266
rect 6802 -6266 6868 -6250
rect 6802 -6283 6818 -6266
rect 6594 -6300 6677 -6283
rect 6477 -6338 6677 -6300
rect 6735 -6300 6818 -6283
rect 6852 -6283 6868 -6266
rect 7060 -6266 7126 -6250
rect 7060 -6283 7076 -6266
rect 6852 -6300 6935 -6283
rect 6735 -6338 6935 -6300
rect 6993 -6300 7076 -6283
rect 7110 -6283 7126 -6266
rect 7924 -6266 7990 -6250
rect 7924 -6283 7940 -6266
rect 7110 -6300 7193 -6283
rect 6993 -6338 7193 -6300
rect 7857 -6300 7940 -6283
rect 7974 -6283 7990 -6266
rect 8182 -6266 8248 -6250
rect 8182 -6283 8198 -6266
rect 7974 -6300 8057 -6283
rect 7857 -6338 8057 -6300
rect 8115 -6300 8198 -6283
rect 8232 -6283 8248 -6266
rect 8440 -6266 8506 -6250
rect 8440 -6283 8456 -6266
rect 8232 -6300 8315 -6283
rect 8115 -6338 8315 -6300
rect 8373 -6300 8456 -6283
rect 8490 -6283 8506 -6266
rect 8698 -6266 8764 -6250
rect 8698 -6283 8714 -6266
rect 8490 -6300 8573 -6283
rect 8373 -6338 8573 -6300
rect 8631 -6300 8714 -6283
rect 8748 -6283 8764 -6266
rect 8956 -6266 9022 -6250
rect 8956 -6283 8972 -6266
rect 8748 -6300 8831 -6283
rect 8631 -6338 8831 -6300
rect 8889 -6300 8972 -6283
rect 9006 -6283 9022 -6266
rect 9214 -6266 9280 -6250
rect 9214 -6283 9230 -6266
rect 9006 -6300 9089 -6283
rect 8889 -6338 9089 -6300
rect 9147 -6300 9230 -6283
rect 9264 -6283 9280 -6266
rect 9472 -6266 9538 -6250
rect 9472 -6283 9488 -6266
rect 9264 -6300 9347 -6283
rect 9147 -6338 9347 -6300
rect 9405 -6300 9488 -6283
rect 9522 -6283 9538 -6266
rect 9730 -6266 9796 -6250
rect 9730 -6283 9746 -6266
rect 9522 -6300 9605 -6283
rect 9405 -6338 9605 -6300
rect 9663 -6300 9746 -6283
rect 9780 -6283 9796 -6266
rect 10587 -6265 10653 -6249
rect 10587 -6282 10603 -6265
rect 9780 -6300 9863 -6283
rect 9663 -6338 9863 -6300
rect 10520 -6299 10603 -6282
rect 10637 -6282 10653 -6265
rect 10845 -6265 10911 -6249
rect 10845 -6282 10861 -6265
rect 10637 -6299 10720 -6282
rect 10520 -6337 10720 -6299
rect 10778 -6299 10861 -6282
rect 10895 -6282 10911 -6265
rect 11103 -6265 11169 -6249
rect 11103 -6282 11119 -6265
rect 10895 -6299 10978 -6282
rect 10778 -6337 10978 -6299
rect 11036 -6299 11119 -6282
rect 11153 -6282 11169 -6265
rect 11361 -6265 11427 -6249
rect 11361 -6282 11377 -6265
rect 11153 -6299 11236 -6282
rect 11036 -6337 11236 -6299
rect 11294 -6299 11377 -6282
rect 11411 -6282 11427 -6265
rect 11619 -6265 11685 -6249
rect 11619 -6282 11635 -6265
rect 11411 -6299 11494 -6282
rect 11294 -6337 11494 -6299
rect 11552 -6299 11635 -6282
rect 11669 -6282 11685 -6265
rect 11877 -6265 11943 -6249
rect 11877 -6282 11893 -6265
rect 11669 -6299 11752 -6282
rect 11552 -6337 11752 -6299
rect 11810 -6299 11893 -6282
rect 11927 -6282 11943 -6265
rect 12135 -6265 12201 -6249
rect 12135 -6282 12151 -6265
rect 11927 -6299 12010 -6282
rect 11810 -6337 12010 -6299
rect 12068 -6299 12151 -6282
rect 12185 -6282 12201 -6265
rect 12393 -6265 12459 -6249
rect 12393 -6282 12409 -6265
rect 12185 -6299 12268 -6282
rect 12068 -6337 12268 -6299
rect 12326 -6299 12409 -6282
rect 12443 -6282 12459 -6265
rect 12443 -6299 12526 -6282
rect 12326 -6337 12526 -6299
rect 5187 -6576 5387 -6538
rect 5187 -6593 5270 -6576
rect 5254 -6610 5270 -6593
rect 5304 -6593 5387 -6576
rect 5445 -6576 5645 -6538
rect 5445 -6593 5528 -6576
rect 5304 -6610 5320 -6593
rect 5254 -6626 5320 -6610
rect 5512 -6610 5528 -6593
rect 5562 -6593 5645 -6576
rect 5703 -6576 5903 -6538
rect 5703 -6593 5786 -6576
rect 5562 -6610 5578 -6593
rect 5512 -6626 5578 -6610
rect 5770 -6610 5786 -6593
rect 5820 -6593 5903 -6576
rect 5961 -6576 6161 -6538
rect 5961 -6593 6044 -6576
rect 5820 -6610 5836 -6593
rect 5770 -6626 5836 -6610
rect 6028 -6610 6044 -6593
rect 6078 -6593 6161 -6576
rect 6219 -6576 6419 -6538
rect 6219 -6593 6302 -6576
rect 6078 -6610 6094 -6593
rect 6028 -6626 6094 -6610
rect 6286 -6610 6302 -6593
rect 6336 -6593 6419 -6576
rect 6477 -6576 6677 -6538
rect 6477 -6593 6560 -6576
rect 6336 -6610 6352 -6593
rect 6286 -6626 6352 -6610
rect 6544 -6610 6560 -6593
rect 6594 -6593 6677 -6576
rect 6735 -6576 6935 -6538
rect 6735 -6593 6818 -6576
rect 6594 -6610 6610 -6593
rect 6544 -6626 6610 -6610
rect 6802 -6610 6818 -6593
rect 6852 -6593 6935 -6576
rect 6993 -6576 7193 -6538
rect 6993 -6593 7076 -6576
rect 6852 -6610 6868 -6593
rect 6802 -6626 6868 -6610
rect 7060 -6610 7076 -6593
rect 7110 -6593 7193 -6576
rect 7857 -6576 8057 -6538
rect 7857 -6593 7940 -6576
rect 7110 -6610 7126 -6593
rect 7060 -6626 7126 -6610
rect 7924 -6610 7940 -6593
rect 7974 -6593 8057 -6576
rect 8115 -6576 8315 -6538
rect 8115 -6593 8198 -6576
rect 7974 -6610 7990 -6593
rect 7924 -6626 7990 -6610
rect 8182 -6610 8198 -6593
rect 8232 -6593 8315 -6576
rect 8373 -6576 8573 -6538
rect 8373 -6593 8456 -6576
rect 8232 -6610 8248 -6593
rect 8182 -6626 8248 -6610
rect 8440 -6610 8456 -6593
rect 8490 -6593 8573 -6576
rect 8631 -6576 8831 -6538
rect 8631 -6593 8714 -6576
rect 8490 -6610 8506 -6593
rect 8440 -6626 8506 -6610
rect 8698 -6610 8714 -6593
rect 8748 -6593 8831 -6576
rect 8889 -6576 9089 -6538
rect 8889 -6593 8972 -6576
rect 8748 -6610 8764 -6593
rect 8698 -6626 8764 -6610
rect 8956 -6610 8972 -6593
rect 9006 -6593 9089 -6576
rect 9147 -6576 9347 -6538
rect 9147 -6593 9230 -6576
rect 9006 -6610 9022 -6593
rect 8956 -6626 9022 -6610
rect 9214 -6610 9230 -6593
rect 9264 -6593 9347 -6576
rect 9405 -6576 9605 -6538
rect 9405 -6593 9488 -6576
rect 9264 -6610 9280 -6593
rect 9214 -6626 9280 -6610
rect 9472 -6610 9488 -6593
rect 9522 -6593 9605 -6576
rect 9663 -6576 9863 -6538
rect 9663 -6593 9746 -6576
rect 9522 -6610 9538 -6593
rect 9472 -6626 9538 -6610
rect 9730 -6610 9746 -6593
rect 9780 -6593 9863 -6576
rect 10520 -6575 10720 -6537
rect 10520 -6592 10603 -6575
rect 9780 -6610 9796 -6593
rect 9730 -6626 9796 -6610
rect 10587 -6609 10603 -6592
rect 10637 -6592 10720 -6575
rect 10778 -6575 10978 -6537
rect 10778 -6592 10861 -6575
rect 10637 -6609 10653 -6592
rect 10587 -6625 10653 -6609
rect 10845 -6609 10861 -6592
rect 10895 -6592 10978 -6575
rect 11036 -6575 11236 -6537
rect 11036 -6592 11119 -6575
rect 10895 -6609 10911 -6592
rect 10845 -6625 10911 -6609
rect 11103 -6609 11119 -6592
rect 11153 -6592 11236 -6575
rect 11294 -6575 11494 -6537
rect 11294 -6592 11377 -6575
rect 11153 -6609 11169 -6592
rect 11103 -6625 11169 -6609
rect 11361 -6609 11377 -6592
rect 11411 -6592 11494 -6575
rect 11552 -6575 11752 -6537
rect 11552 -6592 11635 -6575
rect 11411 -6609 11427 -6592
rect 11361 -6625 11427 -6609
rect 11619 -6609 11635 -6592
rect 11669 -6592 11752 -6575
rect 11810 -6575 12010 -6537
rect 11810 -6592 11893 -6575
rect 11669 -6609 11685 -6592
rect 11619 -6625 11685 -6609
rect 11877 -6609 11893 -6592
rect 11927 -6592 12010 -6575
rect 12068 -6575 12268 -6537
rect 12068 -6592 12151 -6575
rect 11927 -6609 11943 -6592
rect 11877 -6625 11943 -6609
rect 12135 -6609 12151 -6592
rect 12185 -6592 12268 -6575
rect 12326 -6575 12526 -6537
rect 12326 -6592 12409 -6575
rect 12185 -6609 12201 -6592
rect 12135 -6625 12201 -6609
rect 12393 -6609 12409 -6592
rect 12443 -6592 12526 -6575
rect 12443 -6609 12459 -6592
rect 12393 -6625 12459 -6609
rect 5254 -6684 5320 -6668
rect 5254 -6701 5270 -6684
rect 5187 -6718 5270 -6701
rect 5304 -6701 5320 -6684
rect 5512 -6684 5578 -6668
rect 5512 -6701 5528 -6684
rect 5304 -6718 5387 -6701
rect 5187 -6756 5387 -6718
rect 5445 -6718 5528 -6701
rect 5562 -6701 5578 -6684
rect 5770 -6684 5836 -6668
rect 5770 -6701 5786 -6684
rect 5562 -6718 5645 -6701
rect 5445 -6756 5645 -6718
rect 5703 -6718 5786 -6701
rect 5820 -6701 5836 -6684
rect 6028 -6684 6094 -6668
rect 6028 -6701 6044 -6684
rect 5820 -6718 5903 -6701
rect 5703 -6756 5903 -6718
rect 5961 -6718 6044 -6701
rect 6078 -6701 6094 -6684
rect 6286 -6684 6352 -6668
rect 6286 -6701 6302 -6684
rect 6078 -6718 6161 -6701
rect 5961 -6756 6161 -6718
rect 6219 -6718 6302 -6701
rect 6336 -6701 6352 -6684
rect 6544 -6684 6610 -6668
rect 6544 -6701 6560 -6684
rect 6336 -6718 6419 -6701
rect 6219 -6756 6419 -6718
rect 6477 -6718 6560 -6701
rect 6594 -6701 6610 -6684
rect 6802 -6684 6868 -6668
rect 6802 -6701 6818 -6684
rect 6594 -6718 6677 -6701
rect 6477 -6756 6677 -6718
rect 6735 -6718 6818 -6701
rect 6852 -6701 6868 -6684
rect 7060 -6684 7126 -6668
rect 7060 -6701 7076 -6684
rect 6852 -6718 6935 -6701
rect 6735 -6756 6935 -6718
rect 6993 -6718 7076 -6701
rect 7110 -6701 7126 -6684
rect 7924 -6684 7990 -6668
rect 7924 -6701 7940 -6684
rect 7110 -6718 7193 -6701
rect 6993 -6756 7193 -6718
rect 7857 -6718 7940 -6701
rect 7974 -6701 7990 -6684
rect 8182 -6684 8248 -6668
rect 8182 -6701 8198 -6684
rect 7974 -6718 8057 -6701
rect 7857 -6756 8057 -6718
rect 8115 -6718 8198 -6701
rect 8232 -6701 8248 -6684
rect 8440 -6684 8506 -6668
rect 8440 -6701 8456 -6684
rect 8232 -6718 8315 -6701
rect 8115 -6756 8315 -6718
rect 8373 -6718 8456 -6701
rect 8490 -6701 8506 -6684
rect 8698 -6684 8764 -6668
rect 8698 -6701 8714 -6684
rect 8490 -6718 8573 -6701
rect 8373 -6756 8573 -6718
rect 8631 -6718 8714 -6701
rect 8748 -6701 8764 -6684
rect 8956 -6684 9022 -6668
rect 8956 -6701 8972 -6684
rect 8748 -6718 8831 -6701
rect 8631 -6756 8831 -6718
rect 8889 -6718 8972 -6701
rect 9006 -6701 9022 -6684
rect 9214 -6684 9280 -6668
rect 9214 -6701 9230 -6684
rect 9006 -6718 9089 -6701
rect 8889 -6756 9089 -6718
rect 9147 -6718 9230 -6701
rect 9264 -6701 9280 -6684
rect 9472 -6684 9538 -6668
rect 9472 -6701 9488 -6684
rect 9264 -6718 9347 -6701
rect 9147 -6756 9347 -6718
rect 9405 -6718 9488 -6701
rect 9522 -6701 9538 -6684
rect 9730 -6684 9796 -6668
rect 9730 -6701 9746 -6684
rect 9522 -6718 9605 -6701
rect 9405 -6756 9605 -6718
rect 9663 -6718 9746 -6701
rect 9780 -6701 9796 -6684
rect 10587 -6683 10653 -6667
rect 10587 -6700 10603 -6683
rect 9780 -6718 9863 -6701
rect 9663 -6756 9863 -6718
rect 10520 -6717 10603 -6700
rect 10637 -6700 10653 -6683
rect 10845 -6683 10911 -6667
rect 10845 -6700 10861 -6683
rect 10637 -6717 10720 -6700
rect 10520 -6755 10720 -6717
rect 10778 -6717 10861 -6700
rect 10895 -6700 10911 -6683
rect 11103 -6683 11169 -6667
rect 11103 -6700 11119 -6683
rect 10895 -6717 10978 -6700
rect 10778 -6755 10978 -6717
rect 11036 -6717 11119 -6700
rect 11153 -6700 11169 -6683
rect 11361 -6683 11427 -6667
rect 11361 -6700 11377 -6683
rect 11153 -6717 11236 -6700
rect 11036 -6755 11236 -6717
rect 11294 -6717 11377 -6700
rect 11411 -6700 11427 -6683
rect 11619 -6683 11685 -6667
rect 11619 -6700 11635 -6683
rect 11411 -6717 11494 -6700
rect 11294 -6755 11494 -6717
rect 11552 -6717 11635 -6700
rect 11669 -6700 11685 -6683
rect 11877 -6683 11943 -6667
rect 11877 -6700 11893 -6683
rect 11669 -6717 11752 -6700
rect 11552 -6755 11752 -6717
rect 11810 -6717 11893 -6700
rect 11927 -6700 11943 -6683
rect 12135 -6683 12201 -6667
rect 12135 -6700 12151 -6683
rect 11927 -6717 12010 -6700
rect 11810 -6755 12010 -6717
rect 12068 -6717 12151 -6700
rect 12185 -6700 12201 -6683
rect 12393 -6683 12459 -6667
rect 12393 -6700 12409 -6683
rect 12185 -6717 12268 -6700
rect 12068 -6755 12268 -6717
rect 12326 -6717 12409 -6700
rect 12443 -6700 12459 -6683
rect 12443 -6717 12526 -6700
rect 12326 -6755 12526 -6717
rect 5187 -6994 5387 -6956
rect 5187 -7011 5270 -6994
rect 5254 -7028 5270 -7011
rect 5304 -7011 5387 -6994
rect 5445 -6994 5645 -6956
rect 5445 -7011 5528 -6994
rect 5304 -7028 5320 -7011
rect 5254 -7044 5320 -7028
rect 5512 -7028 5528 -7011
rect 5562 -7011 5645 -6994
rect 5703 -6994 5903 -6956
rect 5703 -7011 5786 -6994
rect 5562 -7028 5578 -7011
rect 5512 -7044 5578 -7028
rect 5770 -7028 5786 -7011
rect 5820 -7011 5903 -6994
rect 5961 -6994 6161 -6956
rect 5961 -7011 6044 -6994
rect 5820 -7028 5836 -7011
rect 5770 -7044 5836 -7028
rect 6028 -7028 6044 -7011
rect 6078 -7011 6161 -6994
rect 6219 -6994 6419 -6956
rect 6219 -7011 6302 -6994
rect 6078 -7028 6094 -7011
rect 6028 -7044 6094 -7028
rect 6286 -7028 6302 -7011
rect 6336 -7011 6419 -6994
rect 6477 -6994 6677 -6956
rect 6477 -7011 6560 -6994
rect 6336 -7028 6352 -7011
rect 6286 -7044 6352 -7028
rect 6544 -7028 6560 -7011
rect 6594 -7011 6677 -6994
rect 6735 -6994 6935 -6956
rect 6735 -7011 6818 -6994
rect 6594 -7028 6610 -7011
rect 6544 -7044 6610 -7028
rect 6802 -7028 6818 -7011
rect 6852 -7011 6935 -6994
rect 6993 -6994 7193 -6956
rect 6993 -7011 7076 -6994
rect 6852 -7028 6868 -7011
rect 6802 -7044 6868 -7028
rect 7060 -7028 7076 -7011
rect 7110 -7011 7193 -6994
rect 7857 -6994 8057 -6956
rect 7857 -7011 7940 -6994
rect 7110 -7028 7126 -7011
rect 7060 -7044 7126 -7028
rect 7924 -7028 7940 -7011
rect 7974 -7011 8057 -6994
rect 8115 -6994 8315 -6956
rect 8115 -7011 8198 -6994
rect 7974 -7028 7990 -7011
rect 7924 -7044 7990 -7028
rect 8182 -7028 8198 -7011
rect 8232 -7011 8315 -6994
rect 8373 -6994 8573 -6956
rect 8373 -7011 8456 -6994
rect 8232 -7028 8248 -7011
rect 8182 -7044 8248 -7028
rect 8440 -7028 8456 -7011
rect 8490 -7011 8573 -6994
rect 8631 -6994 8831 -6956
rect 8631 -7011 8714 -6994
rect 8490 -7028 8506 -7011
rect 8440 -7044 8506 -7028
rect 8698 -7028 8714 -7011
rect 8748 -7011 8831 -6994
rect 8889 -6994 9089 -6956
rect 8889 -7011 8972 -6994
rect 8748 -7028 8764 -7011
rect 8698 -7044 8764 -7028
rect 8956 -7028 8972 -7011
rect 9006 -7011 9089 -6994
rect 9147 -6994 9347 -6956
rect 9147 -7011 9230 -6994
rect 9006 -7028 9022 -7011
rect 8956 -7044 9022 -7028
rect 9214 -7028 9230 -7011
rect 9264 -7011 9347 -6994
rect 9405 -6994 9605 -6956
rect 9405 -7011 9488 -6994
rect 9264 -7028 9280 -7011
rect 9214 -7044 9280 -7028
rect 9472 -7028 9488 -7011
rect 9522 -7011 9605 -6994
rect 9663 -6994 9863 -6956
rect 9663 -7011 9746 -6994
rect 9522 -7028 9538 -7011
rect 9472 -7044 9538 -7028
rect 9730 -7028 9746 -7011
rect 9780 -7011 9863 -6994
rect 10520 -6993 10720 -6955
rect 10520 -7010 10603 -6993
rect 9780 -7028 9796 -7011
rect 9730 -7044 9796 -7028
rect 10587 -7027 10603 -7010
rect 10637 -7010 10720 -6993
rect 10778 -6993 10978 -6955
rect 10778 -7010 10861 -6993
rect 10637 -7027 10653 -7010
rect 10587 -7043 10653 -7027
rect 10845 -7027 10861 -7010
rect 10895 -7010 10978 -6993
rect 11036 -6993 11236 -6955
rect 11036 -7010 11119 -6993
rect 10895 -7027 10911 -7010
rect 10845 -7043 10911 -7027
rect 11103 -7027 11119 -7010
rect 11153 -7010 11236 -6993
rect 11294 -6993 11494 -6955
rect 11294 -7010 11377 -6993
rect 11153 -7027 11169 -7010
rect 11103 -7043 11169 -7027
rect 11361 -7027 11377 -7010
rect 11411 -7010 11494 -6993
rect 11552 -6993 11752 -6955
rect 11552 -7010 11635 -6993
rect 11411 -7027 11427 -7010
rect 11361 -7043 11427 -7027
rect 11619 -7027 11635 -7010
rect 11669 -7010 11752 -6993
rect 11810 -6993 12010 -6955
rect 11810 -7010 11893 -6993
rect 11669 -7027 11685 -7010
rect 11619 -7043 11685 -7027
rect 11877 -7027 11893 -7010
rect 11927 -7010 12010 -6993
rect 12068 -6993 12268 -6955
rect 12068 -7010 12151 -6993
rect 11927 -7027 11943 -7010
rect 11877 -7043 11943 -7027
rect 12135 -7027 12151 -7010
rect 12185 -7010 12268 -6993
rect 12326 -6993 12526 -6955
rect 12326 -7010 12409 -6993
rect 12185 -7027 12201 -7010
rect 12135 -7043 12201 -7027
rect 12393 -7027 12409 -7010
rect 12443 -7010 12526 -6993
rect 12443 -7027 12459 -7010
rect 12393 -7043 12459 -7027
rect 5254 -7102 5320 -7086
rect 5254 -7119 5270 -7102
rect 5187 -7136 5270 -7119
rect 5304 -7119 5320 -7102
rect 5512 -7102 5578 -7086
rect 5512 -7119 5528 -7102
rect 5304 -7136 5387 -7119
rect 5187 -7174 5387 -7136
rect 5445 -7136 5528 -7119
rect 5562 -7119 5578 -7102
rect 5770 -7102 5836 -7086
rect 5770 -7119 5786 -7102
rect 5562 -7136 5645 -7119
rect 5445 -7174 5645 -7136
rect 5703 -7136 5786 -7119
rect 5820 -7119 5836 -7102
rect 6028 -7102 6094 -7086
rect 6028 -7119 6044 -7102
rect 5820 -7136 5903 -7119
rect 5703 -7174 5903 -7136
rect 5961 -7136 6044 -7119
rect 6078 -7119 6094 -7102
rect 6286 -7102 6352 -7086
rect 6286 -7119 6302 -7102
rect 6078 -7136 6161 -7119
rect 5961 -7174 6161 -7136
rect 6219 -7136 6302 -7119
rect 6336 -7119 6352 -7102
rect 6544 -7102 6610 -7086
rect 6544 -7119 6560 -7102
rect 6336 -7136 6419 -7119
rect 6219 -7174 6419 -7136
rect 6477 -7136 6560 -7119
rect 6594 -7119 6610 -7102
rect 6802 -7102 6868 -7086
rect 6802 -7119 6818 -7102
rect 6594 -7136 6677 -7119
rect 6477 -7174 6677 -7136
rect 6735 -7136 6818 -7119
rect 6852 -7119 6868 -7102
rect 7060 -7102 7126 -7086
rect 7060 -7119 7076 -7102
rect 6852 -7136 6935 -7119
rect 6735 -7174 6935 -7136
rect 6993 -7136 7076 -7119
rect 7110 -7119 7126 -7102
rect 7924 -7102 7990 -7086
rect 7924 -7119 7940 -7102
rect 7110 -7136 7193 -7119
rect 6993 -7174 7193 -7136
rect 7857 -7136 7940 -7119
rect 7974 -7119 7990 -7102
rect 8182 -7102 8248 -7086
rect 8182 -7119 8198 -7102
rect 7974 -7136 8057 -7119
rect 7857 -7174 8057 -7136
rect 8115 -7136 8198 -7119
rect 8232 -7119 8248 -7102
rect 8440 -7102 8506 -7086
rect 8440 -7119 8456 -7102
rect 8232 -7136 8315 -7119
rect 8115 -7174 8315 -7136
rect 8373 -7136 8456 -7119
rect 8490 -7119 8506 -7102
rect 8698 -7102 8764 -7086
rect 8698 -7119 8714 -7102
rect 8490 -7136 8573 -7119
rect 8373 -7174 8573 -7136
rect 8631 -7136 8714 -7119
rect 8748 -7119 8764 -7102
rect 8956 -7102 9022 -7086
rect 8956 -7119 8972 -7102
rect 8748 -7136 8831 -7119
rect 8631 -7174 8831 -7136
rect 8889 -7136 8972 -7119
rect 9006 -7119 9022 -7102
rect 9214 -7102 9280 -7086
rect 9214 -7119 9230 -7102
rect 9006 -7136 9089 -7119
rect 8889 -7174 9089 -7136
rect 9147 -7136 9230 -7119
rect 9264 -7119 9280 -7102
rect 9472 -7102 9538 -7086
rect 9472 -7119 9488 -7102
rect 9264 -7136 9347 -7119
rect 9147 -7174 9347 -7136
rect 9405 -7136 9488 -7119
rect 9522 -7119 9538 -7102
rect 9730 -7102 9796 -7086
rect 9730 -7119 9746 -7102
rect 9522 -7136 9605 -7119
rect 9405 -7174 9605 -7136
rect 9663 -7136 9746 -7119
rect 9780 -7119 9796 -7102
rect 10587 -7101 10653 -7085
rect 10587 -7118 10603 -7101
rect 9780 -7136 9863 -7119
rect 9663 -7174 9863 -7136
rect 10520 -7135 10603 -7118
rect 10637 -7118 10653 -7101
rect 10845 -7101 10911 -7085
rect 10845 -7118 10861 -7101
rect 10637 -7135 10720 -7118
rect 10520 -7173 10720 -7135
rect 10778 -7135 10861 -7118
rect 10895 -7118 10911 -7101
rect 11103 -7101 11169 -7085
rect 11103 -7118 11119 -7101
rect 10895 -7135 10978 -7118
rect 10778 -7173 10978 -7135
rect 11036 -7135 11119 -7118
rect 11153 -7118 11169 -7101
rect 11361 -7101 11427 -7085
rect 11361 -7118 11377 -7101
rect 11153 -7135 11236 -7118
rect 11036 -7173 11236 -7135
rect 11294 -7135 11377 -7118
rect 11411 -7118 11427 -7101
rect 11619 -7101 11685 -7085
rect 11619 -7118 11635 -7101
rect 11411 -7135 11494 -7118
rect 11294 -7173 11494 -7135
rect 11552 -7135 11635 -7118
rect 11669 -7118 11685 -7101
rect 11877 -7101 11943 -7085
rect 11877 -7118 11893 -7101
rect 11669 -7135 11752 -7118
rect 11552 -7173 11752 -7135
rect 11810 -7135 11893 -7118
rect 11927 -7118 11943 -7101
rect 12135 -7101 12201 -7085
rect 12135 -7118 12151 -7101
rect 11927 -7135 12010 -7118
rect 11810 -7173 12010 -7135
rect 12068 -7135 12151 -7118
rect 12185 -7118 12201 -7101
rect 12393 -7101 12459 -7085
rect 12393 -7118 12409 -7101
rect 12185 -7135 12268 -7118
rect 12068 -7173 12268 -7135
rect 12326 -7135 12409 -7118
rect 12443 -7118 12459 -7101
rect 12443 -7135 12526 -7118
rect 12326 -7173 12526 -7135
rect 5187 -7412 5387 -7374
rect 5187 -7429 5270 -7412
rect 5254 -7446 5270 -7429
rect 5304 -7429 5387 -7412
rect 5445 -7412 5645 -7374
rect 5445 -7429 5528 -7412
rect 5304 -7446 5320 -7429
rect 5254 -7462 5320 -7446
rect 5512 -7446 5528 -7429
rect 5562 -7429 5645 -7412
rect 5703 -7412 5903 -7374
rect 5703 -7429 5786 -7412
rect 5562 -7446 5578 -7429
rect 5512 -7462 5578 -7446
rect 5770 -7446 5786 -7429
rect 5820 -7429 5903 -7412
rect 5961 -7412 6161 -7374
rect 5961 -7429 6044 -7412
rect 5820 -7446 5836 -7429
rect 5770 -7462 5836 -7446
rect 6028 -7446 6044 -7429
rect 6078 -7429 6161 -7412
rect 6219 -7412 6419 -7374
rect 6219 -7429 6302 -7412
rect 6078 -7446 6094 -7429
rect 6028 -7462 6094 -7446
rect 6286 -7446 6302 -7429
rect 6336 -7429 6419 -7412
rect 6477 -7412 6677 -7374
rect 6477 -7429 6560 -7412
rect 6336 -7446 6352 -7429
rect 6286 -7462 6352 -7446
rect 6544 -7446 6560 -7429
rect 6594 -7429 6677 -7412
rect 6735 -7412 6935 -7374
rect 6735 -7429 6818 -7412
rect 6594 -7446 6610 -7429
rect 6544 -7462 6610 -7446
rect 6802 -7446 6818 -7429
rect 6852 -7429 6935 -7412
rect 6993 -7412 7193 -7374
rect 6993 -7429 7076 -7412
rect 6852 -7446 6868 -7429
rect 6802 -7462 6868 -7446
rect 7060 -7446 7076 -7429
rect 7110 -7429 7193 -7412
rect 7857 -7412 8057 -7374
rect 7857 -7429 7940 -7412
rect 7110 -7446 7126 -7429
rect 7060 -7462 7126 -7446
rect 7924 -7446 7940 -7429
rect 7974 -7429 8057 -7412
rect 8115 -7412 8315 -7374
rect 8115 -7429 8198 -7412
rect 7974 -7446 7990 -7429
rect 7924 -7462 7990 -7446
rect 8182 -7446 8198 -7429
rect 8232 -7429 8315 -7412
rect 8373 -7412 8573 -7374
rect 8373 -7429 8456 -7412
rect 8232 -7446 8248 -7429
rect 8182 -7462 8248 -7446
rect 8440 -7446 8456 -7429
rect 8490 -7429 8573 -7412
rect 8631 -7412 8831 -7374
rect 8631 -7429 8714 -7412
rect 8490 -7446 8506 -7429
rect 8440 -7462 8506 -7446
rect 8698 -7446 8714 -7429
rect 8748 -7429 8831 -7412
rect 8889 -7412 9089 -7374
rect 8889 -7429 8972 -7412
rect 8748 -7446 8764 -7429
rect 8698 -7462 8764 -7446
rect 8956 -7446 8972 -7429
rect 9006 -7429 9089 -7412
rect 9147 -7412 9347 -7374
rect 9147 -7429 9230 -7412
rect 9006 -7446 9022 -7429
rect 8956 -7462 9022 -7446
rect 9214 -7446 9230 -7429
rect 9264 -7429 9347 -7412
rect 9405 -7412 9605 -7374
rect 9405 -7429 9488 -7412
rect 9264 -7446 9280 -7429
rect 9214 -7462 9280 -7446
rect 9472 -7446 9488 -7429
rect 9522 -7429 9605 -7412
rect 9663 -7412 9863 -7374
rect 9663 -7429 9746 -7412
rect 9522 -7446 9538 -7429
rect 9472 -7462 9538 -7446
rect 9730 -7446 9746 -7429
rect 9780 -7429 9863 -7412
rect 10520 -7411 10720 -7373
rect 10520 -7428 10603 -7411
rect 9780 -7446 9796 -7429
rect 9730 -7462 9796 -7446
rect 10587 -7445 10603 -7428
rect 10637 -7428 10720 -7411
rect 10778 -7411 10978 -7373
rect 10778 -7428 10861 -7411
rect 10637 -7445 10653 -7428
rect 10587 -7461 10653 -7445
rect 10845 -7445 10861 -7428
rect 10895 -7428 10978 -7411
rect 11036 -7411 11236 -7373
rect 11036 -7428 11119 -7411
rect 10895 -7445 10911 -7428
rect 10845 -7461 10911 -7445
rect 11103 -7445 11119 -7428
rect 11153 -7428 11236 -7411
rect 11294 -7411 11494 -7373
rect 11294 -7428 11377 -7411
rect 11153 -7445 11169 -7428
rect 11103 -7461 11169 -7445
rect 11361 -7445 11377 -7428
rect 11411 -7428 11494 -7411
rect 11552 -7411 11752 -7373
rect 11552 -7428 11635 -7411
rect 11411 -7445 11427 -7428
rect 11361 -7461 11427 -7445
rect 11619 -7445 11635 -7428
rect 11669 -7428 11752 -7411
rect 11810 -7411 12010 -7373
rect 11810 -7428 11893 -7411
rect 11669 -7445 11685 -7428
rect 11619 -7461 11685 -7445
rect 11877 -7445 11893 -7428
rect 11927 -7428 12010 -7411
rect 12068 -7411 12268 -7373
rect 12068 -7428 12151 -7411
rect 11927 -7445 11943 -7428
rect 11877 -7461 11943 -7445
rect 12135 -7445 12151 -7428
rect 12185 -7428 12268 -7411
rect 12326 -7411 12526 -7373
rect 12326 -7428 12409 -7411
rect 12185 -7445 12201 -7428
rect 12135 -7461 12201 -7445
rect 12393 -7445 12409 -7428
rect 12443 -7428 12526 -7411
rect 12443 -7445 12459 -7428
rect 12393 -7461 12459 -7445
rect 5254 -7520 5320 -7504
rect 5254 -7537 5270 -7520
rect 5187 -7554 5270 -7537
rect 5304 -7537 5320 -7520
rect 5512 -7520 5578 -7504
rect 5512 -7537 5528 -7520
rect 5304 -7554 5387 -7537
rect 5187 -7592 5387 -7554
rect 5445 -7554 5528 -7537
rect 5562 -7537 5578 -7520
rect 5770 -7520 5836 -7504
rect 5770 -7537 5786 -7520
rect 5562 -7554 5645 -7537
rect 5445 -7592 5645 -7554
rect 5703 -7554 5786 -7537
rect 5820 -7537 5836 -7520
rect 6028 -7520 6094 -7504
rect 6028 -7537 6044 -7520
rect 5820 -7554 5903 -7537
rect 5703 -7592 5903 -7554
rect 5961 -7554 6044 -7537
rect 6078 -7537 6094 -7520
rect 6286 -7520 6352 -7504
rect 6286 -7537 6302 -7520
rect 6078 -7554 6161 -7537
rect 5961 -7592 6161 -7554
rect 6219 -7554 6302 -7537
rect 6336 -7537 6352 -7520
rect 6544 -7520 6610 -7504
rect 6544 -7537 6560 -7520
rect 6336 -7554 6419 -7537
rect 6219 -7592 6419 -7554
rect 6477 -7554 6560 -7537
rect 6594 -7537 6610 -7520
rect 6802 -7520 6868 -7504
rect 6802 -7537 6818 -7520
rect 6594 -7554 6677 -7537
rect 6477 -7592 6677 -7554
rect 6735 -7554 6818 -7537
rect 6852 -7537 6868 -7520
rect 7060 -7520 7126 -7504
rect 7060 -7537 7076 -7520
rect 6852 -7554 6935 -7537
rect 6735 -7592 6935 -7554
rect 6993 -7554 7076 -7537
rect 7110 -7537 7126 -7520
rect 7924 -7520 7990 -7504
rect 7924 -7537 7940 -7520
rect 7110 -7554 7193 -7537
rect 6993 -7592 7193 -7554
rect 7857 -7554 7940 -7537
rect 7974 -7537 7990 -7520
rect 8182 -7520 8248 -7504
rect 8182 -7537 8198 -7520
rect 7974 -7554 8057 -7537
rect 7857 -7592 8057 -7554
rect 8115 -7554 8198 -7537
rect 8232 -7537 8248 -7520
rect 8440 -7520 8506 -7504
rect 8440 -7537 8456 -7520
rect 8232 -7554 8315 -7537
rect 8115 -7592 8315 -7554
rect 8373 -7554 8456 -7537
rect 8490 -7537 8506 -7520
rect 8698 -7520 8764 -7504
rect 8698 -7537 8714 -7520
rect 8490 -7554 8573 -7537
rect 8373 -7592 8573 -7554
rect 8631 -7554 8714 -7537
rect 8748 -7537 8764 -7520
rect 8956 -7520 9022 -7504
rect 8956 -7537 8972 -7520
rect 8748 -7554 8831 -7537
rect 8631 -7592 8831 -7554
rect 8889 -7554 8972 -7537
rect 9006 -7537 9022 -7520
rect 9214 -7520 9280 -7504
rect 9214 -7537 9230 -7520
rect 9006 -7554 9089 -7537
rect 8889 -7592 9089 -7554
rect 9147 -7554 9230 -7537
rect 9264 -7537 9280 -7520
rect 9472 -7520 9538 -7504
rect 9472 -7537 9488 -7520
rect 9264 -7554 9347 -7537
rect 9147 -7592 9347 -7554
rect 9405 -7554 9488 -7537
rect 9522 -7537 9538 -7520
rect 9730 -7520 9796 -7504
rect 9730 -7537 9746 -7520
rect 9522 -7554 9605 -7537
rect 9405 -7592 9605 -7554
rect 9663 -7554 9746 -7537
rect 9780 -7537 9796 -7520
rect 10587 -7519 10653 -7503
rect 10587 -7536 10603 -7519
rect 9780 -7554 9863 -7537
rect 9663 -7592 9863 -7554
rect 10520 -7553 10603 -7536
rect 10637 -7536 10653 -7519
rect 10845 -7519 10911 -7503
rect 10845 -7536 10861 -7519
rect 10637 -7553 10720 -7536
rect 10520 -7591 10720 -7553
rect 10778 -7553 10861 -7536
rect 10895 -7536 10911 -7519
rect 11103 -7519 11169 -7503
rect 11103 -7536 11119 -7519
rect 10895 -7553 10978 -7536
rect 10778 -7591 10978 -7553
rect 11036 -7553 11119 -7536
rect 11153 -7536 11169 -7519
rect 11361 -7519 11427 -7503
rect 11361 -7536 11377 -7519
rect 11153 -7553 11236 -7536
rect 11036 -7591 11236 -7553
rect 11294 -7553 11377 -7536
rect 11411 -7536 11427 -7519
rect 11619 -7519 11685 -7503
rect 11619 -7536 11635 -7519
rect 11411 -7553 11494 -7536
rect 11294 -7591 11494 -7553
rect 11552 -7553 11635 -7536
rect 11669 -7536 11685 -7519
rect 11877 -7519 11943 -7503
rect 11877 -7536 11893 -7519
rect 11669 -7553 11752 -7536
rect 11552 -7591 11752 -7553
rect 11810 -7553 11893 -7536
rect 11927 -7536 11943 -7519
rect 12135 -7519 12201 -7503
rect 12135 -7536 12151 -7519
rect 11927 -7553 12010 -7536
rect 11810 -7591 12010 -7553
rect 12068 -7553 12151 -7536
rect 12185 -7536 12201 -7519
rect 12393 -7519 12459 -7503
rect 12393 -7536 12409 -7519
rect 12185 -7553 12268 -7536
rect 12068 -7591 12268 -7553
rect 12326 -7553 12409 -7536
rect 12443 -7536 12459 -7519
rect 12443 -7553 12526 -7536
rect 12326 -7591 12526 -7553
rect 5187 -7830 5387 -7792
rect 5187 -7847 5270 -7830
rect 5254 -7864 5270 -7847
rect 5304 -7847 5387 -7830
rect 5445 -7830 5645 -7792
rect 5445 -7847 5528 -7830
rect 5304 -7864 5320 -7847
rect 5254 -7880 5320 -7864
rect 5512 -7864 5528 -7847
rect 5562 -7847 5645 -7830
rect 5703 -7830 5903 -7792
rect 5703 -7847 5786 -7830
rect 5562 -7864 5578 -7847
rect 5512 -7880 5578 -7864
rect 5770 -7864 5786 -7847
rect 5820 -7847 5903 -7830
rect 5961 -7830 6161 -7792
rect 5961 -7847 6044 -7830
rect 5820 -7864 5836 -7847
rect 5770 -7880 5836 -7864
rect 6028 -7864 6044 -7847
rect 6078 -7847 6161 -7830
rect 6219 -7830 6419 -7792
rect 6219 -7847 6302 -7830
rect 6078 -7864 6094 -7847
rect 6028 -7880 6094 -7864
rect 6286 -7864 6302 -7847
rect 6336 -7847 6419 -7830
rect 6477 -7830 6677 -7792
rect 6477 -7847 6560 -7830
rect 6336 -7864 6352 -7847
rect 6286 -7880 6352 -7864
rect 6544 -7864 6560 -7847
rect 6594 -7847 6677 -7830
rect 6735 -7830 6935 -7792
rect 6735 -7847 6818 -7830
rect 6594 -7864 6610 -7847
rect 6544 -7880 6610 -7864
rect 6802 -7864 6818 -7847
rect 6852 -7847 6935 -7830
rect 6993 -7830 7193 -7792
rect 6993 -7847 7076 -7830
rect 6852 -7864 6868 -7847
rect 6802 -7880 6868 -7864
rect 7060 -7864 7076 -7847
rect 7110 -7847 7193 -7830
rect 7857 -7830 8057 -7792
rect 7857 -7847 7940 -7830
rect 7110 -7864 7126 -7847
rect 7060 -7880 7126 -7864
rect 7924 -7864 7940 -7847
rect 7974 -7847 8057 -7830
rect 8115 -7830 8315 -7792
rect 8115 -7847 8198 -7830
rect 7974 -7864 7990 -7847
rect 7924 -7880 7990 -7864
rect 8182 -7864 8198 -7847
rect 8232 -7847 8315 -7830
rect 8373 -7830 8573 -7792
rect 8373 -7847 8456 -7830
rect 8232 -7864 8248 -7847
rect 8182 -7880 8248 -7864
rect 8440 -7864 8456 -7847
rect 8490 -7847 8573 -7830
rect 8631 -7830 8831 -7792
rect 8631 -7847 8714 -7830
rect 8490 -7864 8506 -7847
rect 8440 -7880 8506 -7864
rect 8698 -7864 8714 -7847
rect 8748 -7847 8831 -7830
rect 8889 -7830 9089 -7792
rect 8889 -7847 8972 -7830
rect 8748 -7864 8764 -7847
rect 8698 -7880 8764 -7864
rect 8956 -7864 8972 -7847
rect 9006 -7847 9089 -7830
rect 9147 -7830 9347 -7792
rect 9147 -7847 9230 -7830
rect 9006 -7864 9022 -7847
rect 8956 -7880 9022 -7864
rect 9214 -7864 9230 -7847
rect 9264 -7847 9347 -7830
rect 9405 -7830 9605 -7792
rect 9405 -7847 9488 -7830
rect 9264 -7864 9280 -7847
rect 9214 -7880 9280 -7864
rect 9472 -7864 9488 -7847
rect 9522 -7847 9605 -7830
rect 9663 -7830 9863 -7792
rect 9663 -7847 9746 -7830
rect 9522 -7864 9538 -7847
rect 9472 -7880 9538 -7864
rect 9730 -7864 9746 -7847
rect 9780 -7847 9863 -7830
rect 10520 -7829 10720 -7791
rect 10520 -7846 10603 -7829
rect 9780 -7864 9796 -7847
rect 9730 -7880 9796 -7864
rect 10587 -7863 10603 -7846
rect 10637 -7846 10720 -7829
rect 10778 -7829 10978 -7791
rect 10778 -7846 10861 -7829
rect 10637 -7863 10653 -7846
rect 10587 -7879 10653 -7863
rect 10845 -7863 10861 -7846
rect 10895 -7846 10978 -7829
rect 11036 -7829 11236 -7791
rect 11036 -7846 11119 -7829
rect 10895 -7863 10911 -7846
rect 10845 -7879 10911 -7863
rect 11103 -7863 11119 -7846
rect 11153 -7846 11236 -7829
rect 11294 -7829 11494 -7791
rect 11294 -7846 11377 -7829
rect 11153 -7863 11169 -7846
rect 11103 -7879 11169 -7863
rect 11361 -7863 11377 -7846
rect 11411 -7846 11494 -7829
rect 11552 -7829 11752 -7791
rect 11552 -7846 11635 -7829
rect 11411 -7863 11427 -7846
rect 11361 -7879 11427 -7863
rect 11619 -7863 11635 -7846
rect 11669 -7846 11752 -7829
rect 11810 -7829 12010 -7791
rect 11810 -7846 11893 -7829
rect 11669 -7863 11685 -7846
rect 11619 -7879 11685 -7863
rect 11877 -7863 11893 -7846
rect 11927 -7846 12010 -7829
rect 12068 -7829 12268 -7791
rect 12068 -7846 12151 -7829
rect 11927 -7863 11943 -7846
rect 11877 -7879 11943 -7863
rect 12135 -7863 12151 -7846
rect 12185 -7846 12268 -7829
rect 12326 -7829 12526 -7791
rect 12326 -7846 12409 -7829
rect 12185 -7863 12201 -7846
rect 12135 -7879 12201 -7863
rect 12393 -7863 12409 -7846
rect 12443 -7846 12526 -7829
rect 12443 -7863 12459 -7846
rect 12393 -7879 12459 -7863
rect 5134 -8172 5200 -8156
rect 5134 -8189 5150 -8172
rect 5067 -8206 5150 -8189
rect 5184 -8189 5200 -8172
rect 5674 -8172 5740 -8156
rect 5674 -8189 5690 -8172
rect 5184 -8206 5267 -8189
rect 5067 -8244 5267 -8206
rect 5607 -8206 5690 -8189
rect 5724 -8189 5740 -8172
rect 6154 -8172 6220 -8156
rect 6154 -8189 6170 -8172
rect 5724 -8206 5807 -8189
rect 5607 -8244 5807 -8206
rect 6087 -8206 6170 -8189
rect 6204 -8189 6220 -8172
rect 6657 -8170 6723 -8154
rect 6657 -8187 6673 -8170
rect 6204 -8206 6287 -8189
rect 6087 -8244 6287 -8206
rect 6590 -8204 6673 -8187
rect 6707 -8187 6723 -8170
rect 7167 -8160 7233 -8144
rect 7167 -8177 7183 -8160
rect 6707 -8204 6790 -8187
rect 6590 -8242 6790 -8204
rect 7100 -8194 7183 -8177
rect 7217 -8177 7233 -8160
rect 7804 -8172 7870 -8156
rect 7217 -8194 7300 -8177
rect 7804 -8189 7820 -8172
rect 7100 -8232 7300 -8194
rect 7737 -8206 7820 -8189
rect 7854 -8189 7870 -8172
rect 8344 -8172 8410 -8156
rect 8344 -8189 8360 -8172
rect 7854 -8206 7937 -8189
rect 7737 -8244 7937 -8206
rect 8277 -8206 8360 -8189
rect 8394 -8189 8410 -8172
rect 8824 -8172 8890 -8156
rect 8824 -8189 8840 -8172
rect 8394 -8206 8477 -8189
rect 8277 -8244 8477 -8206
rect 8757 -8206 8840 -8189
rect 8874 -8189 8890 -8172
rect 9327 -8170 9393 -8154
rect 9327 -8187 9343 -8170
rect 8874 -8206 8957 -8189
rect 8757 -8244 8957 -8206
rect 9260 -8204 9343 -8187
rect 9377 -8187 9393 -8170
rect 9837 -8160 9903 -8144
rect 9837 -8177 9853 -8160
rect 9377 -8204 9460 -8187
rect 9260 -8242 9460 -8204
rect 9770 -8194 9853 -8177
rect 9887 -8177 9903 -8160
rect 10467 -8171 10533 -8155
rect 9887 -8194 9970 -8177
rect 10467 -8188 10483 -8171
rect 9770 -8232 9970 -8194
rect 10400 -8205 10483 -8188
rect 10517 -8188 10533 -8171
rect 11007 -8171 11073 -8155
rect 11007 -8188 11023 -8171
rect 10517 -8205 10600 -8188
rect 5067 -8482 5267 -8444
rect 5067 -8499 5150 -8482
rect 5134 -8516 5150 -8499
rect 5184 -8499 5267 -8482
rect 5607 -8482 5807 -8444
rect 5607 -8499 5690 -8482
rect 5184 -8516 5200 -8499
rect 5134 -8532 5200 -8516
rect 5674 -8516 5690 -8499
rect 5724 -8499 5807 -8482
rect 6087 -8482 6287 -8444
rect 6087 -8499 6170 -8482
rect 5724 -8516 5740 -8499
rect 5674 -8532 5740 -8516
rect 6154 -8516 6170 -8499
rect 6204 -8499 6287 -8482
rect 6590 -8480 6790 -8442
rect 6590 -8497 6673 -8480
rect 6204 -8516 6220 -8499
rect 6154 -8532 6220 -8516
rect 6657 -8514 6673 -8497
rect 6707 -8497 6790 -8480
rect 7100 -8470 7300 -8432
rect 10400 -8243 10600 -8205
rect 10940 -8205 11023 -8188
rect 11057 -8188 11073 -8171
rect 11487 -8171 11553 -8155
rect 11487 -8188 11503 -8171
rect 11057 -8205 11140 -8188
rect 10940 -8243 11140 -8205
rect 11420 -8205 11503 -8188
rect 11537 -8188 11553 -8171
rect 11990 -8169 12056 -8153
rect 11990 -8186 12006 -8169
rect 11537 -8205 11620 -8188
rect 11420 -8243 11620 -8205
rect 11923 -8203 12006 -8186
rect 12040 -8186 12056 -8169
rect 12500 -8159 12566 -8143
rect 12500 -8176 12516 -8159
rect 12040 -8203 12123 -8186
rect 11923 -8241 12123 -8203
rect 12433 -8193 12516 -8176
rect 12550 -8176 12566 -8159
rect 12550 -8193 12633 -8176
rect 12433 -8231 12633 -8193
rect 7100 -8487 7183 -8470
rect 6707 -8514 6723 -8497
rect 6657 -8530 6723 -8514
rect 7167 -8504 7183 -8487
rect 7217 -8487 7300 -8470
rect 7737 -8482 7937 -8444
rect 7217 -8504 7233 -8487
rect 7737 -8499 7820 -8482
rect 7167 -8520 7233 -8504
rect 7804 -8516 7820 -8499
rect 7854 -8499 7937 -8482
rect 8277 -8482 8477 -8444
rect 8277 -8499 8360 -8482
rect 7854 -8516 7870 -8499
rect 7804 -8532 7870 -8516
rect 8344 -8516 8360 -8499
rect 8394 -8499 8477 -8482
rect 8757 -8482 8957 -8444
rect 8757 -8499 8840 -8482
rect 8394 -8516 8410 -8499
rect 8344 -8532 8410 -8516
rect 8824 -8516 8840 -8499
rect 8874 -8499 8957 -8482
rect 9260 -8480 9460 -8442
rect 9260 -8497 9343 -8480
rect 8874 -8516 8890 -8499
rect 8824 -8532 8890 -8516
rect 9327 -8514 9343 -8497
rect 9377 -8497 9460 -8480
rect 9770 -8470 9970 -8432
rect 9770 -8487 9853 -8470
rect 9377 -8514 9393 -8497
rect 9327 -8530 9393 -8514
rect 9837 -8504 9853 -8487
rect 9887 -8487 9970 -8470
rect 10400 -8481 10600 -8443
rect 9887 -8504 9903 -8487
rect 10400 -8498 10483 -8481
rect 9837 -8520 9903 -8504
rect 10467 -8515 10483 -8498
rect 10517 -8498 10600 -8481
rect 10940 -8481 11140 -8443
rect 10940 -8498 11023 -8481
rect 10517 -8515 10533 -8498
rect 10467 -8531 10533 -8515
rect 11007 -8515 11023 -8498
rect 11057 -8498 11140 -8481
rect 11420 -8481 11620 -8443
rect 11420 -8498 11503 -8481
rect 11057 -8515 11073 -8498
rect 11007 -8531 11073 -8515
rect 11487 -8515 11503 -8498
rect 11537 -8498 11620 -8481
rect 11923 -8479 12123 -8441
rect 11923 -8496 12006 -8479
rect 11537 -8515 11553 -8498
rect 11487 -8531 11553 -8515
rect 11990 -8513 12006 -8496
rect 12040 -8496 12123 -8479
rect 12433 -8469 12633 -8431
rect 12433 -8486 12516 -8469
rect 12040 -8513 12056 -8496
rect 11990 -8529 12056 -8513
rect 12500 -8503 12516 -8486
rect 12550 -8486 12633 -8469
rect 12550 -8503 12566 -8486
rect 12500 -8519 12566 -8503
rect 14064 8623 15664 8639
rect 14064 8589 14080 8623
rect 15448 8589 15664 8623
rect 14064 8551 15664 8589
rect 15722 8623 17322 8639
rect 15722 8589 15941 8623
rect 17306 8589 17322 8623
rect 15722 8551 17322 8589
rect 14064 7113 15664 7151
rect 14064 7079 14080 7113
rect 15448 7079 15664 7113
rect 14064 7041 15664 7079
rect 15722 7113 17322 7151
rect 15722 7079 15941 7113
rect 17306 7079 17322 7113
rect 15722 7041 17322 7079
rect 14064 5603 15664 5641
rect 14064 5569 14080 5603
rect 15448 5569 15664 5603
rect 14064 5531 15664 5569
rect 15722 5603 17322 5641
rect 15722 5569 15941 5603
rect 17306 5569 17322 5603
rect 15722 5531 17322 5569
rect 14064 4093 15664 4131
rect 14064 4059 14080 4093
rect 15448 4059 15664 4093
rect 14064 4021 15664 4059
rect 15722 4093 17322 4131
rect 15722 4059 15941 4093
rect 17306 4059 17322 4093
rect 15722 4021 17322 4059
rect 14064 2583 15664 2621
rect 14064 2549 14080 2583
rect 15448 2549 15664 2583
rect 14064 2511 15664 2549
rect 15722 2583 17322 2621
rect 15722 2549 15941 2583
rect 17306 2549 17322 2583
rect 15722 2511 17322 2549
rect 14064 1073 15664 1111
rect 14064 1039 14080 1073
rect 15448 1039 15664 1073
rect 14064 1001 15664 1039
rect 15722 1073 17322 1111
rect 15722 1039 15941 1073
rect 17306 1039 17322 1073
rect 15722 1001 17322 1039
rect 14064 -437 15664 -399
rect 14064 -471 14080 -437
rect 15448 -471 15664 -437
rect 14064 -509 15664 -471
rect 15722 -437 17322 -399
rect 15722 -471 15941 -437
rect 17306 -471 17322 -437
rect 15722 -509 17322 -471
rect 14064 -1947 15664 -1909
rect 14064 -1981 14080 -1947
rect 15448 -1981 15664 -1947
rect 14064 -2019 15664 -1981
rect 15722 -1947 17322 -1909
rect 15722 -1981 15941 -1947
rect 17306 -1981 17322 -1947
rect 15722 -2019 17322 -1981
rect 14064 -3457 15664 -3419
rect 14064 -3491 14080 -3457
rect 15448 -3491 15664 -3457
rect 14064 -3529 15664 -3491
rect 15722 -3457 17322 -3419
rect 15722 -3491 15941 -3457
rect 17306 -3491 17322 -3457
rect 15722 -3529 17322 -3491
rect 14064 -4967 15664 -4929
rect 14064 -5001 14080 -4967
rect 15448 -5001 15664 -4967
rect 14064 -5039 15664 -5001
rect 15722 -4967 17322 -4929
rect 15722 -5001 15941 -4967
rect 17306 -5001 17322 -4967
rect 15722 -5039 17322 -5001
rect 14064 -6477 15664 -6439
rect 14064 -6511 14080 -6477
rect 15448 -6511 15664 -6477
rect 14064 -6549 15664 -6511
rect 15722 -6477 17322 -6439
rect 15722 -6511 15941 -6477
rect 17306 -6511 17322 -6477
rect 15722 -6549 17322 -6511
rect 14064 -7987 15664 -7949
rect 14064 -8021 14080 -7987
rect 15448 -8021 15664 -7987
rect 14064 -8059 15664 -8021
rect 15722 -7987 17322 -7949
rect 15722 -8021 15941 -7987
rect 17306 -8021 17322 -7987
rect 15722 -8059 17322 -8021
rect 14064 -9497 15664 -9459
rect 14064 -9531 14080 -9497
rect 15448 -9531 15664 -9497
rect 14064 -9547 15664 -9531
rect 15722 -9497 17322 -9459
rect 15722 -9531 15941 -9497
rect 17306 -9531 17322 -9497
rect 15722 -9547 17322 -9531
<< polycont >>
rect 459 8588 1824 8622
rect 2318 8588 3685 8622
rect 459 7078 1824 7112
rect 2318 7078 3685 7112
rect 459 5568 1824 5602
rect 2318 5568 3685 5602
rect 459 4058 1824 4092
rect 2318 4058 3685 4092
rect 459 2548 1824 2582
rect 2318 2548 3685 2582
rect 459 1038 1824 1072
rect 2318 1038 3685 1072
rect 459 -472 1824 -438
rect 2318 -472 3685 -438
rect 459 -1982 1824 -1948
rect 2318 -1982 3685 -1948
rect 459 -3492 1824 -3458
rect 2318 -3492 3685 -3458
rect 459 -5002 1824 -4968
rect 2318 -5002 3685 -4968
rect 459 -6512 1824 -6478
rect 2318 -6512 3685 -6478
rect 459 -8022 1824 -7988
rect 2318 -8022 3685 -7988
rect 459 -9532 1824 -9498
rect 2318 -9532 3685 -9498
rect 5544 8545 5578 8579
rect 6204 8545 6238 8579
rect 6674 8545 6708 8579
rect 7277 8544 7311 8578
rect 7535 8544 7569 8578
rect 7793 8544 7827 8578
rect 8051 8544 8085 8578
rect 8309 8544 8343 8578
rect 9092 8544 9126 8578
rect 9350 8544 9384 8578
rect 9608 8544 9642 8578
rect 9866 8544 9900 8578
rect 10124 8544 10158 8578
rect 10898 8544 10932 8578
rect 11156 8544 11190 8578
rect 11414 8544 11448 8578
rect 11672 8544 11706 8578
rect 11930 8544 11964 8578
rect 5544 8217 5578 8251
rect 6204 8217 6238 8251
rect 6674 8217 6708 8251
rect 7277 8216 7311 8250
rect 7535 8216 7569 8250
rect 7793 8216 7827 8250
rect 8051 8216 8085 8250
rect 8309 8216 8343 8250
rect 9092 8216 9126 8250
rect 9350 8216 9384 8250
rect 9608 8216 9642 8250
rect 9866 8216 9900 8250
rect 10124 8216 10158 8250
rect 10898 8216 10932 8250
rect 11156 8216 11190 8250
rect 11414 8216 11448 8250
rect 11672 8216 11706 8250
rect 11930 8216 11964 8250
rect 5436 7574 5502 7612
rect 6088 7571 6242 7605
rect 6822 7574 6888 7612
rect 7192 7574 7258 7612
rect 7614 7574 7680 7612
rect 8036 7574 8102 7612
rect 8758 7571 8912 7605
rect 9536 7574 9602 7612
rect 9906 7574 9972 7612
rect 10328 7574 10394 7612
rect 10750 7574 10816 7612
rect 11421 7572 11575 7606
rect 12190 7574 12256 7612
rect 6088 7333 6242 7367
rect 8758 7333 8912 7367
rect 11421 7334 11575 7368
rect 5270 6575 5304 6609
rect 5528 6575 5562 6609
rect 5786 6575 5820 6609
rect 6044 6575 6078 6609
rect 6302 6575 6336 6609
rect 6560 6575 6594 6609
rect 6818 6575 6852 6609
rect 7076 6575 7110 6609
rect 7940 6575 7974 6609
rect 8198 6575 8232 6609
rect 8456 6575 8490 6609
rect 8714 6575 8748 6609
rect 8972 6575 9006 6609
rect 9230 6575 9264 6609
rect 9488 6575 9522 6609
rect 9746 6575 9780 6609
rect 10603 6576 10637 6610
rect 10861 6576 10895 6610
rect 11119 6576 11153 6610
rect 11377 6576 11411 6610
rect 11635 6576 11669 6610
rect 11893 6576 11927 6610
rect 12151 6576 12185 6610
rect 12409 6576 12443 6610
rect 5270 6265 5304 6299
rect 5528 6265 5562 6299
rect 5786 6265 5820 6299
rect 6044 6265 6078 6299
rect 6302 6265 6336 6299
rect 6560 6265 6594 6299
rect 6818 6265 6852 6299
rect 7076 6265 7110 6299
rect 7940 6265 7974 6299
rect 8198 6265 8232 6299
rect 8456 6265 8490 6299
rect 8714 6265 8748 6299
rect 8972 6265 9006 6299
rect 9230 6265 9264 6299
rect 9488 6265 9522 6299
rect 9746 6265 9780 6299
rect 10603 6266 10637 6300
rect 10861 6266 10895 6300
rect 11119 6266 11153 6300
rect 11377 6266 11411 6300
rect 11635 6266 11669 6300
rect 11893 6266 11927 6300
rect 12151 6266 12185 6300
rect 12409 6266 12443 6300
rect 5270 6157 5304 6191
rect 5528 6157 5562 6191
rect 5786 6157 5820 6191
rect 6044 6157 6078 6191
rect 6302 6157 6336 6191
rect 6560 6157 6594 6191
rect 6818 6157 6852 6191
rect 7076 6157 7110 6191
rect 7940 6157 7974 6191
rect 8198 6157 8232 6191
rect 8456 6157 8490 6191
rect 8714 6157 8748 6191
rect 8972 6157 9006 6191
rect 9230 6157 9264 6191
rect 9488 6157 9522 6191
rect 9746 6157 9780 6191
rect 10603 6158 10637 6192
rect 10861 6158 10895 6192
rect 11119 6158 11153 6192
rect 11377 6158 11411 6192
rect 11635 6158 11669 6192
rect 11893 6158 11927 6192
rect 12151 6158 12185 6192
rect 12409 6158 12443 6192
rect 5270 5847 5304 5881
rect 5528 5847 5562 5881
rect 5786 5847 5820 5881
rect 6044 5847 6078 5881
rect 6302 5847 6336 5881
rect 6560 5847 6594 5881
rect 6818 5847 6852 5881
rect 7076 5847 7110 5881
rect 7940 5847 7974 5881
rect 8198 5847 8232 5881
rect 8456 5847 8490 5881
rect 8714 5847 8748 5881
rect 8972 5847 9006 5881
rect 9230 5847 9264 5881
rect 9488 5847 9522 5881
rect 9746 5847 9780 5881
rect 10603 5848 10637 5882
rect 10861 5848 10895 5882
rect 11119 5848 11153 5882
rect 11377 5848 11411 5882
rect 11635 5848 11669 5882
rect 11893 5848 11927 5882
rect 12151 5848 12185 5882
rect 12409 5848 12443 5882
rect 5270 5739 5304 5773
rect 5528 5739 5562 5773
rect 5786 5739 5820 5773
rect 6044 5739 6078 5773
rect 6302 5739 6336 5773
rect 6560 5739 6594 5773
rect 6818 5739 6852 5773
rect 7076 5739 7110 5773
rect 7940 5739 7974 5773
rect 8198 5739 8232 5773
rect 8456 5739 8490 5773
rect 8714 5739 8748 5773
rect 8972 5739 9006 5773
rect 9230 5739 9264 5773
rect 9488 5739 9522 5773
rect 9746 5739 9780 5773
rect 10603 5740 10637 5774
rect 10861 5740 10895 5774
rect 11119 5740 11153 5774
rect 11377 5740 11411 5774
rect 11635 5740 11669 5774
rect 11893 5740 11927 5774
rect 12151 5740 12185 5774
rect 12409 5740 12443 5774
rect 5270 5429 5304 5463
rect 5528 5429 5562 5463
rect 5786 5429 5820 5463
rect 6044 5429 6078 5463
rect 6302 5429 6336 5463
rect 6560 5429 6594 5463
rect 6818 5429 6852 5463
rect 7076 5429 7110 5463
rect 7940 5429 7974 5463
rect 8198 5429 8232 5463
rect 8456 5429 8490 5463
rect 8714 5429 8748 5463
rect 8972 5429 9006 5463
rect 9230 5429 9264 5463
rect 9488 5429 9522 5463
rect 9746 5429 9780 5463
rect 10603 5430 10637 5464
rect 10861 5430 10895 5464
rect 11119 5430 11153 5464
rect 11377 5430 11411 5464
rect 11635 5430 11669 5464
rect 11893 5430 11927 5464
rect 12151 5430 12185 5464
rect 12409 5430 12443 5464
rect 5270 5321 5304 5355
rect 5528 5321 5562 5355
rect 5786 5321 5820 5355
rect 6044 5321 6078 5355
rect 6302 5321 6336 5355
rect 6560 5321 6594 5355
rect 6818 5321 6852 5355
rect 7076 5321 7110 5355
rect 7940 5321 7974 5355
rect 8198 5321 8232 5355
rect 8456 5321 8490 5355
rect 8714 5321 8748 5355
rect 8972 5321 9006 5355
rect 9230 5321 9264 5355
rect 9488 5321 9522 5355
rect 9746 5321 9780 5355
rect 10603 5322 10637 5356
rect 10861 5322 10895 5356
rect 11119 5322 11153 5356
rect 11377 5322 11411 5356
rect 11635 5322 11669 5356
rect 11893 5322 11927 5356
rect 12151 5322 12185 5356
rect 12409 5322 12443 5356
rect 5270 5011 5304 5045
rect 5528 5011 5562 5045
rect 5786 5011 5820 5045
rect 6044 5011 6078 5045
rect 6302 5011 6336 5045
rect 6560 5011 6594 5045
rect 6818 5011 6852 5045
rect 7076 5011 7110 5045
rect 7940 5011 7974 5045
rect 8198 5011 8232 5045
rect 8456 5011 8490 5045
rect 8714 5011 8748 5045
rect 8972 5011 9006 5045
rect 9230 5011 9264 5045
rect 9488 5011 9522 5045
rect 9746 5011 9780 5045
rect 10603 5012 10637 5046
rect 10861 5012 10895 5046
rect 11119 5012 11153 5046
rect 11377 5012 11411 5046
rect 11635 5012 11669 5046
rect 11893 5012 11927 5046
rect 12151 5012 12185 5046
rect 12409 5012 12443 5046
rect 5270 4903 5304 4937
rect 5528 4903 5562 4937
rect 5786 4903 5820 4937
rect 6044 4903 6078 4937
rect 6302 4903 6336 4937
rect 6560 4903 6594 4937
rect 6818 4903 6852 4937
rect 7076 4903 7110 4937
rect 7940 4903 7974 4937
rect 8198 4903 8232 4937
rect 8456 4903 8490 4937
rect 8714 4903 8748 4937
rect 8972 4903 9006 4937
rect 9230 4903 9264 4937
rect 9488 4903 9522 4937
rect 9746 4903 9780 4937
rect 10603 4904 10637 4938
rect 10861 4904 10895 4938
rect 11119 4904 11153 4938
rect 11377 4904 11411 4938
rect 11635 4904 11669 4938
rect 11893 4904 11927 4938
rect 12151 4904 12185 4938
rect 12409 4904 12443 4938
rect 5270 4593 5304 4627
rect 5528 4593 5562 4627
rect 5786 4593 5820 4627
rect 6044 4593 6078 4627
rect 6302 4593 6336 4627
rect 6560 4593 6594 4627
rect 6818 4593 6852 4627
rect 7076 4593 7110 4627
rect 7940 4593 7974 4627
rect 8198 4593 8232 4627
rect 8456 4593 8490 4627
rect 8714 4593 8748 4627
rect 8972 4593 9006 4627
rect 9230 4593 9264 4627
rect 9488 4593 9522 4627
rect 9746 4593 9780 4627
rect 10603 4594 10637 4628
rect 10861 4594 10895 4628
rect 11119 4594 11153 4628
rect 11377 4594 11411 4628
rect 11635 4594 11669 4628
rect 11893 4594 11927 4628
rect 12151 4594 12185 4628
rect 12409 4594 12443 4628
rect 5270 4485 5304 4519
rect 5528 4485 5562 4519
rect 5786 4485 5820 4519
rect 6044 4485 6078 4519
rect 6302 4485 6336 4519
rect 6560 4485 6594 4519
rect 6818 4485 6852 4519
rect 7076 4485 7110 4519
rect 7940 4485 7974 4519
rect 8198 4485 8232 4519
rect 8456 4485 8490 4519
rect 8714 4485 8748 4519
rect 8972 4485 9006 4519
rect 9230 4485 9264 4519
rect 9488 4485 9522 4519
rect 9746 4485 9780 4519
rect 10603 4486 10637 4520
rect 10861 4486 10895 4520
rect 11119 4486 11153 4520
rect 11377 4486 11411 4520
rect 11635 4486 11669 4520
rect 11893 4486 11927 4520
rect 12151 4486 12185 4520
rect 12409 4486 12443 4520
rect 5270 4175 5304 4209
rect 5528 4175 5562 4209
rect 5786 4175 5820 4209
rect 6044 4175 6078 4209
rect 6302 4175 6336 4209
rect 6560 4175 6594 4209
rect 6818 4175 6852 4209
rect 7076 4175 7110 4209
rect 7940 4175 7974 4209
rect 8198 4175 8232 4209
rect 8456 4175 8490 4209
rect 8714 4175 8748 4209
rect 8972 4175 9006 4209
rect 9230 4175 9264 4209
rect 9488 4175 9522 4209
rect 9746 4175 9780 4209
rect 10603 4176 10637 4210
rect 10861 4176 10895 4210
rect 11119 4176 11153 4210
rect 11377 4176 11411 4210
rect 11635 4176 11669 4210
rect 11893 4176 11927 4210
rect 12151 4176 12185 4210
rect 12409 4176 12443 4210
rect 5270 4067 5304 4101
rect 5528 4067 5562 4101
rect 5786 4067 5820 4101
rect 6044 4067 6078 4101
rect 6302 4067 6336 4101
rect 6560 4067 6594 4101
rect 6818 4067 6852 4101
rect 7076 4067 7110 4101
rect 7940 4067 7974 4101
rect 8198 4067 8232 4101
rect 8456 4067 8490 4101
rect 8714 4067 8748 4101
rect 8972 4067 9006 4101
rect 9230 4067 9264 4101
rect 9488 4067 9522 4101
rect 9746 4067 9780 4101
rect 10603 4068 10637 4102
rect 10861 4068 10895 4102
rect 11119 4068 11153 4102
rect 11377 4068 11411 4102
rect 11635 4068 11669 4102
rect 11893 4068 11927 4102
rect 12151 4068 12185 4102
rect 12409 4068 12443 4102
rect 5270 3757 5304 3791
rect 5528 3757 5562 3791
rect 5786 3757 5820 3791
rect 6044 3757 6078 3791
rect 6302 3757 6336 3791
rect 6560 3757 6594 3791
rect 6818 3757 6852 3791
rect 7076 3757 7110 3791
rect 7940 3757 7974 3791
rect 8198 3757 8232 3791
rect 8456 3757 8490 3791
rect 8714 3757 8748 3791
rect 8972 3757 9006 3791
rect 9230 3757 9264 3791
rect 9488 3757 9522 3791
rect 9746 3757 9780 3791
rect 10603 3758 10637 3792
rect 10861 3758 10895 3792
rect 11119 3758 11153 3792
rect 11377 3758 11411 3792
rect 11635 3758 11669 3792
rect 11893 3758 11927 3792
rect 12151 3758 12185 3792
rect 12409 3758 12443 3792
rect 5150 3415 5184 3449
rect 5690 3415 5724 3449
rect 6170 3415 6204 3449
rect 6673 3417 6707 3451
rect 7183 3427 7217 3461
rect 7820 3415 7854 3449
rect 8360 3415 8394 3449
rect 8840 3415 8874 3449
rect 9343 3417 9377 3451
rect 9853 3427 9887 3461
rect 10483 3416 10517 3450
rect 5150 3105 5184 3139
rect 5690 3105 5724 3139
rect 6170 3105 6204 3139
rect 6673 3107 6707 3141
rect 11023 3416 11057 3450
rect 11503 3416 11537 3450
rect 12006 3418 12040 3452
rect 12516 3428 12550 3462
rect 7183 3117 7217 3151
rect 7820 3105 7854 3139
rect 8360 3105 8394 3139
rect 8840 3105 8874 3139
rect 9343 3107 9377 3141
rect 9853 3117 9887 3151
rect 10483 3106 10517 3140
rect 11023 3106 11057 3140
rect 11503 3106 11537 3140
rect 12006 3108 12040 3142
rect 12516 3118 12550 3152
rect 5436 1892 5502 1930
rect 6080 1889 6234 1923
rect 6822 1891 6888 1929
rect 7192 1891 7258 1929
rect 7614 1891 7680 1929
rect 8036 1891 8102 1929
rect 8757 1889 8911 1923
rect 9536 1895 9602 1933
rect 9906 1895 9972 1933
rect 10328 1895 10394 1933
rect 10750 1895 10816 1933
rect 11421 1890 11575 1924
rect 12134 1892 12200 1930
rect 6080 1651 6234 1685
rect 8757 1651 8911 1685
rect 11421 1652 11575 1686
rect 5270 858 5304 892
rect 5528 858 5562 892
rect 5786 858 5820 892
rect 6044 858 6078 892
rect 6302 858 6336 892
rect 6560 858 6594 892
rect 6818 858 6852 892
rect 7076 858 7110 892
rect 7940 858 7974 892
rect 8198 858 8232 892
rect 8456 858 8490 892
rect 8714 858 8748 892
rect 8972 858 9006 892
rect 9230 858 9264 892
rect 9488 858 9522 892
rect 9746 858 9780 892
rect 10603 859 10637 893
rect 10861 859 10895 893
rect 11119 859 11153 893
rect 11377 859 11411 893
rect 11635 859 11669 893
rect 11893 859 11927 893
rect 12151 859 12185 893
rect 12409 859 12443 893
rect 5270 548 5304 582
rect 5528 548 5562 582
rect 5786 548 5820 582
rect 6044 548 6078 582
rect 6302 548 6336 582
rect 6560 548 6594 582
rect 6818 548 6852 582
rect 7076 548 7110 582
rect 7940 548 7974 582
rect 8198 548 8232 582
rect 8456 548 8490 582
rect 8714 548 8748 582
rect 8972 548 9006 582
rect 9230 548 9264 582
rect 9488 548 9522 582
rect 9746 548 9780 582
rect 10603 549 10637 583
rect 10861 549 10895 583
rect 11119 549 11153 583
rect 11377 549 11411 583
rect 11635 549 11669 583
rect 11893 549 11927 583
rect 12151 549 12185 583
rect 12409 549 12443 583
rect 5270 440 5304 474
rect 5528 440 5562 474
rect 5786 440 5820 474
rect 6044 440 6078 474
rect 6302 440 6336 474
rect 6560 440 6594 474
rect 6818 440 6852 474
rect 7076 440 7110 474
rect 7940 440 7974 474
rect 8198 440 8232 474
rect 8456 440 8490 474
rect 8714 440 8748 474
rect 8972 440 9006 474
rect 9230 440 9264 474
rect 9488 440 9522 474
rect 9746 440 9780 474
rect 10603 441 10637 475
rect 10861 441 10895 475
rect 11119 441 11153 475
rect 11377 441 11411 475
rect 11635 441 11669 475
rect 11893 441 11927 475
rect 12151 441 12185 475
rect 12409 441 12443 475
rect 5270 130 5304 164
rect 5528 130 5562 164
rect 5786 130 5820 164
rect 6044 130 6078 164
rect 6302 130 6336 164
rect 6560 130 6594 164
rect 6818 130 6852 164
rect 7076 130 7110 164
rect 7940 130 7974 164
rect 8198 130 8232 164
rect 8456 130 8490 164
rect 8714 130 8748 164
rect 8972 130 9006 164
rect 9230 130 9264 164
rect 9488 130 9522 164
rect 9746 130 9780 164
rect 10603 131 10637 165
rect 10861 131 10895 165
rect 11119 131 11153 165
rect 11377 131 11411 165
rect 11635 131 11669 165
rect 11893 131 11927 165
rect 12151 131 12185 165
rect 12409 131 12443 165
rect 5270 22 5304 56
rect 5528 22 5562 56
rect 5786 22 5820 56
rect 6044 22 6078 56
rect 6302 22 6336 56
rect 6560 22 6594 56
rect 6818 22 6852 56
rect 7076 22 7110 56
rect 7940 22 7974 56
rect 8198 22 8232 56
rect 8456 22 8490 56
rect 8714 22 8748 56
rect 8972 22 9006 56
rect 9230 22 9264 56
rect 9488 22 9522 56
rect 9746 22 9780 56
rect 10603 23 10637 57
rect 10861 23 10895 57
rect 11119 23 11153 57
rect 11377 23 11411 57
rect 11635 23 11669 57
rect 11893 23 11927 57
rect 12151 23 12185 57
rect 12409 23 12443 57
rect 5270 -288 5304 -254
rect 5528 -288 5562 -254
rect 5786 -288 5820 -254
rect 6044 -288 6078 -254
rect 6302 -288 6336 -254
rect 6560 -288 6594 -254
rect 6818 -288 6852 -254
rect 7076 -288 7110 -254
rect 7940 -288 7974 -254
rect 8198 -288 8232 -254
rect 8456 -288 8490 -254
rect 8714 -288 8748 -254
rect 8972 -288 9006 -254
rect 9230 -288 9264 -254
rect 9488 -288 9522 -254
rect 9746 -288 9780 -254
rect 10603 -287 10637 -253
rect 10861 -287 10895 -253
rect 11119 -287 11153 -253
rect 11377 -287 11411 -253
rect 11635 -287 11669 -253
rect 11893 -287 11927 -253
rect 12151 -287 12185 -253
rect 12409 -287 12443 -253
rect 5270 -396 5304 -362
rect 5528 -396 5562 -362
rect 5786 -396 5820 -362
rect 6044 -396 6078 -362
rect 6302 -396 6336 -362
rect 6560 -396 6594 -362
rect 6818 -396 6852 -362
rect 7076 -396 7110 -362
rect 7940 -396 7974 -362
rect 8198 -396 8232 -362
rect 8456 -396 8490 -362
rect 8714 -396 8748 -362
rect 8972 -396 9006 -362
rect 9230 -396 9264 -362
rect 9488 -396 9522 -362
rect 9746 -396 9780 -362
rect 10603 -395 10637 -361
rect 10861 -395 10895 -361
rect 11119 -395 11153 -361
rect 11377 -395 11411 -361
rect 11635 -395 11669 -361
rect 11893 -395 11927 -361
rect 12151 -395 12185 -361
rect 12409 -395 12443 -361
rect 5270 -706 5304 -672
rect 5528 -706 5562 -672
rect 5786 -706 5820 -672
rect 6044 -706 6078 -672
rect 6302 -706 6336 -672
rect 6560 -706 6594 -672
rect 6818 -706 6852 -672
rect 7076 -706 7110 -672
rect 7940 -706 7974 -672
rect 8198 -706 8232 -672
rect 8456 -706 8490 -672
rect 8714 -706 8748 -672
rect 8972 -706 9006 -672
rect 9230 -706 9264 -672
rect 9488 -706 9522 -672
rect 9746 -706 9780 -672
rect 10603 -705 10637 -671
rect 10861 -705 10895 -671
rect 11119 -705 11153 -671
rect 11377 -705 11411 -671
rect 11635 -705 11669 -671
rect 11893 -705 11927 -671
rect 12151 -705 12185 -671
rect 12409 -705 12443 -671
rect 5270 -814 5304 -780
rect 5528 -814 5562 -780
rect 5786 -814 5820 -780
rect 6044 -814 6078 -780
rect 6302 -814 6336 -780
rect 6560 -814 6594 -780
rect 6818 -814 6852 -780
rect 7076 -814 7110 -780
rect 7940 -814 7974 -780
rect 8198 -814 8232 -780
rect 8456 -814 8490 -780
rect 8714 -814 8748 -780
rect 8972 -814 9006 -780
rect 9230 -814 9264 -780
rect 9488 -814 9522 -780
rect 9746 -814 9780 -780
rect 10603 -813 10637 -779
rect 10861 -813 10895 -779
rect 11119 -813 11153 -779
rect 11377 -813 11411 -779
rect 11635 -813 11669 -779
rect 11893 -813 11927 -779
rect 12151 -813 12185 -779
rect 12409 -813 12443 -779
rect 5270 -1124 5304 -1090
rect 5528 -1124 5562 -1090
rect 5786 -1124 5820 -1090
rect 6044 -1124 6078 -1090
rect 6302 -1124 6336 -1090
rect 6560 -1124 6594 -1090
rect 6818 -1124 6852 -1090
rect 7076 -1124 7110 -1090
rect 7940 -1124 7974 -1090
rect 8198 -1124 8232 -1090
rect 8456 -1124 8490 -1090
rect 8714 -1124 8748 -1090
rect 8972 -1124 9006 -1090
rect 9230 -1124 9264 -1090
rect 9488 -1124 9522 -1090
rect 9746 -1124 9780 -1090
rect 10603 -1123 10637 -1089
rect 10861 -1123 10895 -1089
rect 11119 -1123 11153 -1089
rect 11377 -1123 11411 -1089
rect 11635 -1123 11669 -1089
rect 11893 -1123 11927 -1089
rect 12151 -1123 12185 -1089
rect 12409 -1123 12443 -1089
rect 5270 -1232 5304 -1198
rect 5528 -1232 5562 -1198
rect 5786 -1232 5820 -1198
rect 6044 -1232 6078 -1198
rect 6302 -1232 6336 -1198
rect 6560 -1232 6594 -1198
rect 6818 -1232 6852 -1198
rect 7076 -1232 7110 -1198
rect 7940 -1232 7974 -1198
rect 8198 -1232 8232 -1198
rect 8456 -1232 8490 -1198
rect 8714 -1232 8748 -1198
rect 8972 -1232 9006 -1198
rect 9230 -1232 9264 -1198
rect 9488 -1232 9522 -1198
rect 9746 -1232 9780 -1198
rect 10603 -1231 10637 -1197
rect 10861 -1231 10895 -1197
rect 11119 -1231 11153 -1197
rect 11377 -1231 11411 -1197
rect 11635 -1231 11669 -1197
rect 11893 -1231 11927 -1197
rect 12151 -1231 12185 -1197
rect 12409 -1231 12443 -1197
rect 5270 -1542 5304 -1508
rect 5528 -1542 5562 -1508
rect 5786 -1542 5820 -1508
rect 6044 -1542 6078 -1508
rect 6302 -1542 6336 -1508
rect 6560 -1542 6594 -1508
rect 6818 -1542 6852 -1508
rect 7076 -1542 7110 -1508
rect 7940 -1542 7974 -1508
rect 8198 -1542 8232 -1508
rect 8456 -1542 8490 -1508
rect 8714 -1542 8748 -1508
rect 8972 -1542 9006 -1508
rect 9230 -1542 9264 -1508
rect 9488 -1542 9522 -1508
rect 9746 -1542 9780 -1508
rect 10603 -1541 10637 -1507
rect 10861 -1541 10895 -1507
rect 11119 -1541 11153 -1507
rect 11377 -1541 11411 -1507
rect 11635 -1541 11669 -1507
rect 11893 -1541 11927 -1507
rect 12151 -1541 12185 -1507
rect 12409 -1541 12443 -1507
rect 5270 -1650 5304 -1616
rect 5528 -1650 5562 -1616
rect 5786 -1650 5820 -1616
rect 6044 -1650 6078 -1616
rect 6302 -1650 6336 -1616
rect 6560 -1650 6594 -1616
rect 6818 -1650 6852 -1616
rect 7076 -1650 7110 -1616
rect 7940 -1650 7974 -1616
rect 8198 -1650 8232 -1616
rect 8456 -1650 8490 -1616
rect 8714 -1650 8748 -1616
rect 8972 -1650 9006 -1616
rect 9230 -1650 9264 -1616
rect 9488 -1650 9522 -1616
rect 9746 -1650 9780 -1616
rect 10603 -1649 10637 -1615
rect 10861 -1649 10895 -1615
rect 11119 -1649 11153 -1615
rect 11377 -1649 11411 -1615
rect 11635 -1649 11669 -1615
rect 11893 -1649 11927 -1615
rect 12151 -1649 12185 -1615
rect 12409 -1649 12443 -1615
rect 5270 -1960 5304 -1926
rect 5528 -1960 5562 -1926
rect 5786 -1960 5820 -1926
rect 6044 -1960 6078 -1926
rect 6302 -1960 6336 -1926
rect 6560 -1960 6594 -1926
rect 6818 -1960 6852 -1926
rect 7076 -1960 7110 -1926
rect 7940 -1960 7974 -1926
rect 8198 -1960 8232 -1926
rect 8456 -1960 8490 -1926
rect 8714 -1960 8748 -1926
rect 8972 -1960 9006 -1926
rect 9230 -1960 9264 -1926
rect 9488 -1960 9522 -1926
rect 9746 -1960 9780 -1926
rect 10603 -1959 10637 -1925
rect 10861 -1959 10895 -1925
rect 11119 -1959 11153 -1925
rect 11377 -1959 11411 -1925
rect 11635 -1959 11669 -1925
rect 11893 -1959 11927 -1925
rect 12151 -1959 12185 -1925
rect 12409 -1959 12443 -1925
rect 5150 -2302 5184 -2268
rect 5690 -2302 5724 -2268
rect 6170 -2302 6204 -2268
rect 6673 -2300 6707 -2266
rect 7183 -2290 7217 -2256
rect 7820 -2302 7854 -2268
rect 8360 -2302 8394 -2268
rect 8840 -2302 8874 -2268
rect 9343 -2300 9377 -2266
rect 9853 -2290 9887 -2256
rect 10483 -2301 10517 -2267
rect 5150 -2612 5184 -2578
rect 5690 -2612 5724 -2578
rect 6170 -2612 6204 -2578
rect 6673 -2610 6707 -2576
rect 11023 -2301 11057 -2267
rect 11503 -2301 11537 -2267
rect 12006 -2299 12040 -2265
rect 12516 -2289 12550 -2255
rect 7183 -2600 7217 -2566
rect 7820 -2612 7854 -2578
rect 8360 -2612 8394 -2578
rect 8840 -2612 8874 -2578
rect 9343 -2610 9377 -2576
rect 9853 -2600 9887 -2566
rect 10483 -2611 10517 -2577
rect 11023 -2611 11057 -2577
rect 11503 -2611 11537 -2577
rect 12006 -2609 12040 -2575
rect 12516 -2599 12550 -2565
rect 12726 -3402 12760 -3368
rect 5481 -4032 5547 -3994
rect 6088 -4036 6242 -4002
rect 6822 -4034 6888 -3996
rect 7192 -4034 7258 -3996
rect 7614 -4034 7680 -3996
rect 8036 -4034 8102 -3996
rect 8758 -4036 8912 -4002
rect 9523 -4034 9589 -3996
rect 9893 -4034 9959 -3996
rect 10315 -4034 10381 -3996
rect 10737 -4034 10803 -3996
rect 11421 -4035 11575 -4001
rect 6088 -4274 6242 -4240
rect 8758 -4274 8912 -4240
rect 11421 -4273 11575 -4239
rect 13116 -3404 13150 -3370
rect 12726 -3866 12760 -3832
rect 13116 -3868 13150 -3834
rect 12730 -4198 12764 -4164
rect 13120 -4198 13154 -4164
rect 12730 -4392 12764 -4358
rect 13120 -4392 13154 -4358
rect 5270 -5046 5304 -5012
rect 5528 -5046 5562 -5012
rect 5786 -5046 5820 -5012
rect 6044 -5046 6078 -5012
rect 6302 -5046 6336 -5012
rect 6560 -5046 6594 -5012
rect 6818 -5046 6852 -5012
rect 7076 -5046 7110 -5012
rect 7940 -5046 7974 -5012
rect 8198 -5046 8232 -5012
rect 8456 -5046 8490 -5012
rect 8714 -5046 8748 -5012
rect 8972 -5046 9006 -5012
rect 9230 -5046 9264 -5012
rect 9488 -5046 9522 -5012
rect 9746 -5046 9780 -5012
rect 10603 -5045 10637 -5011
rect 10861 -5045 10895 -5011
rect 11119 -5045 11153 -5011
rect 11377 -5045 11411 -5011
rect 11635 -5045 11669 -5011
rect 11893 -5045 11927 -5011
rect 12151 -5045 12185 -5011
rect 12409 -5045 12443 -5011
rect 5270 -5356 5304 -5322
rect 5528 -5356 5562 -5322
rect 5786 -5356 5820 -5322
rect 6044 -5356 6078 -5322
rect 6302 -5356 6336 -5322
rect 6560 -5356 6594 -5322
rect 6818 -5356 6852 -5322
rect 7076 -5356 7110 -5322
rect 7940 -5356 7974 -5322
rect 8198 -5356 8232 -5322
rect 8456 -5356 8490 -5322
rect 8714 -5356 8748 -5322
rect 8972 -5356 9006 -5322
rect 9230 -5356 9264 -5322
rect 9488 -5356 9522 -5322
rect 9746 -5356 9780 -5322
rect 10603 -5355 10637 -5321
rect 10861 -5355 10895 -5321
rect 11119 -5355 11153 -5321
rect 11377 -5355 11411 -5321
rect 11635 -5355 11669 -5321
rect 11893 -5355 11927 -5321
rect 12151 -5355 12185 -5321
rect 12409 -5355 12443 -5321
rect 5270 -5464 5304 -5430
rect 5528 -5464 5562 -5430
rect 5786 -5464 5820 -5430
rect 6044 -5464 6078 -5430
rect 6302 -5464 6336 -5430
rect 6560 -5464 6594 -5430
rect 6818 -5464 6852 -5430
rect 7076 -5464 7110 -5430
rect 7940 -5464 7974 -5430
rect 8198 -5464 8232 -5430
rect 8456 -5464 8490 -5430
rect 8714 -5464 8748 -5430
rect 8972 -5464 9006 -5430
rect 9230 -5464 9264 -5430
rect 9488 -5464 9522 -5430
rect 9746 -5464 9780 -5430
rect 10603 -5463 10637 -5429
rect 10861 -5463 10895 -5429
rect 11119 -5463 11153 -5429
rect 11377 -5463 11411 -5429
rect 11635 -5463 11669 -5429
rect 11893 -5463 11927 -5429
rect 12151 -5463 12185 -5429
rect 12409 -5463 12443 -5429
rect 5270 -5774 5304 -5740
rect 5528 -5774 5562 -5740
rect 5786 -5774 5820 -5740
rect 6044 -5774 6078 -5740
rect 6302 -5774 6336 -5740
rect 6560 -5774 6594 -5740
rect 6818 -5774 6852 -5740
rect 7076 -5774 7110 -5740
rect 7940 -5774 7974 -5740
rect 8198 -5774 8232 -5740
rect 8456 -5774 8490 -5740
rect 8714 -5774 8748 -5740
rect 8972 -5774 9006 -5740
rect 9230 -5774 9264 -5740
rect 9488 -5774 9522 -5740
rect 9746 -5774 9780 -5740
rect 10603 -5773 10637 -5739
rect 10861 -5773 10895 -5739
rect 11119 -5773 11153 -5739
rect 11377 -5773 11411 -5739
rect 11635 -5773 11669 -5739
rect 11893 -5773 11927 -5739
rect 12151 -5773 12185 -5739
rect 12409 -5773 12443 -5739
rect 5270 -5882 5304 -5848
rect 5528 -5882 5562 -5848
rect 5786 -5882 5820 -5848
rect 6044 -5882 6078 -5848
rect 6302 -5882 6336 -5848
rect 6560 -5882 6594 -5848
rect 6818 -5882 6852 -5848
rect 7076 -5882 7110 -5848
rect 7940 -5882 7974 -5848
rect 8198 -5882 8232 -5848
rect 8456 -5882 8490 -5848
rect 8714 -5882 8748 -5848
rect 8972 -5882 9006 -5848
rect 9230 -5882 9264 -5848
rect 9488 -5882 9522 -5848
rect 9746 -5882 9780 -5848
rect 10603 -5881 10637 -5847
rect 10861 -5881 10895 -5847
rect 11119 -5881 11153 -5847
rect 11377 -5881 11411 -5847
rect 11635 -5881 11669 -5847
rect 11893 -5881 11927 -5847
rect 12151 -5881 12185 -5847
rect 12409 -5881 12443 -5847
rect 5270 -6192 5304 -6158
rect 5528 -6192 5562 -6158
rect 5786 -6192 5820 -6158
rect 6044 -6192 6078 -6158
rect 6302 -6192 6336 -6158
rect 6560 -6192 6594 -6158
rect 6818 -6192 6852 -6158
rect 7076 -6192 7110 -6158
rect 7940 -6192 7974 -6158
rect 8198 -6192 8232 -6158
rect 8456 -6192 8490 -6158
rect 8714 -6192 8748 -6158
rect 8972 -6192 9006 -6158
rect 9230 -6192 9264 -6158
rect 9488 -6192 9522 -6158
rect 9746 -6192 9780 -6158
rect 10603 -6191 10637 -6157
rect 10861 -6191 10895 -6157
rect 11119 -6191 11153 -6157
rect 11377 -6191 11411 -6157
rect 11635 -6191 11669 -6157
rect 11893 -6191 11927 -6157
rect 12151 -6191 12185 -6157
rect 12409 -6191 12443 -6157
rect 5270 -6300 5304 -6266
rect 5528 -6300 5562 -6266
rect 5786 -6300 5820 -6266
rect 6044 -6300 6078 -6266
rect 6302 -6300 6336 -6266
rect 6560 -6300 6594 -6266
rect 6818 -6300 6852 -6266
rect 7076 -6300 7110 -6266
rect 7940 -6300 7974 -6266
rect 8198 -6300 8232 -6266
rect 8456 -6300 8490 -6266
rect 8714 -6300 8748 -6266
rect 8972 -6300 9006 -6266
rect 9230 -6300 9264 -6266
rect 9488 -6300 9522 -6266
rect 9746 -6300 9780 -6266
rect 10603 -6299 10637 -6265
rect 10861 -6299 10895 -6265
rect 11119 -6299 11153 -6265
rect 11377 -6299 11411 -6265
rect 11635 -6299 11669 -6265
rect 11893 -6299 11927 -6265
rect 12151 -6299 12185 -6265
rect 12409 -6299 12443 -6265
rect 5270 -6610 5304 -6576
rect 5528 -6610 5562 -6576
rect 5786 -6610 5820 -6576
rect 6044 -6610 6078 -6576
rect 6302 -6610 6336 -6576
rect 6560 -6610 6594 -6576
rect 6818 -6610 6852 -6576
rect 7076 -6610 7110 -6576
rect 7940 -6610 7974 -6576
rect 8198 -6610 8232 -6576
rect 8456 -6610 8490 -6576
rect 8714 -6610 8748 -6576
rect 8972 -6610 9006 -6576
rect 9230 -6610 9264 -6576
rect 9488 -6610 9522 -6576
rect 9746 -6610 9780 -6576
rect 10603 -6609 10637 -6575
rect 10861 -6609 10895 -6575
rect 11119 -6609 11153 -6575
rect 11377 -6609 11411 -6575
rect 11635 -6609 11669 -6575
rect 11893 -6609 11927 -6575
rect 12151 -6609 12185 -6575
rect 12409 -6609 12443 -6575
rect 5270 -6718 5304 -6684
rect 5528 -6718 5562 -6684
rect 5786 -6718 5820 -6684
rect 6044 -6718 6078 -6684
rect 6302 -6718 6336 -6684
rect 6560 -6718 6594 -6684
rect 6818 -6718 6852 -6684
rect 7076 -6718 7110 -6684
rect 7940 -6718 7974 -6684
rect 8198 -6718 8232 -6684
rect 8456 -6718 8490 -6684
rect 8714 -6718 8748 -6684
rect 8972 -6718 9006 -6684
rect 9230 -6718 9264 -6684
rect 9488 -6718 9522 -6684
rect 9746 -6718 9780 -6684
rect 10603 -6717 10637 -6683
rect 10861 -6717 10895 -6683
rect 11119 -6717 11153 -6683
rect 11377 -6717 11411 -6683
rect 11635 -6717 11669 -6683
rect 11893 -6717 11927 -6683
rect 12151 -6717 12185 -6683
rect 12409 -6717 12443 -6683
rect 5270 -7028 5304 -6994
rect 5528 -7028 5562 -6994
rect 5786 -7028 5820 -6994
rect 6044 -7028 6078 -6994
rect 6302 -7028 6336 -6994
rect 6560 -7028 6594 -6994
rect 6818 -7028 6852 -6994
rect 7076 -7028 7110 -6994
rect 7940 -7028 7974 -6994
rect 8198 -7028 8232 -6994
rect 8456 -7028 8490 -6994
rect 8714 -7028 8748 -6994
rect 8972 -7028 9006 -6994
rect 9230 -7028 9264 -6994
rect 9488 -7028 9522 -6994
rect 9746 -7028 9780 -6994
rect 10603 -7027 10637 -6993
rect 10861 -7027 10895 -6993
rect 11119 -7027 11153 -6993
rect 11377 -7027 11411 -6993
rect 11635 -7027 11669 -6993
rect 11893 -7027 11927 -6993
rect 12151 -7027 12185 -6993
rect 12409 -7027 12443 -6993
rect 5270 -7136 5304 -7102
rect 5528 -7136 5562 -7102
rect 5786 -7136 5820 -7102
rect 6044 -7136 6078 -7102
rect 6302 -7136 6336 -7102
rect 6560 -7136 6594 -7102
rect 6818 -7136 6852 -7102
rect 7076 -7136 7110 -7102
rect 7940 -7136 7974 -7102
rect 8198 -7136 8232 -7102
rect 8456 -7136 8490 -7102
rect 8714 -7136 8748 -7102
rect 8972 -7136 9006 -7102
rect 9230 -7136 9264 -7102
rect 9488 -7136 9522 -7102
rect 9746 -7136 9780 -7102
rect 10603 -7135 10637 -7101
rect 10861 -7135 10895 -7101
rect 11119 -7135 11153 -7101
rect 11377 -7135 11411 -7101
rect 11635 -7135 11669 -7101
rect 11893 -7135 11927 -7101
rect 12151 -7135 12185 -7101
rect 12409 -7135 12443 -7101
rect 5270 -7446 5304 -7412
rect 5528 -7446 5562 -7412
rect 5786 -7446 5820 -7412
rect 6044 -7446 6078 -7412
rect 6302 -7446 6336 -7412
rect 6560 -7446 6594 -7412
rect 6818 -7446 6852 -7412
rect 7076 -7446 7110 -7412
rect 7940 -7446 7974 -7412
rect 8198 -7446 8232 -7412
rect 8456 -7446 8490 -7412
rect 8714 -7446 8748 -7412
rect 8972 -7446 9006 -7412
rect 9230 -7446 9264 -7412
rect 9488 -7446 9522 -7412
rect 9746 -7446 9780 -7412
rect 10603 -7445 10637 -7411
rect 10861 -7445 10895 -7411
rect 11119 -7445 11153 -7411
rect 11377 -7445 11411 -7411
rect 11635 -7445 11669 -7411
rect 11893 -7445 11927 -7411
rect 12151 -7445 12185 -7411
rect 12409 -7445 12443 -7411
rect 5270 -7554 5304 -7520
rect 5528 -7554 5562 -7520
rect 5786 -7554 5820 -7520
rect 6044 -7554 6078 -7520
rect 6302 -7554 6336 -7520
rect 6560 -7554 6594 -7520
rect 6818 -7554 6852 -7520
rect 7076 -7554 7110 -7520
rect 7940 -7554 7974 -7520
rect 8198 -7554 8232 -7520
rect 8456 -7554 8490 -7520
rect 8714 -7554 8748 -7520
rect 8972 -7554 9006 -7520
rect 9230 -7554 9264 -7520
rect 9488 -7554 9522 -7520
rect 9746 -7554 9780 -7520
rect 10603 -7553 10637 -7519
rect 10861 -7553 10895 -7519
rect 11119 -7553 11153 -7519
rect 11377 -7553 11411 -7519
rect 11635 -7553 11669 -7519
rect 11893 -7553 11927 -7519
rect 12151 -7553 12185 -7519
rect 12409 -7553 12443 -7519
rect 5270 -7864 5304 -7830
rect 5528 -7864 5562 -7830
rect 5786 -7864 5820 -7830
rect 6044 -7864 6078 -7830
rect 6302 -7864 6336 -7830
rect 6560 -7864 6594 -7830
rect 6818 -7864 6852 -7830
rect 7076 -7864 7110 -7830
rect 7940 -7864 7974 -7830
rect 8198 -7864 8232 -7830
rect 8456 -7864 8490 -7830
rect 8714 -7864 8748 -7830
rect 8972 -7864 9006 -7830
rect 9230 -7864 9264 -7830
rect 9488 -7864 9522 -7830
rect 9746 -7864 9780 -7830
rect 10603 -7863 10637 -7829
rect 10861 -7863 10895 -7829
rect 11119 -7863 11153 -7829
rect 11377 -7863 11411 -7829
rect 11635 -7863 11669 -7829
rect 11893 -7863 11927 -7829
rect 12151 -7863 12185 -7829
rect 12409 -7863 12443 -7829
rect 5150 -8206 5184 -8172
rect 5690 -8206 5724 -8172
rect 6170 -8206 6204 -8172
rect 6673 -8204 6707 -8170
rect 7183 -8194 7217 -8160
rect 7820 -8206 7854 -8172
rect 8360 -8206 8394 -8172
rect 8840 -8206 8874 -8172
rect 9343 -8204 9377 -8170
rect 9853 -8194 9887 -8160
rect 10483 -8205 10517 -8171
rect 5150 -8516 5184 -8482
rect 5690 -8516 5724 -8482
rect 6170 -8516 6204 -8482
rect 6673 -8514 6707 -8480
rect 11023 -8205 11057 -8171
rect 11503 -8205 11537 -8171
rect 12006 -8203 12040 -8169
rect 12516 -8193 12550 -8159
rect 7183 -8504 7217 -8470
rect 7820 -8516 7854 -8482
rect 8360 -8516 8394 -8482
rect 8840 -8516 8874 -8482
rect 9343 -8514 9377 -8480
rect 9853 -8504 9887 -8470
rect 10483 -8515 10517 -8481
rect 11023 -8515 11057 -8481
rect 11503 -8515 11537 -8481
rect 12006 -8513 12040 -8479
rect 12516 -8503 12550 -8469
rect 14080 8589 15448 8623
rect 15941 8589 17306 8623
rect 14080 7079 15448 7113
rect 15941 7079 17306 7113
rect 14080 5569 15448 5603
rect 15941 5569 17306 5603
rect 14080 4059 15448 4093
rect 15941 4059 17306 4093
rect 14080 2549 15448 2583
rect 15941 2549 17306 2583
rect 14080 1039 15448 1073
rect 15941 1039 17306 1073
rect 14080 -471 15448 -437
rect 15941 -471 17306 -437
rect 14080 -1981 15448 -1947
rect 15941 -1981 17306 -1947
rect 14080 -3491 15448 -3457
rect 15941 -3491 17306 -3457
rect 14080 -5001 15448 -4967
rect 15941 -5001 17306 -4967
rect 14080 -6511 15448 -6477
rect 15941 -6511 17306 -6477
rect 14080 -8021 15448 -7987
rect 15941 -8021 17306 -7987
rect 14080 -9531 15448 -9497
rect 15941 -9531 17306 -9497
<< locali >>
rect 500 8930 17271 9162
rect 500 8902 17272 8930
rect 503 8660 3651 8902
rect 503 8622 1824 8660
rect 2046 8658 2096 8660
rect 443 8588 459 8622
rect 397 8538 431 8554
rect 397 7146 431 7162
rect 503 7112 1824 8588
rect 2318 8622 3651 8660
rect 3685 8588 3701 8622
rect 2038 8538 2108 8560
rect 2038 8518 2055 8538
rect 443 7078 459 7112
rect 397 7028 431 7044
rect 397 5636 431 5652
rect 503 5602 1824 7078
rect 443 5568 459 5602
rect 397 5518 431 5534
rect 397 4126 431 4142
rect 503 4092 1824 5568
rect 443 4058 459 4092
rect 397 4008 431 4024
rect 397 2616 431 2632
rect 503 2582 1824 4058
rect 443 2548 459 2582
rect 397 2498 431 2514
rect 397 1106 431 1122
rect 503 1072 1824 2548
rect 443 1038 459 1072
rect 397 988 431 1004
rect 397 -404 431 -388
rect 503 -438 1824 1038
rect 443 -472 459 -438
rect 397 -522 431 -506
rect 397 -1914 431 -1898
rect 503 -1948 1824 -472
rect 443 -1982 459 -1948
rect 397 -2032 431 -2016
rect 397 -3424 431 -3408
rect 503 -3458 1824 -1982
rect 443 -3492 459 -3458
rect 397 -3542 431 -3526
rect 397 -4934 431 -4918
rect 503 -4968 1824 -3492
rect 443 -5002 459 -4968
rect 397 -5052 431 -5036
rect 397 -6444 431 -6428
rect 503 -6478 1824 -5002
rect 443 -6512 459 -6478
rect 397 -6562 431 -6546
rect 397 -7954 431 -7938
rect 503 -7988 1824 -6512
rect 443 -8022 459 -7988
rect 397 -8072 431 -8056
rect 397 -9464 431 -9448
rect 503 -9498 1824 -8022
rect 443 -9532 459 -9498
rect 503 -9548 1824 -9532
rect 2046 7162 2055 8518
rect 2089 8518 2108 8538
rect 2089 7162 2096 8518
rect 2046 7028 2096 7162
rect 2046 5652 2055 7028
rect 2089 5652 2096 7028
rect 2046 5518 2096 5652
rect 2046 4142 2055 5518
rect 2089 4142 2096 5518
rect 2046 4008 2096 4142
rect 2046 2632 2055 4008
rect 2089 2632 2096 4008
rect 2046 2498 2096 2632
rect 2046 1122 2055 2498
rect 2089 1122 2096 2498
rect 2046 988 2096 1122
rect 2046 -388 2055 988
rect 2089 -388 2096 988
rect 2046 -522 2096 -388
rect 2046 -1898 2055 -522
rect 2089 -1898 2096 -522
rect 2046 -2032 2096 -1898
rect 2046 -3408 2055 -2032
rect 2089 -3408 2096 -2032
rect 2046 -3542 2096 -3408
rect 2046 -4918 2055 -3542
rect 2089 -4918 2096 -3542
rect 2046 -5052 2096 -4918
rect 2046 -6428 2055 -5052
rect 2089 -6428 2096 -5052
rect 2046 -6562 2096 -6428
rect 2046 -7938 2055 -6562
rect 2089 -7938 2096 -6562
rect 2046 -8072 2096 -7938
rect 2046 -9448 2055 -8072
rect 2089 -9448 2096 -8072
rect 2046 -9548 2096 -9448
rect 2318 8502 3651 8588
rect 3713 8538 3747 8554
rect 2318 7112 3647 8502
rect 3713 7146 3747 7162
rect 3685 7078 3701 7112
rect 2318 5602 3647 7078
rect 3713 7028 3747 7044
rect 3713 5636 3747 5652
rect 3685 5568 3701 5602
rect 2318 4092 3647 5568
rect 3713 5518 3747 5534
rect 3713 4126 3747 4142
rect 3685 4058 3701 4092
rect 2318 2582 3647 4058
rect 3713 4008 3747 4024
rect 3713 2616 3747 2632
rect 3685 2548 3701 2582
rect 2318 1072 3647 2548
rect 3713 2498 3747 2514
rect 3713 1106 3747 1122
rect 3685 1038 3701 1072
rect 2318 -438 3647 1038
rect 3713 988 3747 1004
rect 3713 -404 3747 -388
rect 3685 -472 3701 -438
rect 2318 -1948 3647 -472
rect 3713 -522 3747 -506
rect 3713 -1914 3747 -1898
rect 3685 -1982 3701 -1948
rect 2318 -3458 3647 -1982
rect 3713 -2032 3747 -2016
rect 3713 -3424 3747 -3408
rect 3685 -3492 3701 -3458
rect 2318 -4968 3647 -3492
rect 3713 -3542 3747 -3526
rect 3713 -4934 3747 -4918
rect 3685 -5002 3701 -4968
rect 2318 -6478 3647 -5002
rect 3713 -5052 3747 -5036
rect 3713 -6444 3747 -6428
rect 3685 -6512 3701 -6478
rect 2318 -7988 3647 -6512
rect 3713 -6562 3747 -6546
rect 3713 -7954 3747 -7938
rect 3685 -8022 3701 -7988
rect 2318 -9498 3647 -8022
rect 3713 -8072 3747 -8056
rect 3713 -9464 3747 -9448
rect 3685 -9532 3701 -9498
rect 2318 -9548 3647 -9532
rect 4498 8052 4820 8902
rect 6056 8794 10038 8803
rect 6056 8699 6194 8794
rect 6822 8790 10038 8794
rect 6822 8699 8974 8790
rect 6056 8695 8974 8699
rect 9602 8695 10038 8790
rect 6056 8633 10038 8695
rect 10750 8671 11844 8672
rect 6060 8632 8223 8633
rect 8944 8632 10038 8633
rect 6060 8631 7129 8632
rect 5400 8614 5453 8615
rect 5400 8579 5730 8614
rect 5400 8545 5544 8579
rect 5578 8545 5730 8579
rect 5400 8500 5730 8545
rect 6060 8508 6113 8631
rect 6188 8545 6204 8579
rect 6238 8545 6254 8579
rect 6658 8570 6674 8579
rect 6529 8545 6674 8570
rect 6708 8570 6724 8579
rect 7123 8578 8490 8595
rect 6708 8545 6859 8570
rect 6060 8500 6114 8508
rect 5401 8490 5730 8500
rect 5401 8454 5416 8490
rect 5450 8486 5730 8490
rect 5450 8454 5673 8486
rect 5401 8450 5673 8454
rect 5707 8450 5730 8486
rect 5401 8416 5730 8450
rect 5401 8380 5415 8416
rect 5449 8380 5673 8416
rect 5707 8380 5730 8416
rect 5401 8343 5730 8380
rect 5401 8307 5415 8343
rect 5449 8307 5672 8343
rect 5706 8307 5730 8343
rect 5401 8251 5730 8307
rect 6061 8490 6114 8500
rect 6061 8454 6076 8490
rect 6110 8454 6114 8490
rect 6061 8416 6114 8454
rect 6061 8380 6075 8416
rect 6109 8380 6114 8416
rect 6061 8343 6114 8380
rect 6061 8307 6075 8343
rect 6109 8307 6114 8343
rect 6061 8274 6114 8307
rect 6328 8486 6388 8502
rect 6328 8450 6333 8486
rect 6367 8450 6388 8486
rect 6328 8416 6388 8450
rect 6328 8380 6333 8416
rect 6367 8380 6388 8416
rect 6328 8343 6388 8380
rect 6328 8307 6332 8343
rect 6366 8307 6388 8343
rect 6328 8296 6388 8307
rect 6529 8490 6859 8545
rect 6529 8454 6546 8490
rect 6580 8486 6859 8490
rect 6580 8454 6803 8486
rect 6529 8450 6803 8454
rect 6837 8450 6859 8486
rect 6529 8416 6859 8450
rect 6529 8380 6545 8416
rect 6579 8380 6803 8416
rect 6837 8380 6859 8416
rect 6529 8343 6859 8380
rect 6529 8307 6545 8343
rect 6579 8307 6802 8343
rect 6836 8307 6859 8343
rect 6529 8296 6859 8307
rect 7123 8544 7277 8578
rect 7311 8544 7535 8578
rect 7569 8544 7793 8578
rect 7827 8544 8051 8578
rect 8085 8544 8309 8578
rect 8343 8544 8490 8578
rect 7123 8486 8490 8544
rect 7123 8450 7148 8486
rect 7182 8450 7406 8486
rect 7440 8450 7664 8486
rect 7698 8450 7922 8486
rect 7956 8450 8180 8486
rect 8214 8450 8438 8486
rect 8472 8450 8490 8486
rect 7123 8415 8490 8450
rect 7123 8379 7148 8415
rect 7182 8379 7406 8415
rect 7440 8379 7664 8415
rect 7698 8379 7922 8415
rect 7956 8379 8180 8415
rect 8214 8379 8438 8415
rect 8472 8379 8490 8415
rect 7123 8344 8490 8379
rect 7123 8308 7148 8344
rect 7182 8308 7406 8344
rect 7440 8308 7664 8344
rect 7698 8308 7922 8344
rect 7956 8308 8180 8344
rect 8214 8308 8438 8344
rect 8472 8308 8490 8344
rect 5401 8217 5544 8251
rect 5578 8217 5730 8251
rect 6188 8217 6204 8251
rect 6238 8217 6254 8251
rect 5401 8171 5730 8217
rect 6328 8052 6390 8296
rect 6529 8251 6860 8296
rect 6529 8217 6674 8251
rect 6708 8217 6860 8251
rect 6529 8172 6860 8217
rect 7123 8250 8490 8308
rect 8944 8486 9004 8632
rect 9076 8544 9092 8578
rect 9126 8544 9142 8578
rect 9334 8544 9350 8578
rect 9384 8544 9400 8578
rect 8944 8450 8963 8486
rect 8997 8450 9004 8486
rect 8944 8415 9004 8450
rect 8944 8379 8963 8415
rect 8997 8379 9004 8415
rect 8944 8344 9004 8379
rect 8944 8308 8963 8344
rect 8997 8308 9004 8344
rect 8944 8273 9004 8308
rect 9212 8486 9263 8516
rect 9212 8450 9221 8486
rect 9255 8450 9263 8486
rect 9212 8415 9263 8450
rect 9212 8379 9221 8415
rect 9255 8379 9263 8415
rect 9212 8344 9263 8379
rect 9212 8308 9221 8344
rect 9255 8308 9263 8344
rect 7123 8216 7277 8250
rect 7311 8216 7535 8250
rect 7569 8216 7793 8250
rect 7827 8216 8051 8250
rect 8085 8216 8309 8250
rect 8343 8216 8490 8250
rect 9076 8216 9092 8250
rect 9126 8216 9142 8250
rect 7123 8191 8490 8216
rect 7397 8172 7448 8191
rect 7914 8172 7965 8191
rect 8430 8172 8481 8191
rect 6529 8126 6859 8172
rect 9212 8159 9263 8308
rect 9470 8486 9521 8632
rect 9592 8544 9608 8578
rect 9642 8544 9658 8578
rect 9850 8544 9866 8578
rect 9900 8544 9916 8578
rect 9470 8450 9479 8486
rect 9513 8450 9521 8486
rect 9470 8415 9521 8450
rect 9470 8379 9479 8415
rect 9513 8379 9521 8415
rect 9470 8344 9521 8379
rect 9470 8308 9479 8344
rect 9513 8308 9521 8344
rect 9470 8277 9521 8308
rect 9729 8486 9780 8518
rect 9986 8503 10038 8632
rect 10749 8578 12108 8671
rect 10108 8544 10124 8578
rect 10158 8544 10174 8578
rect 10749 8544 10898 8578
rect 10932 8544 11156 8578
rect 11190 8544 11414 8578
rect 11448 8544 11672 8578
rect 11706 8544 11930 8578
rect 11964 8544 12108 8578
rect 9729 8450 9737 8486
rect 9771 8450 9780 8486
rect 9729 8415 9780 8450
rect 9729 8379 9737 8415
rect 9771 8379 9780 8415
rect 9729 8344 9780 8379
rect 9729 8308 9737 8344
rect 9771 8308 9780 8344
rect 9334 8216 9350 8250
rect 9384 8216 9400 8250
rect 9592 8216 9608 8250
rect 9642 8216 9658 8250
rect 9729 8160 9780 8308
rect 9987 8486 10038 8503
rect 9987 8450 9995 8486
rect 10029 8450 10038 8486
rect 9987 8415 10038 8450
rect 9987 8379 9995 8415
rect 10029 8379 10038 8415
rect 9987 8344 10038 8379
rect 9987 8308 9995 8344
rect 10029 8308 10038 8344
rect 9987 8277 10038 8308
rect 10245 8486 10296 8517
rect 10245 8450 10253 8486
rect 10287 8450 10296 8486
rect 10245 8415 10296 8450
rect 10245 8379 10253 8415
rect 10287 8379 10296 8415
rect 10245 8344 10296 8379
rect 10245 8308 10253 8344
rect 10287 8308 10296 8344
rect 9850 8216 9866 8250
rect 9900 8216 9916 8250
rect 10108 8216 10124 8250
rect 10158 8216 10174 8250
rect 9729 8159 9789 8160
rect 10245 8159 10296 8308
rect 9212 8052 10296 8159
rect 10749 8486 12108 8544
rect 10749 8450 10769 8486
rect 10803 8450 11027 8486
rect 11061 8450 11285 8486
rect 11319 8450 11543 8486
rect 11577 8450 11801 8486
rect 11835 8450 12059 8486
rect 12093 8450 12108 8486
rect 10749 8415 12108 8450
rect 10749 8379 10769 8415
rect 10803 8379 11027 8415
rect 11061 8379 11285 8415
rect 11319 8379 11543 8415
rect 11577 8379 11801 8415
rect 11835 8379 12059 8415
rect 12093 8379 12108 8415
rect 10749 8344 12108 8379
rect 10749 8308 10769 8344
rect 10803 8308 11027 8344
rect 11061 8308 11285 8344
rect 11319 8308 11543 8344
rect 11577 8308 11801 8344
rect 11835 8308 12059 8344
rect 12093 8308 12108 8344
rect 10749 8250 12108 8308
rect 10749 8216 10898 8250
rect 10932 8216 11156 8250
rect 11190 8216 11414 8250
rect 11448 8216 11672 8250
rect 11706 8216 11930 8250
rect 11964 8216 12108 8250
rect 10749 8109 12108 8216
rect 12846 8052 13168 8902
rect 14124 8668 17272 8902
rect 4498 8050 12508 8052
rect 12544 8050 13168 8052
rect 4498 7844 13168 8050
rect 4498 7842 4820 7844
rect 4508 7652 4670 7842
rect 4507 7638 4670 7652
rect 4507 7314 4669 7638
rect 5340 7612 5612 7642
rect 5692 7616 5756 7844
rect 8360 7652 8424 7844
rect 5340 7574 5436 7612
rect 5502 7574 5612 7612
rect 4512 6806 4662 7314
rect 5340 7488 5612 7574
rect 5340 7486 5544 7488
rect 5340 7450 5358 7486
rect 5396 7452 5544 7486
rect 5582 7452 5612 7488
rect 5396 7450 5612 7452
rect 5340 7414 5612 7450
rect 5693 7486 5755 7616
rect 6726 7612 6998 7642
rect 6072 7571 6088 7605
rect 6242 7571 6258 7605
rect 6726 7574 6822 7612
rect 6888 7574 6998 7612
rect 5693 7452 5719 7486
rect 5753 7452 5755 7486
rect 5693 7381 5755 7452
rect 6577 7486 6622 7502
rect 6611 7452 6622 7486
rect 6072 7333 6088 7367
rect 6242 7333 6258 7367
rect 6577 7224 6622 7452
rect 6726 7488 6998 7574
rect 6726 7486 6930 7488
rect 6726 7450 6744 7486
rect 6782 7452 6930 7486
rect 6968 7452 6998 7488
rect 6782 7450 6998 7452
rect 6726 7414 6998 7450
rect 7096 7612 7368 7642
rect 7096 7574 7192 7612
rect 7258 7574 7368 7612
rect 7096 7488 7368 7574
rect 7096 7486 7300 7488
rect 7096 7450 7114 7486
rect 7152 7452 7300 7486
rect 7338 7452 7368 7488
rect 7152 7450 7368 7452
rect 7096 7414 7368 7450
rect 7518 7612 7790 7642
rect 7518 7574 7614 7612
rect 7680 7574 7790 7612
rect 7518 7488 7790 7574
rect 7518 7486 7722 7488
rect 7518 7450 7536 7486
rect 7574 7452 7722 7486
rect 7760 7452 7790 7488
rect 7574 7450 7790 7452
rect 7518 7414 7790 7450
rect 7940 7612 8212 7642
rect 8360 7640 8425 7652
rect 7940 7574 8036 7612
rect 8102 7574 8212 7612
rect 7940 7488 8212 7574
rect 7940 7486 8144 7488
rect 7940 7450 7958 7486
rect 7996 7452 8144 7486
rect 8182 7452 8212 7488
rect 7996 7450 8212 7452
rect 7940 7414 8212 7450
rect 8363 7486 8425 7640
rect 9440 7612 9712 7642
rect 8742 7571 8758 7605
rect 8912 7571 8928 7605
rect 9440 7574 9536 7612
rect 9602 7574 9712 7612
rect 8363 7452 8389 7486
rect 8423 7452 8425 7486
rect 8363 7381 8425 7452
rect 9247 7486 9292 7502
rect 9281 7452 9292 7486
rect 8742 7333 8758 7367
rect 8912 7333 8928 7367
rect 9247 7242 9292 7452
rect 9440 7488 9712 7574
rect 9440 7486 9644 7488
rect 9440 7450 9458 7486
rect 9496 7452 9644 7486
rect 9682 7452 9712 7488
rect 9496 7450 9712 7452
rect 9440 7414 9712 7450
rect 9810 7612 10082 7642
rect 9810 7574 9906 7612
rect 9972 7574 10082 7612
rect 9810 7488 10082 7574
rect 9810 7486 10014 7488
rect 9810 7450 9828 7486
rect 9866 7452 10014 7486
rect 10052 7452 10082 7488
rect 9866 7450 10082 7452
rect 9810 7414 10082 7450
rect 10232 7612 10504 7642
rect 10232 7574 10328 7612
rect 10394 7574 10504 7612
rect 10232 7488 10504 7574
rect 10232 7486 10436 7488
rect 10232 7450 10250 7486
rect 10288 7452 10436 7486
rect 10474 7452 10504 7488
rect 10288 7450 10504 7452
rect 10232 7414 10504 7450
rect 10654 7612 10926 7642
rect 10654 7574 10750 7612
rect 10816 7574 10926 7612
rect 10654 7488 10926 7574
rect 10654 7486 10858 7488
rect 10654 7450 10672 7486
rect 10710 7452 10858 7486
rect 10896 7452 10926 7488
rect 10710 7450 10926 7452
rect 10654 7414 10926 7450
rect 11026 7624 11090 7844
rect 12090 7842 13168 7844
rect 12090 7840 12402 7842
rect 12846 7836 13168 7842
rect 13010 7644 13166 7836
rect 11026 7487 11088 7624
rect 12094 7612 12366 7642
rect 11405 7572 11421 7606
rect 11575 7572 11591 7606
rect 12094 7574 12190 7612
rect 12256 7574 12366 7612
rect 13010 7606 13167 7644
rect 11026 7453 11052 7487
rect 11086 7453 11088 7487
rect 11026 7382 11088 7453
rect 11910 7487 11955 7503
rect 11944 7453 11955 7487
rect 11405 7334 11421 7368
rect 11575 7334 11591 7368
rect 6576 7220 6622 7224
rect 4507 6697 4662 6806
rect 6576 6818 6621 7220
rect 9246 6818 9292 7242
rect 11910 7220 11955 7453
rect 12094 7488 12366 7574
rect 12094 7486 12298 7488
rect 12094 7450 12112 7486
rect 12150 7452 12298 7486
rect 12336 7452 12366 7488
rect 12150 7450 12366 7452
rect 12094 7414 12366 7450
rect 6576 6807 8917 6818
rect 6576 6728 8783 6807
rect 8878 6728 8917 6807
rect 6576 6713 8917 6728
rect 6576 6711 7247 6713
rect 8654 6712 8917 6713
rect 9246 6807 11575 6818
rect 9246 6728 11456 6807
rect 11551 6728 11575 6807
rect 9246 6713 11575 6728
rect 9246 6711 9922 6713
rect 11327 6712 11575 6713
rect 11909 6817 11955 7220
rect 13011 7215 13167 7606
rect 13015 7050 13165 7215
rect 12668 6920 12882 6966
rect 12668 6817 12692 6920
rect 11909 6742 12692 6817
rect 12860 6742 12882 6920
rect 11909 6712 12882 6742
rect 4512 2800 4662 6697
rect 5254 6575 5270 6609
rect 5304 6575 5320 6609
rect 5512 6575 5528 6609
rect 5562 6575 5578 6609
rect 5770 6575 5786 6609
rect 5820 6575 5836 6609
rect 6028 6575 6044 6609
rect 6078 6575 6094 6609
rect 6286 6575 6302 6609
rect 6336 6575 6352 6609
rect 6544 6575 6560 6609
rect 6594 6575 6610 6609
rect 6802 6575 6818 6609
rect 6852 6575 6868 6609
rect 7060 6575 7076 6609
rect 7110 6575 7126 6609
rect 5135 6525 5180 6569
rect 5135 6489 5141 6525
rect 5175 6489 5180 6525
rect 5135 6455 5180 6489
rect 5135 6419 5141 6455
rect 5175 6419 5180 6455
rect 5135 6385 5180 6419
rect 5135 6349 5141 6385
rect 5175 6349 5180 6385
rect 5135 6107 5180 6349
rect 5393 6525 5438 6569
rect 5393 6489 5399 6525
rect 5433 6489 5438 6525
rect 5393 6455 5438 6489
rect 5393 6419 5399 6455
rect 5433 6419 5438 6455
rect 5393 6385 5438 6419
rect 5393 6349 5399 6385
rect 5433 6349 5438 6385
rect 5254 6265 5270 6299
rect 5304 6265 5320 6299
rect 5254 6157 5270 6191
rect 5304 6157 5320 6191
rect 5135 6071 5141 6107
rect 5175 6071 5180 6107
rect 5135 6037 5180 6071
rect 5135 6001 5141 6037
rect 5175 6001 5180 6037
rect 5135 5967 5180 6001
rect 5135 5931 5141 5967
rect 5175 5931 5180 5967
rect 5135 5689 5180 5931
rect 5393 6107 5438 6349
rect 5650 6525 5695 6569
rect 5650 6489 5657 6525
rect 5691 6489 5695 6525
rect 5650 6455 5695 6489
rect 5650 6419 5657 6455
rect 5691 6419 5695 6455
rect 5650 6384 5695 6419
rect 5650 6348 5657 6384
rect 5691 6348 5695 6384
rect 5512 6265 5528 6299
rect 5562 6265 5578 6299
rect 5512 6157 5528 6191
rect 5562 6157 5578 6191
rect 5393 6071 5399 6107
rect 5433 6071 5438 6107
rect 5393 6037 5438 6071
rect 5393 6001 5399 6037
rect 5433 6001 5438 6037
rect 5393 5967 5438 6001
rect 5393 5931 5399 5967
rect 5433 5931 5438 5967
rect 5254 5847 5270 5881
rect 5304 5847 5320 5881
rect 5254 5739 5270 5773
rect 5304 5739 5320 5773
rect 5135 5653 5141 5689
rect 5175 5653 5180 5689
rect 5135 5619 5180 5653
rect 5135 5583 5141 5619
rect 5175 5583 5180 5619
rect 5135 5549 5180 5583
rect 5135 5513 5141 5549
rect 5175 5513 5180 5549
rect 5135 5271 5180 5513
rect 5393 5689 5438 5931
rect 5650 6107 5695 6348
rect 5910 6525 5955 6569
rect 5910 6489 5915 6525
rect 5949 6489 5955 6525
rect 5910 6455 5955 6489
rect 5910 6419 5915 6455
rect 5949 6419 5955 6455
rect 5910 6385 5955 6419
rect 5910 6349 5915 6385
rect 5949 6349 5955 6385
rect 5770 6265 5786 6299
rect 5820 6265 5836 6299
rect 5770 6157 5786 6191
rect 5820 6157 5836 6191
rect 5650 6071 5657 6107
rect 5691 6071 5695 6107
rect 5650 6037 5695 6071
rect 5650 6001 5657 6037
rect 5691 6001 5695 6037
rect 5650 5966 5695 6001
rect 5650 5930 5657 5966
rect 5691 5930 5695 5966
rect 5512 5847 5528 5881
rect 5562 5847 5578 5881
rect 5512 5739 5528 5773
rect 5562 5739 5578 5773
rect 5393 5653 5399 5689
rect 5433 5653 5438 5689
rect 5393 5619 5438 5653
rect 5393 5583 5399 5619
rect 5433 5583 5438 5619
rect 5393 5549 5438 5583
rect 5393 5513 5399 5549
rect 5433 5513 5438 5549
rect 5254 5429 5270 5463
rect 5304 5429 5320 5463
rect 5254 5321 5270 5355
rect 5304 5321 5320 5355
rect 5135 5235 5141 5271
rect 5175 5235 5180 5271
rect 5135 5201 5180 5235
rect 5135 5165 5141 5201
rect 5175 5165 5180 5201
rect 5135 5131 5180 5165
rect 5135 5095 5141 5131
rect 5175 5095 5180 5131
rect 5135 4853 5180 5095
rect 5393 5271 5438 5513
rect 5650 5689 5695 5930
rect 5910 6107 5955 6349
rect 6168 6525 6213 6569
rect 6168 6489 6173 6525
rect 6207 6489 6213 6525
rect 6168 6455 6213 6489
rect 6168 6419 6173 6455
rect 6207 6419 6213 6455
rect 6168 6385 6213 6419
rect 6168 6349 6173 6385
rect 6207 6349 6213 6385
rect 6028 6265 6044 6299
rect 6078 6265 6094 6299
rect 6028 6157 6044 6191
rect 6078 6157 6094 6191
rect 5910 6071 5915 6107
rect 5949 6071 5955 6107
rect 5910 6037 5955 6071
rect 5910 6001 5915 6037
rect 5949 6001 5955 6037
rect 5910 5967 5955 6001
rect 5910 5931 5915 5967
rect 5949 5931 5955 5967
rect 5770 5847 5786 5881
rect 5820 5847 5836 5881
rect 5770 5739 5786 5773
rect 5820 5739 5836 5773
rect 5650 5653 5657 5689
rect 5691 5653 5695 5689
rect 5650 5619 5695 5653
rect 5650 5583 5657 5619
rect 5691 5583 5695 5619
rect 5650 5548 5695 5583
rect 5650 5512 5657 5548
rect 5691 5512 5695 5548
rect 5512 5429 5528 5463
rect 5562 5429 5578 5463
rect 5512 5321 5528 5355
rect 5562 5321 5578 5355
rect 5393 5235 5399 5271
rect 5433 5235 5438 5271
rect 5393 5201 5438 5235
rect 5393 5165 5399 5201
rect 5433 5165 5438 5201
rect 5393 5131 5438 5165
rect 5393 5095 5399 5131
rect 5433 5095 5438 5131
rect 5254 5011 5270 5045
rect 5304 5011 5320 5045
rect 5254 4903 5270 4937
rect 5304 4903 5320 4937
rect 5135 4817 5141 4853
rect 5175 4817 5180 4853
rect 5135 4783 5180 4817
rect 5135 4747 5141 4783
rect 5175 4747 5180 4783
rect 5135 4713 5180 4747
rect 5135 4677 5141 4713
rect 5175 4677 5180 4713
rect 5135 4435 5180 4677
rect 5393 4853 5438 5095
rect 5650 5271 5695 5512
rect 5910 5689 5955 5931
rect 6168 6107 6213 6349
rect 6425 6525 6470 6569
rect 6425 6489 6431 6525
rect 6465 6489 6470 6525
rect 6425 6455 6470 6489
rect 6425 6419 6431 6455
rect 6465 6419 6470 6455
rect 6425 6385 6470 6419
rect 6425 6349 6431 6385
rect 6465 6349 6470 6385
rect 6286 6265 6302 6299
rect 6336 6265 6352 6299
rect 6286 6157 6302 6191
rect 6336 6157 6352 6191
rect 6168 6071 6173 6107
rect 6207 6071 6213 6107
rect 6168 6037 6213 6071
rect 6168 6001 6173 6037
rect 6207 6001 6213 6037
rect 6168 5967 6213 6001
rect 6168 5931 6173 5967
rect 6207 5931 6213 5967
rect 6028 5847 6044 5881
rect 6078 5847 6094 5881
rect 6028 5739 6044 5773
rect 6078 5739 6094 5773
rect 5910 5653 5915 5689
rect 5949 5653 5955 5689
rect 5910 5619 5955 5653
rect 5910 5583 5915 5619
rect 5949 5583 5955 5619
rect 5910 5549 5955 5583
rect 5910 5513 5915 5549
rect 5949 5513 5955 5549
rect 5770 5429 5786 5463
rect 5820 5429 5836 5463
rect 5770 5321 5786 5355
rect 5820 5321 5836 5355
rect 5650 5235 5657 5271
rect 5691 5235 5695 5271
rect 5650 5201 5695 5235
rect 5650 5165 5657 5201
rect 5691 5165 5695 5201
rect 5650 5130 5695 5165
rect 5650 5094 5657 5130
rect 5691 5094 5695 5130
rect 5512 5011 5528 5045
rect 5562 5011 5578 5045
rect 5512 4903 5528 4937
rect 5562 4903 5578 4937
rect 5393 4817 5399 4853
rect 5433 4817 5438 4853
rect 5393 4783 5438 4817
rect 5393 4747 5399 4783
rect 5433 4747 5438 4783
rect 5393 4713 5438 4747
rect 5393 4677 5399 4713
rect 5433 4677 5438 4713
rect 5254 4593 5270 4627
rect 5304 4593 5320 4627
rect 5254 4485 5270 4519
rect 5304 4485 5320 4519
rect 5135 4399 5141 4435
rect 5175 4399 5180 4435
rect 5135 4365 5180 4399
rect 5135 4329 5141 4365
rect 5175 4329 5180 4365
rect 5135 4295 5180 4329
rect 5135 4259 5141 4295
rect 5175 4259 5180 4295
rect 5135 4017 5180 4259
rect 5393 4435 5438 4677
rect 5650 4853 5695 5094
rect 5910 5271 5955 5513
rect 6168 5689 6213 5931
rect 6425 6107 6470 6349
rect 6682 6525 6727 6569
rect 6682 6489 6689 6525
rect 6723 6489 6727 6525
rect 6682 6455 6727 6489
rect 6682 6419 6689 6455
rect 6723 6419 6727 6455
rect 6682 6385 6727 6419
rect 6682 6349 6689 6385
rect 6723 6349 6727 6385
rect 6544 6265 6560 6299
rect 6594 6265 6610 6299
rect 6544 6157 6560 6191
rect 6594 6157 6610 6191
rect 6425 6071 6431 6107
rect 6465 6071 6470 6107
rect 6425 6037 6470 6071
rect 6425 6001 6431 6037
rect 6465 6001 6470 6037
rect 6425 5967 6470 6001
rect 6425 5931 6431 5967
rect 6465 5931 6470 5967
rect 6286 5847 6302 5881
rect 6336 5847 6352 5881
rect 6286 5739 6302 5773
rect 6336 5739 6352 5773
rect 6168 5653 6173 5689
rect 6207 5653 6213 5689
rect 6168 5619 6213 5653
rect 6168 5583 6173 5619
rect 6207 5583 6213 5619
rect 6168 5549 6213 5583
rect 6168 5513 6173 5549
rect 6207 5513 6213 5549
rect 6028 5429 6044 5463
rect 6078 5429 6094 5463
rect 6028 5321 6044 5355
rect 6078 5321 6094 5355
rect 5910 5235 5915 5271
rect 5949 5235 5955 5271
rect 5910 5201 5955 5235
rect 5910 5165 5915 5201
rect 5949 5165 5955 5201
rect 5910 5131 5955 5165
rect 5910 5095 5915 5131
rect 5949 5095 5955 5131
rect 5770 5011 5786 5045
rect 5820 5011 5836 5045
rect 5770 4903 5786 4937
rect 5820 4903 5836 4937
rect 5650 4817 5657 4853
rect 5691 4817 5695 4853
rect 5650 4783 5695 4817
rect 5650 4747 5657 4783
rect 5691 4747 5695 4783
rect 5650 4712 5695 4747
rect 5650 4676 5657 4712
rect 5691 4676 5695 4712
rect 5512 4593 5528 4627
rect 5562 4593 5578 4627
rect 5512 4485 5528 4519
rect 5562 4485 5578 4519
rect 5393 4399 5399 4435
rect 5433 4399 5438 4435
rect 5393 4365 5438 4399
rect 5393 4329 5399 4365
rect 5433 4329 5438 4365
rect 5393 4295 5438 4329
rect 5393 4259 5399 4295
rect 5433 4259 5438 4295
rect 5254 4175 5270 4209
rect 5304 4175 5320 4209
rect 5254 4067 5270 4101
rect 5304 4067 5320 4101
rect 5135 3981 5141 4017
rect 5175 3981 5180 4017
rect 5135 3947 5180 3981
rect 5135 3911 5141 3947
rect 5175 3911 5180 3947
rect 5135 3877 5180 3911
rect 5135 3841 5141 3877
rect 5175 3841 5180 3877
rect 5135 3599 5180 3841
rect 5393 4017 5438 4259
rect 5650 4435 5695 4676
rect 5910 4853 5955 5095
rect 6168 5271 6213 5513
rect 6425 5689 6470 5931
rect 6682 6107 6727 6349
rect 6941 6525 6986 6569
rect 6941 6489 6947 6525
rect 6981 6489 6986 6525
rect 6941 6455 6986 6489
rect 6941 6419 6947 6455
rect 6981 6419 6986 6455
rect 6941 6385 6986 6419
rect 6941 6349 6947 6385
rect 6981 6349 6986 6385
rect 6802 6265 6818 6299
rect 6852 6265 6868 6299
rect 6802 6157 6818 6191
rect 6852 6157 6868 6191
rect 6682 6071 6689 6107
rect 6723 6071 6727 6107
rect 6682 6037 6727 6071
rect 6682 6001 6689 6037
rect 6723 6001 6727 6037
rect 6682 5967 6727 6001
rect 6682 5931 6689 5967
rect 6723 5931 6727 5967
rect 6544 5847 6560 5881
rect 6594 5847 6610 5881
rect 6544 5739 6560 5773
rect 6594 5739 6610 5773
rect 6425 5653 6431 5689
rect 6465 5653 6470 5689
rect 6425 5619 6470 5653
rect 6425 5583 6431 5619
rect 6465 5583 6470 5619
rect 6425 5549 6470 5583
rect 6425 5513 6431 5549
rect 6465 5513 6470 5549
rect 6286 5429 6302 5463
rect 6336 5429 6352 5463
rect 6286 5321 6302 5355
rect 6336 5321 6352 5355
rect 6168 5235 6173 5271
rect 6207 5235 6213 5271
rect 6168 5201 6213 5235
rect 6168 5165 6173 5201
rect 6207 5165 6213 5201
rect 6168 5131 6213 5165
rect 6168 5095 6173 5131
rect 6207 5095 6213 5131
rect 6028 5011 6044 5045
rect 6078 5011 6094 5045
rect 6028 4903 6044 4937
rect 6078 4903 6094 4937
rect 5910 4817 5915 4853
rect 5949 4817 5955 4853
rect 5910 4783 5955 4817
rect 5910 4747 5915 4783
rect 5949 4747 5955 4783
rect 5910 4713 5955 4747
rect 5910 4677 5915 4713
rect 5949 4677 5955 4713
rect 5770 4593 5786 4627
rect 5820 4593 5836 4627
rect 5770 4485 5786 4519
rect 5820 4485 5836 4519
rect 5650 4399 5657 4435
rect 5691 4399 5695 4435
rect 5650 4365 5695 4399
rect 5650 4329 5657 4365
rect 5691 4329 5695 4365
rect 5650 4294 5695 4329
rect 5650 4258 5657 4294
rect 5691 4258 5695 4294
rect 5512 4175 5528 4209
rect 5562 4175 5578 4209
rect 5512 4067 5528 4101
rect 5562 4067 5578 4101
rect 5393 3981 5399 4017
rect 5433 3981 5438 4017
rect 5393 3947 5438 3981
rect 5393 3911 5399 3947
rect 5433 3911 5438 3947
rect 5393 3877 5438 3911
rect 5393 3841 5399 3877
rect 5433 3841 5438 3877
rect 5254 3757 5270 3791
rect 5304 3757 5320 3791
rect 5393 3723 5438 3841
rect 5650 4017 5695 4258
rect 5910 4435 5955 4677
rect 6168 4853 6213 5095
rect 6425 5271 6470 5513
rect 6682 5689 6727 5931
rect 6941 6107 6986 6349
rect 7199 6525 7244 6711
rect 7924 6575 7940 6609
rect 7974 6575 7990 6609
rect 8182 6575 8198 6609
rect 8232 6575 8248 6609
rect 8440 6575 8456 6609
rect 8490 6575 8506 6609
rect 8698 6575 8714 6609
rect 8748 6575 8764 6609
rect 8956 6575 8972 6609
rect 9006 6575 9022 6609
rect 9214 6575 9230 6609
rect 9264 6575 9280 6609
rect 9472 6575 9488 6609
rect 9522 6575 9538 6609
rect 9730 6575 9746 6609
rect 9780 6575 9796 6609
rect 7199 6489 7205 6525
rect 7239 6489 7244 6525
rect 7199 6455 7244 6489
rect 7199 6419 7205 6455
rect 7239 6419 7244 6455
rect 7199 6385 7244 6419
rect 7199 6349 7205 6385
rect 7239 6349 7244 6385
rect 7060 6265 7076 6299
rect 7110 6265 7126 6299
rect 7060 6157 7076 6191
rect 7110 6157 7126 6191
rect 6941 6071 6947 6107
rect 6981 6071 6986 6107
rect 6941 6037 6986 6071
rect 6941 6001 6947 6037
rect 6981 6001 6986 6037
rect 6941 5967 6986 6001
rect 6941 5931 6947 5967
rect 6981 5931 6986 5967
rect 6802 5847 6818 5881
rect 6852 5847 6868 5881
rect 6802 5739 6818 5773
rect 6852 5739 6868 5773
rect 6682 5653 6689 5689
rect 6723 5653 6727 5689
rect 6682 5619 6727 5653
rect 6682 5583 6689 5619
rect 6723 5583 6727 5619
rect 6682 5549 6727 5583
rect 6682 5513 6689 5549
rect 6723 5513 6727 5549
rect 6544 5429 6560 5463
rect 6594 5429 6610 5463
rect 6544 5321 6560 5355
rect 6594 5321 6610 5355
rect 6425 5235 6431 5271
rect 6465 5235 6470 5271
rect 6425 5201 6470 5235
rect 6425 5165 6431 5201
rect 6465 5165 6470 5201
rect 6425 5131 6470 5165
rect 6425 5095 6431 5131
rect 6465 5095 6470 5131
rect 6286 5011 6302 5045
rect 6336 5011 6352 5045
rect 6286 4903 6302 4937
rect 6336 4903 6352 4937
rect 6168 4817 6173 4853
rect 6207 4817 6213 4853
rect 6168 4783 6213 4817
rect 6168 4747 6173 4783
rect 6207 4747 6213 4783
rect 6168 4713 6213 4747
rect 6168 4677 6173 4713
rect 6207 4677 6213 4713
rect 6028 4593 6044 4627
rect 6078 4593 6094 4627
rect 6028 4485 6044 4519
rect 6078 4485 6094 4519
rect 5910 4399 5915 4435
rect 5949 4399 5955 4435
rect 5910 4365 5955 4399
rect 5910 4329 5915 4365
rect 5949 4329 5955 4365
rect 5910 4295 5955 4329
rect 5910 4259 5915 4295
rect 5949 4259 5955 4295
rect 5770 4175 5786 4209
rect 5820 4175 5836 4209
rect 5770 4067 5786 4101
rect 5820 4067 5836 4101
rect 5650 3981 5657 4017
rect 5691 3981 5695 4017
rect 5650 3947 5695 3981
rect 5650 3911 5657 3947
rect 5691 3911 5695 3947
rect 5650 3876 5695 3911
rect 5650 3840 5657 3876
rect 5691 3840 5695 3876
rect 5512 3757 5528 3791
rect 5562 3757 5578 3791
rect 5650 3723 5695 3840
rect 5910 4017 5955 4259
rect 6168 4435 6213 4677
rect 6425 4853 6470 5095
rect 6682 5271 6727 5513
rect 6941 5689 6986 5931
rect 7199 6107 7244 6349
rect 7199 6071 7205 6107
rect 7239 6071 7244 6107
rect 7199 6037 7244 6071
rect 7199 6001 7205 6037
rect 7239 6001 7244 6037
rect 7199 5967 7244 6001
rect 7199 5931 7205 5967
rect 7239 5931 7244 5967
rect 7060 5847 7076 5881
rect 7110 5847 7126 5881
rect 7060 5739 7076 5773
rect 7110 5739 7126 5773
rect 6941 5653 6947 5689
rect 6981 5653 6986 5689
rect 6941 5619 6986 5653
rect 6941 5583 6947 5619
rect 6981 5583 6986 5619
rect 6941 5549 6986 5583
rect 6941 5513 6947 5549
rect 6981 5513 6986 5549
rect 6802 5429 6818 5463
rect 6852 5429 6868 5463
rect 6802 5321 6818 5355
rect 6852 5321 6868 5355
rect 6682 5235 6689 5271
rect 6723 5235 6727 5271
rect 6682 5201 6727 5235
rect 6682 5165 6689 5201
rect 6723 5165 6727 5201
rect 6682 5131 6727 5165
rect 6682 5095 6689 5131
rect 6723 5095 6727 5131
rect 6544 5011 6560 5045
rect 6594 5011 6610 5045
rect 6544 4903 6560 4937
rect 6594 4903 6610 4937
rect 6425 4817 6431 4853
rect 6465 4817 6470 4853
rect 6425 4783 6470 4817
rect 6425 4747 6431 4783
rect 6465 4747 6470 4783
rect 6425 4713 6470 4747
rect 6425 4677 6431 4713
rect 6465 4677 6470 4713
rect 6286 4593 6302 4627
rect 6336 4593 6352 4627
rect 6286 4485 6302 4519
rect 6336 4485 6352 4519
rect 6168 4399 6173 4435
rect 6207 4399 6213 4435
rect 6168 4365 6213 4399
rect 6168 4329 6173 4365
rect 6207 4329 6213 4365
rect 6168 4295 6213 4329
rect 6168 4259 6173 4295
rect 6207 4259 6213 4295
rect 6028 4175 6044 4209
rect 6078 4175 6094 4209
rect 6028 4067 6044 4101
rect 6078 4067 6094 4101
rect 5910 3981 5915 4017
rect 5949 3981 5955 4017
rect 5910 3947 5955 3981
rect 5910 3911 5915 3947
rect 5949 3911 5955 3947
rect 5910 3877 5955 3911
rect 5910 3841 5915 3877
rect 5949 3841 5955 3877
rect 5770 3757 5786 3791
rect 5820 3757 5836 3791
rect 5910 3723 5955 3841
rect 6168 4017 6213 4259
rect 6425 4435 6470 4677
rect 6682 4853 6727 5095
rect 6941 5271 6986 5513
rect 7199 5689 7244 5931
rect 7199 5653 7205 5689
rect 7239 5653 7244 5689
rect 7199 5619 7244 5653
rect 7199 5583 7205 5619
rect 7239 5583 7244 5619
rect 7199 5549 7244 5583
rect 7199 5513 7205 5549
rect 7239 5513 7244 5549
rect 7060 5429 7076 5463
rect 7110 5429 7126 5463
rect 7060 5321 7076 5355
rect 7110 5321 7126 5355
rect 6941 5235 6947 5271
rect 6981 5235 6986 5271
rect 6941 5201 6986 5235
rect 6941 5165 6947 5201
rect 6981 5165 6986 5201
rect 6941 5131 6986 5165
rect 6941 5095 6947 5131
rect 6981 5095 6986 5131
rect 6802 5011 6818 5045
rect 6852 5011 6868 5045
rect 6802 4903 6818 4937
rect 6852 4903 6868 4937
rect 6682 4817 6689 4853
rect 6723 4817 6727 4853
rect 6682 4783 6727 4817
rect 6682 4747 6689 4783
rect 6723 4747 6727 4783
rect 6682 4713 6727 4747
rect 6682 4677 6689 4713
rect 6723 4677 6727 4713
rect 6544 4593 6560 4627
rect 6594 4593 6610 4627
rect 6544 4485 6560 4519
rect 6594 4485 6610 4519
rect 6425 4399 6431 4435
rect 6465 4399 6470 4435
rect 6425 4365 6470 4399
rect 6425 4329 6431 4365
rect 6465 4329 6470 4365
rect 6425 4295 6470 4329
rect 6425 4259 6431 4295
rect 6465 4259 6470 4295
rect 6286 4175 6302 4209
rect 6336 4175 6352 4209
rect 6286 4067 6302 4101
rect 6336 4067 6352 4101
rect 6168 3981 6173 4017
rect 6207 3981 6213 4017
rect 6168 3947 6213 3981
rect 6168 3911 6173 3947
rect 6207 3911 6213 3947
rect 6168 3877 6213 3911
rect 6168 3841 6173 3877
rect 6207 3841 6213 3877
rect 6028 3757 6044 3791
rect 6078 3757 6094 3791
rect 6168 3723 6213 3841
rect 6425 4017 6470 4259
rect 6682 4435 6727 4677
rect 6941 4853 6986 5095
rect 7199 5271 7244 5513
rect 7199 5235 7205 5271
rect 7239 5235 7244 5271
rect 7199 5201 7244 5235
rect 7199 5165 7205 5201
rect 7239 5165 7244 5201
rect 7199 5131 7244 5165
rect 7199 5095 7205 5131
rect 7239 5095 7244 5131
rect 7060 5011 7076 5045
rect 7110 5011 7126 5045
rect 7060 4903 7076 4937
rect 7110 4903 7126 4937
rect 6941 4817 6947 4853
rect 6981 4817 6986 4853
rect 6941 4783 6986 4817
rect 6941 4747 6947 4783
rect 6981 4747 6986 4783
rect 6941 4713 6986 4747
rect 6941 4677 6947 4713
rect 6981 4677 6986 4713
rect 6802 4593 6818 4627
rect 6852 4593 6868 4627
rect 6802 4485 6818 4519
rect 6852 4485 6868 4519
rect 6682 4399 6689 4435
rect 6723 4399 6727 4435
rect 6682 4365 6727 4399
rect 6682 4329 6689 4365
rect 6723 4329 6727 4365
rect 6682 4295 6727 4329
rect 6682 4259 6689 4295
rect 6723 4259 6727 4295
rect 6544 4175 6560 4209
rect 6594 4175 6610 4209
rect 6544 4067 6560 4101
rect 6594 4067 6610 4101
rect 6425 3981 6431 4017
rect 6465 3981 6470 4017
rect 6425 3947 6470 3981
rect 6425 3911 6431 3947
rect 6465 3911 6470 3947
rect 6425 3877 6470 3911
rect 6425 3841 6431 3877
rect 6465 3841 6470 3877
rect 6286 3757 6302 3791
rect 6336 3757 6352 3791
rect 6425 3723 6470 3841
rect 6682 4017 6727 4259
rect 6941 4435 6986 4677
rect 7199 4853 7244 5095
rect 7199 4817 7205 4853
rect 7239 4817 7244 4853
rect 7199 4783 7244 4817
rect 7199 4747 7205 4783
rect 7239 4747 7244 4783
rect 7199 4713 7244 4747
rect 7199 4677 7205 4713
rect 7239 4677 7244 4713
rect 7060 4593 7076 4627
rect 7110 4593 7126 4627
rect 7060 4485 7076 4519
rect 7110 4485 7126 4519
rect 6941 4399 6947 4435
rect 6981 4399 6986 4435
rect 6941 4365 6986 4399
rect 6941 4329 6947 4365
rect 6981 4329 6986 4365
rect 6941 4295 6986 4329
rect 6941 4259 6947 4295
rect 6981 4259 6986 4295
rect 6802 4175 6818 4209
rect 6852 4175 6868 4209
rect 6802 4067 6818 4101
rect 6852 4067 6868 4101
rect 6682 3981 6689 4017
rect 6723 3981 6727 4017
rect 6682 3947 6727 3981
rect 6682 3911 6689 3947
rect 6723 3911 6727 3947
rect 6682 3877 6727 3911
rect 6682 3841 6689 3877
rect 6723 3841 6727 3877
rect 6544 3757 6560 3791
rect 6594 3757 6610 3791
rect 6682 3723 6727 3841
rect 6941 4017 6986 4259
rect 7199 4435 7244 4677
rect 7199 4399 7205 4435
rect 7239 4399 7244 4435
rect 7199 4365 7244 4399
rect 7199 4329 7205 4365
rect 7239 4329 7244 4365
rect 7199 4295 7244 4329
rect 7199 4259 7205 4295
rect 7239 4259 7244 4295
rect 7060 4175 7076 4209
rect 7110 4175 7126 4209
rect 7060 4067 7076 4101
rect 7110 4067 7126 4101
rect 6941 3981 6947 4017
rect 6981 3981 6986 4017
rect 6941 3947 6986 3981
rect 6941 3911 6947 3947
rect 6981 3911 6986 3947
rect 6941 3877 6986 3911
rect 6941 3841 6947 3877
rect 6981 3841 6986 3877
rect 6802 3757 6818 3791
rect 6852 3757 6868 3791
rect 6941 3723 6986 3841
rect 7199 4017 7244 4259
rect 7199 3981 7205 4017
rect 7239 3981 7244 4017
rect 7199 3947 7244 3981
rect 7199 3911 7205 3947
rect 7239 3911 7244 3947
rect 7199 3877 7244 3911
rect 7199 3841 7205 3877
rect 7239 3841 7244 3877
rect 7060 3757 7076 3791
rect 7110 3757 7126 3791
rect 7199 3723 7244 3841
rect 7805 6525 7850 6569
rect 7805 6489 7811 6525
rect 7845 6489 7850 6525
rect 7805 6455 7850 6489
rect 7805 6419 7811 6455
rect 7845 6419 7850 6455
rect 7805 6385 7850 6419
rect 7805 6349 7811 6385
rect 7845 6349 7850 6385
rect 7805 6107 7850 6349
rect 8063 6525 8108 6569
rect 8063 6489 8069 6525
rect 8103 6489 8108 6525
rect 8063 6455 8108 6489
rect 8063 6419 8069 6455
rect 8103 6419 8108 6455
rect 8063 6385 8108 6419
rect 8063 6349 8069 6385
rect 8103 6349 8108 6385
rect 7924 6265 7940 6299
rect 7974 6265 7990 6299
rect 7924 6157 7940 6191
rect 7974 6157 7990 6191
rect 7805 6071 7811 6107
rect 7845 6071 7850 6107
rect 7805 6037 7850 6071
rect 7805 6001 7811 6037
rect 7845 6001 7850 6037
rect 7805 5967 7850 6001
rect 7805 5931 7811 5967
rect 7845 5931 7850 5967
rect 7805 5689 7850 5931
rect 8063 6107 8108 6349
rect 8320 6525 8365 6569
rect 8320 6489 8327 6525
rect 8361 6489 8365 6525
rect 8320 6455 8365 6489
rect 8320 6419 8327 6455
rect 8361 6419 8365 6455
rect 8320 6384 8365 6419
rect 8320 6348 8327 6384
rect 8361 6348 8365 6384
rect 8182 6265 8198 6299
rect 8232 6265 8248 6299
rect 8182 6157 8198 6191
rect 8232 6157 8248 6191
rect 8063 6071 8069 6107
rect 8103 6071 8108 6107
rect 8063 6037 8108 6071
rect 8063 6001 8069 6037
rect 8103 6001 8108 6037
rect 8063 5967 8108 6001
rect 8063 5931 8069 5967
rect 8103 5931 8108 5967
rect 7924 5847 7940 5881
rect 7974 5847 7990 5881
rect 7924 5739 7940 5773
rect 7974 5739 7990 5773
rect 7805 5653 7811 5689
rect 7845 5653 7850 5689
rect 7805 5619 7850 5653
rect 7805 5583 7811 5619
rect 7845 5583 7850 5619
rect 7805 5549 7850 5583
rect 7805 5513 7811 5549
rect 7845 5513 7850 5549
rect 7805 5271 7850 5513
rect 8063 5689 8108 5931
rect 8320 6107 8365 6348
rect 8580 6525 8625 6569
rect 8580 6489 8585 6525
rect 8619 6489 8625 6525
rect 8580 6455 8625 6489
rect 8580 6419 8585 6455
rect 8619 6419 8625 6455
rect 8580 6385 8625 6419
rect 8580 6349 8585 6385
rect 8619 6349 8625 6385
rect 8440 6265 8456 6299
rect 8490 6265 8506 6299
rect 8440 6157 8456 6191
rect 8490 6157 8506 6191
rect 8320 6071 8327 6107
rect 8361 6071 8365 6107
rect 8320 6037 8365 6071
rect 8320 6001 8327 6037
rect 8361 6001 8365 6037
rect 8320 5966 8365 6001
rect 8320 5930 8327 5966
rect 8361 5930 8365 5966
rect 8182 5847 8198 5881
rect 8232 5847 8248 5881
rect 8182 5739 8198 5773
rect 8232 5739 8248 5773
rect 8063 5653 8069 5689
rect 8103 5653 8108 5689
rect 8063 5619 8108 5653
rect 8063 5583 8069 5619
rect 8103 5583 8108 5619
rect 8063 5549 8108 5583
rect 8063 5513 8069 5549
rect 8103 5513 8108 5549
rect 7924 5429 7940 5463
rect 7974 5429 7990 5463
rect 7924 5321 7940 5355
rect 7974 5321 7990 5355
rect 7805 5235 7811 5271
rect 7845 5235 7850 5271
rect 7805 5201 7850 5235
rect 7805 5165 7811 5201
rect 7845 5165 7850 5201
rect 7805 5131 7850 5165
rect 7805 5095 7811 5131
rect 7845 5095 7850 5131
rect 7805 4853 7850 5095
rect 8063 5271 8108 5513
rect 8320 5689 8365 5930
rect 8580 6107 8625 6349
rect 8838 6525 8883 6569
rect 8838 6489 8843 6525
rect 8877 6489 8883 6525
rect 8838 6455 8883 6489
rect 8838 6419 8843 6455
rect 8877 6419 8883 6455
rect 8838 6385 8883 6419
rect 8838 6349 8843 6385
rect 8877 6349 8883 6385
rect 8698 6265 8714 6299
rect 8748 6265 8764 6299
rect 8698 6157 8714 6191
rect 8748 6157 8764 6191
rect 8580 6071 8585 6107
rect 8619 6071 8625 6107
rect 8580 6037 8625 6071
rect 8580 6001 8585 6037
rect 8619 6001 8625 6037
rect 8580 5967 8625 6001
rect 8580 5931 8585 5967
rect 8619 5931 8625 5967
rect 8440 5847 8456 5881
rect 8490 5847 8506 5881
rect 8440 5739 8456 5773
rect 8490 5739 8506 5773
rect 8320 5653 8327 5689
rect 8361 5653 8365 5689
rect 8320 5619 8365 5653
rect 8320 5583 8327 5619
rect 8361 5583 8365 5619
rect 8320 5548 8365 5583
rect 8320 5512 8327 5548
rect 8361 5512 8365 5548
rect 8182 5429 8198 5463
rect 8232 5429 8248 5463
rect 8182 5321 8198 5355
rect 8232 5321 8248 5355
rect 8063 5235 8069 5271
rect 8103 5235 8108 5271
rect 8063 5201 8108 5235
rect 8063 5165 8069 5201
rect 8103 5165 8108 5201
rect 8063 5131 8108 5165
rect 8063 5095 8069 5131
rect 8103 5095 8108 5131
rect 7924 5011 7940 5045
rect 7974 5011 7990 5045
rect 7924 4903 7940 4937
rect 7974 4903 7990 4937
rect 7805 4817 7811 4853
rect 7845 4817 7850 4853
rect 7805 4783 7850 4817
rect 7805 4747 7811 4783
rect 7845 4747 7850 4783
rect 7805 4713 7850 4747
rect 7805 4677 7811 4713
rect 7845 4677 7850 4713
rect 7805 4435 7850 4677
rect 8063 4853 8108 5095
rect 8320 5271 8365 5512
rect 8580 5689 8625 5931
rect 8838 6107 8883 6349
rect 9095 6525 9140 6569
rect 9095 6489 9101 6525
rect 9135 6489 9140 6525
rect 9095 6455 9140 6489
rect 9095 6419 9101 6455
rect 9135 6419 9140 6455
rect 9095 6385 9140 6419
rect 9095 6349 9101 6385
rect 9135 6349 9140 6385
rect 8956 6265 8972 6299
rect 9006 6265 9022 6299
rect 8956 6157 8972 6191
rect 9006 6157 9022 6191
rect 8838 6071 8843 6107
rect 8877 6071 8883 6107
rect 8838 6037 8883 6071
rect 8838 6001 8843 6037
rect 8877 6001 8883 6037
rect 8838 5967 8883 6001
rect 8838 5931 8843 5967
rect 8877 5931 8883 5967
rect 8698 5847 8714 5881
rect 8748 5847 8764 5881
rect 8698 5739 8714 5773
rect 8748 5739 8764 5773
rect 8580 5653 8585 5689
rect 8619 5653 8625 5689
rect 8580 5619 8625 5653
rect 8580 5583 8585 5619
rect 8619 5583 8625 5619
rect 8580 5549 8625 5583
rect 8580 5513 8585 5549
rect 8619 5513 8625 5549
rect 8440 5429 8456 5463
rect 8490 5429 8506 5463
rect 8440 5321 8456 5355
rect 8490 5321 8506 5355
rect 8320 5235 8327 5271
rect 8361 5235 8365 5271
rect 8320 5201 8365 5235
rect 8320 5165 8327 5201
rect 8361 5165 8365 5201
rect 8320 5130 8365 5165
rect 8320 5094 8327 5130
rect 8361 5094 8365 5130
rect 8182 5011 8198 5045
rect 8232 5011 8248 5045
rect 8182 4903 8198 4937
rect 8232 4903 8248 4937
rect 8063 4817 8069 4853
rect 8103 4817 8108 4853
rect 8063 4783 8108 4817
rect 8063 4747 8069 4783
rect 8103 4747 8108 4783
rect 8063 4713 8108 4747
rect 8063 4677 8069 4713
rect 8103 4677 8108 4713
rect 7924 4593 7940 4627
rect 7974 4593 7990 4627
rect 7924 4485 7940 4519
rect 7974 4485 7990 4519
rect 7805 4399 7811 4435
rect 7845 4399 7850 4435
rect 7805 4365 7850 4399
rect 7805 4329 7811 4365
rect 7845 4329 7850 4365
rect 7805 4295 7850 4329
rect 7805 4259 7811 4295
rect 7845 4259 7850 4295
rect 7805 4017 7850 4259
rect 8063 4435 8108 4677
rect 8320 4853 8365 5094
rect 8580 5271 8625 5513
rect 8838 5689 8883 5931
rect 9095 6107 9140 6349
rect 9352 6525 9397 6569
rect 9352 6489 9359 6525
rect 9393 6489 9397 6525
rect 9352 6455 9397 6489
rect 9352 6419 9359 6455
rect 9393 6419 9397 6455
rect 9352 6385 9397 6419
rect 9352 6349 9359 6385
rect 9393 6349 9397 6385
rect 9214 6265 9230 6299
rect 9264 6265 9280 6299
rect 9214 6157 9230 6191
rect 9264 6157 9280 6191
rect 9095 6071 9101 6107
rect 9135 6071 9140 6107
rect 9095 6037 9140 6071
rect 9095 6001 9101 6037
rect 9135 6001 9140 6037
rect 9095 5967 9140 6001
rect 9095 5931 9101 5967
rect 9135 5931 9140 5967
rect 8956 5847 8972 5881
rect 9006 5847 9022 5881
rect 8956 5739 8972 5773
rect 9006 5739 9022 5773
rect 8838 5653 8843 5689
rect 8877 5653 8883 5689
rect 8838 5619 8883 5653
rect 8838 5583 8843 5619
rect 8877 5583 8883 5619
rect 8838 5549 8883 5583
rect 8838 5513 8843 5549
rect 8877 5513 8883 5549
rect 8698 5429 8714 5463
rect 8748 5429 8764 5463
rect 8698 5321 8714 5355
rect 8748 5321 8764 5355
rect 8580 5235 8585 5271
rect 8619 5235 8625 5271
rect 8580 5201 8625 5235
rect 8580 5165 8585 5201
rect 8619 5165 8625 5201
rect 8580 5131 8625 5165
rect 8580 5095 8585 5131
rect 8619 5095 8625 5131
rect 8440 5011 8456 5045
rect 8490 5011 8506 5045
rect 8440 4903 8456 4937
rect 8490 4903 8506 4937
rect 8320 4817 8327 4853
rect 8361 4817 8365 4853
rect 8320 4783 8365 4817
rect 8320 4747 8327 4783
rect 8361 4747 8365 4783
rect 8320 4712 8365 4747
rect 8320 4676 8327 4712
rect 8361 4676 8365 4712
rect 8182 4593 8198 4627
rect 8232 4593 8248 4627
rect 8182 4485 8198 4519
rect 8232 4485 8248 4519
rect 8063 4399 8069 4435
rect 8103 4399 8108 4435
rect 8063 4365 8108 4399
rect 8063 4329 8069 4365
rect 8103 4329 8108 4365
rect 8063 4295 8108 4329
rect 8063 4259 8069 4295
rect 8103 4259 8108 4295
rect 7924 4175 7940 4209
rect 7974 4175 7990 4209
rect 7924 4067 7940 4101
rect 7974 4067 7990 4101
rect 7805 3981 7811 4017
rect 7845 3981 7850 4017
rect 7805 3947 7850 3981
rect 7805 3911 7811 3947
rect 7845 3911 7850 3947
rect 7805 3877 7850 3911
rect 7805 3841 7811 3877
rect 7845 3841 7850 3877
rect 7805 3599 7850 3841
rect 8063 4017 8108 4259
rect 8320 4435 8365 4676
rect 8580 4853 8625 5095
rect 8838 5271 8883 5513
rect 9095 5689 9140 5931
rect 9352 6107 9397 6349
rect 9611 6525 9656 6569
rect 9611 6489 9617 6525
rect 9651 6489 9656 6525
rect 9611 6455 9656 6489
rect 9611 6419 9617 6455
rect 9651 6419 9656 6455
rect 9611 6385 9656 6419
rect 9611 6349 9617 6385
rect 9651 6349 9656 6385
rect 9472 6265 9488 6299
rect 9522 6265 9538 6299
rect 9472 6157 9488 6191
rect 9522 6157 9538 6191
rect 9352 6071 9359 6107
rect 9393 6071 9397 6107
rect 9352 6037 9397 6071
rect 9352 6001 9359 6037
rect 9393 6001 9397 6037
rect 9352 5967 9397 6001
rect 9352 5931 9359 5967
rect 9393 5931 9397 5967
rect 9214 5847 9230 5881
rect 9264 5847 9280 5881
rect 9214 5739 9230 5773
rect 9264 5739 9280 5773
rect 9095 5653 9101 5689
rect 9135 5653 9140 5689
rect 9095 5619 9140 5653
rect 9095 5583 9101 5619
rect 9135 5583 9140 5619
rect 9095 5549 9140 5583
rect 9095 5513 9101 5549
rect 9135 5513 9140 5549
rect 8956 5429 8972 5463
rect 9006 5429 9022 5463
rect 8956 5321 8972 5355
rect 9006 5321 9022 5355
rect 8838 5235 8843 5271
rect 8877 5235 8883 5271
rect 8838 5201 8883 5235
rect 8838 5165 8843 5201
rect 8877 5165 8883 5201
rect 8838 5131 8883 5165
rect 8838 5095 8843 5131
rect 8877 5095 8883 5131
rect 8698 5011 8714 5045
rect 8748 5011 8764 5045
rect 8698 4903 8714 4937
rect 8748 4903 8764 4937
rect 8580 4817 8585 4853
rect 8619 4817 8625 4853
rect 8580 4783 8625 4817
rect 8580 4747 8585 4783
rect 8619 4747 8625 4783
rect 8580 4713 8625 4747
rect 8580 4677 8585 4713
rect 8619 4677 8625 4713
rect 8440 4593 8456 4627
rect 8490 4593 8506 4627
rect 8440 4485 8456 4519
rect 8490 4485 8506 4519
rect 8320 4399 8327 4435
rect 8361 4399 8365 4435
rect 8320 4365 8365 4399
rect 8320 4329 8327 4365
rect 8361 4329 8365 4365
rect 8320 4294 8365 4329
rect 8320 4258 8327 4294
rect 8361 4258 8365 4294
rect 8182 4175 8198 4209
rect 8232 4175 8248 4209
rect 8182 4067 8198 4101
rect 8232 4067 8248 4101
rect 8063 3981 8069 4017
rect 8103 3981 8108 4017
rect 8063 3947 8108 3981
rect 8063 3911 8069 3947
rect 8103 3911 8108 3947
rect 8063 3877 8108 3911
rect 8063 3841 8069 3877
rect 8103 3841 8108 3877
rect 7924 3757 7940 3791
rect 7974 3757 7990 3791
rect 8063 3723 8108 3841
rect 8320 4017 8365 4258
rect 8580 4435 8625 4677
rect 8838 4853 8883 5095
rect 9095 5271 9140 5513
rect 9352 5689 9397 5931
rect 9611 6107 9656 6349
rect 9869 6525 9914 6711
rect 12528 6710 12577 6712
rect 10587 6576 10603 6610
rect 10637 6576 10653 6610
rect 10845 6576 10861 6610
rect 10895 6576 10911 6610
rect 11103 6576 11119 6610
rect 11153 6576 11169 6610
rect 11361 6576 11377 6610
rect 11411 6576 11427 6610
rect 11619 6576 11635 6610
rect 11669 6576 11685 6610
rect 11877 6576 11893 6610
rect 11927 6576 11943 6610
rect 12135 6576 12151 6610
rect 12185 6576 12201 6610
rect 12393 6576 12409 6610
rect 12443 6576 12459 6610
rect 9869 6489 9875 6525
rect 9909 6489 9914 6525
rect 9869 6455 9914 6489
rect 9869 6419 9875 6455
rect 9909 6419 9914 6455
rect 9869 6385 9914 6419
rect 9869 6349 9875 6385
rect 9909 6349 9914 6385
rect 9730 6265 9746 6299
rect 9780 6265 9796 6299
rect 9730 6157 9746 6191
rect 9780 6157 9796 6191
rect 9611 6071 9617 6107
rect 9651 6071 9656 6107
rect 9611 6037 9656 6071
rect 9611 6001 9617 6037
rect 9651 6001 9656 6037
rect 9611 5967 9656 6001
rect 9611 5931 9617 5967
rect 9651 5931 9656 5967
rect 9472 5847 9488 5881
rect 9522 5847 9538 5881
rect 9472 5739 9488 5773
rect 9522 5739 9538 5773
rect 9352 5653 9359 5689
rect 9393 5653 9397 5689
rect 9352 5619 9397 5653
rect 9352 5583 9359 5619
rect 9393 5583 9397 5619
rect 9352 5549 9397 5583
rect 9352 5513 9359 5549
rect 9393 5513 9397 5549
rect 9214 5429 9230 5463
rect 9264 5429 9280 5463
rect 9214 5321 9230 5355
rect 9264 5321 9280 5355
rect 9095 5235 9101 5271
rect 9135 5235 9140 5271
rect 9095 5201 9140 5235
rect 9095 5165 9101 5201
rect 9135 5165 9140 5201
rect 9095 5131 9140 5165
rect 9095 5095 9101 5131
rect 9135 5095 9140 5131
rect 8956 5011 8972 5045
rect 9006 5011 9022 5045
rect 8956 4903 8972 4937
rect 9006 4903 9022 4937
rect 8838 4817 8843 4853
rect 8877 4817 8883 4853
rect 8838 4783 8883 4817
rect 8838 4747 8843 4783
rect 8877 4747 8883 4783
rect 8838 4713 8883 4747
rect 8838 4677 8843 4713
rect 8877 4677 8883 4713
rect 8698 4593 8714 4627
rect 8748 4593 8764 4627
rect 8698 4485 8714 4519
rect 8748 4485 8764 4519
rect 8580 4399 8585 4435
rect 8619 4399 8625 4435
rect 8580 4365 8625 4399
rect 8580 4329 8585 4365
rect 8619 4329 8625 4365
rect 8580 4295 8625 4329
rect 8580 4259 8585 4295
rect 8619 4259 8625 4295
rect 8440 4175 8456 4209
rect 8490 4175 8506 4209
rect 8440 4067 8456 4101
rect 8490 4067 8506 4101
rect 8320 3981 8327 4017
rect 8361 3981 8365 4017
rect 8320 3947 8365 3981
rect 8320 3911 8327 3947
rect 8361 3911 8365 3947
rect 8320 3876 8365 3911
rect 8320 3840 8327 3876
rect 8361 3840 8365 3876
rect 8182 3757 8198 3791
rect 8232 3757 8248 3791
rect 8320 3723 8365 3840
rect 8580 4017 8625 4259
rect 8838 4435 8883 4677
rect 9095 4853 9140 5095
rect 9352 5271 9397 5513
rect 9611 5689 9656 5931
rect 9869 6107 9914 6349
rect 9869 6071 9875 6107
rect 9909 6071 9914 6107
rect 9869 6037 9914 6071
rect 9869 6001 9875 6037
rect 9909 6001 9914 6037
rect 9869 5967 9914 6001
rect 9869 5931 9875 5967
rect 9909 5931 9914 5967
rect 9730 5847 9746 5881
rect 9780 5847 9796 5881
rect 9730 5739 9746 5773
rect 9780 5739 9796 5773
rect 9611 5653 9617 5689
rect 9651 5653 9656 5689
rect 9611 5619 9656 5653
rect 9611 5583 9617 5619
rect 9651 5583 9656 5619
rect 9611 5549 9656 5583
rect 9611 5513 9617 5549
rect 9651 5513 9656 5549
rect 9472 5429 9488 5463
rect 9522 5429 9538 5463
rect 9472 5321 9488 5355
rect 9522 5321 9538 5355
rect 9352 5235 9359 5271
rect 9393 5235 9397 5271
rect 9352 5201 9397 5235
rect 9352 5165 9359 5201
rect 9393 5165 9397 5201
rect 9352 5131 9397 5165
rect 9352 5095 9359 5131
rect 9393 5095 9397 5131
rect 9214 5011 9230 5045
rect 9264 5011 9280 5045
rect 9214 4903 9230 4937
rect 9264 4903 9280 4937
rect 9095 4817 9101 4853
rect 9135 4817 9140 4853
rect 9095 4783 9140 4817
rect 9095 4747 9101 4783
rect 9135 4747 9140 4783
rect 9095 4713 9140 4747
rect 9095 4677 9101 4713
rect 9135 4677 9140 4713
rect 8956 4593 8972 4627
rect 9006 4593 9022 4627
rect 8956 4485 8972 4519
rect 9006 4485 9022 4519
rect 8838 4399 8843 4435
rect 8877 4399 8883 4435
rect 8838 4365 8883 4399
rect 8838 4329 8843 4365
rect 8877 4329 8883 4365
rect 8838 4295 8883 4329
rect 8838 4259 8843 4295
rect 8877 4259 8883 4295
rect 8698 4175 8714 4209
rect 8748 4175 8764 4209
rect 8698 4067 8714 4101
rect 8748 4067 8764 4101
rect 8580 3981 8585 4017
rect 8619 3981 8625 4017
rect 8580 3947 8625 3981
rect 8580 3911 8585 3947
rect 8619 3911 8625 3947
rect 8580 3877 8625 3911
rect 8580 3841 8585 3877
rect 8619 3841 8625 3877
rect 8440 3757 8456 3791
rect 8490 3757 8506 3791
rect 8580 3723 8625 3841
rect 8838 4017 8883 4259
rect 9095 4435 9140 4677
rect 9352 4853 9397 5095
rect 9611 5271 9656 5513
rect 9869 5689 9914 5931
rect 9869 5653 9875 5689
rect 9909 5653 9914 5689
rect 9869 5619 9914 5653
rect 9869 5583 9875 5619
rect 9909 5583 9914 5619
rect 9869 5549 9914 5583
rect 9869 5513 9875 5549
rect 9909 5513 9914 5549
rect 9730 5429 9746 5463
rect 9780 5429 9796 5463
rect 9730 5321 9746 5355
rect 9780 5321 9796 5355
rect 9611 5235 9617 5271
rect 9651 5235 9656 5271
rect 9611 5201 9656 5235
rect 9611 5165 9617 5201
rect 9651 5165 9656 5201
rect 9611 5131 9656 5165
rect 9611 5095 9617 5131
rect 9651 5095 9656 5131
rect 9472 5011 9488 5045
rect 9522 5011 9538 5045
rect 9472 4903 9488 4937
rect 9522 4903 9538 4937
rect 9352 4817 9359 4853
rect 9393 4817 9397 4853
rect 9352 4783 9397 4817
rect 9352 4747 9359 4783
rect 9393 4747 9397 4783
rect 9352 4713 9397 4747
rect 9352 4677 9359 4713
rect 9393 4677 9397 4713
rect 9214 4593 9230 4627
rect 9264 4593 9280 4627
rect 9214 4485 9230 4519
rect 9264 4485 9280 4519
rect 9095 4399 9101 4435
rect 9135 4399 9140 4435
rect 9095 4365 9140 4399
rect 9095 4329 9101 4365
rect 9135 4329 9140 4365
rect 9095 4295 9140 4329
rect 9095 4259 9101 4295
rect 9135 4259 9140 4295
rect 8956 4175 8972 4209
rect 9006 4175 9022 4209
rect 8956 4067 8972 4101
rect 9006 4067 9022 4101
rect 8838 3981 8843 4017
rect 8877 3981 8883 4017
rect 8838 3947 8883 3981
rect 8838 3911 8843 3947
rect 8877 3911 8883 3947
rect 8838 3877 8883 3911
rect 8838 3841 8843 3877
rect 8877 3841 8883 3877
rect 8698 3757 8714 3791
rect 8748 3757 8764 3791
rect 8838 3723 8883 3841
rect 9095 4017 9140 4259
rect 9352 4435 9397 4677
rect 9611 4853 9656 5095
rect 9869 5271 9914 5513
rect 9869 5235 9875 5271
rect 9909 5235 9914 5271
rect 9869 5201 9914 5235
rect 9869 5165 9875 5201
rect 9909 5165 9914 5201
rect 9869 5131 9914 5165
rect 9869 5095 9875 5131
rect 9909 5095 9914 5131
rect 9730 5011 9746 5045
rect 9780 5011 9796 5045
rect 9730 4903 9746 4937
rect 9780 4903 9796 4937
rect 9611 4817 9617 4853
rect 9651 4817 9656 4853
rect 9611 4783 9656 4817
rect 9611 4747 9617 4783
rect 9651 4747 9656 4783
rect 9611 4713 9656 4747
rect 9611 4677 9617 4713
rect 9651 4677 9656 4713
rect 9472 4593 9488 4627
rect 9522 4593 9538 4627
rect 9472 4485 9488 4519
rect 9522 4485 9538 4519
rect 9352 4399 9359 4435
rect 9393 4399 9397 4435
rect 9352 4365 9397 4399
rect 9352 4329 9359 4365
rect 9393 4329 9397 4365
rect 9352 4295 9397 4329
rect 9352 4259 9359 4295
rect 9393 4259 9397 4295
rect 9214 4175 9230 4209
rect 9264 4175 9280 4209
rect 9214 4067 9230 4101
rect 9264 4067 9280 4101
rect 9095 3981 9101 4017
rect 9135 3981 9140 4017
rect 9095 3947 9140 3981
rect 9095 3911 9101 3947
rect 9135 3911 9140 3947
rect 9095 3877 9140 3911
rect 9095 3841 9101 3877
rect 9135 3841 9140 3877
rect 8956 3757 8972 3791
rect 9006 3757 9022 3791
rect 9095 3723 9140 3841
rect 9352 4017 9397 4259
rect 9611 4435 9656 4677
rect 9869 4853 9914 5095
rect 9869 4817 9875 4853
rect 9909 4817 9914 4853
rect 9869 4783 9914 4817
rect 9869 4747 9875 4783
rect 9909 4747 9914 4783
rect 9869 4713 9914 4747
rect 9869 4677 9875 4713
rect 9909 4677 9914 4713
rect 9730 4593 9746 4627
rect 9780 4593 9796 4627
rect 9730 4485 9746 4519
rect 9780 4485 9796 4519
rect 9611 4399 9617 4435
rect 9651 4399 9656 4435
rect 9611 4365 9656 4399
rect 9611 4329 9617 4365
rect 9651 4329 9656 4365
rect 9611 4295 9656 4329
rect 9611 4259 9617 4295
rect 9651 4259 9656 4295
rect 9472 4175 9488 4209
rect 9522 4175 9538 4209
rect 9472 4067 9488 4101
rect 9522 4067 9538 4101
rect 9352 3981 9359 4017
rect 9393 3981 9397 4017
rect 9352 3947 9397 3981
rect 9352 3911 9359 3947
rect 9393 3911 9397 3947
rect 9352 3877 9397 3911
rect 9352 3841 9359 3877
rect 9393 3841 9397 3877
rect 9214 3757 9230 3791
rect 9264 3757 9280 3791
rect 9352 3723 9397 3841
rect 9611 4017 9656 4259
rect 9869 4435 9914 4677
rect 9869 4399 9875 4435
rect 9909 4399 9914 4435
rect 9869 4365 9914 4399
rect 9869 4329 9875 4365
rect 9909 4329 9914 4365
rect 9869 4295 9914 4329
rect 9869 4259 9875 4295
rect 9909 4259 9914 4295
rect 9730 4175 9746 4209
rect 9780 4175 9796 4209
rect 9730 4067 9746 4101
rect 9780 4067 9796 4101
rect 9611 3981 9617 4017
rect 9651 3981 9656 4017
rect 9611 3947 9656 3981
rect 9611 3911 9617 3947
rect 9651 3911 9656 3947
rect 9611 3877 9656 3911
rect 9611 3841 9617 3877
rect 9651 3841 9656 3877
rect 9472 3757 9488 3791
rect 9522 3757 9538 3791
rect 9611 3723 9656 3841
rect 9869 4017 9914 4259
rect 9869 3981 9875 4017
rect 9909 3981 9914 4017
rect 9869 3947 9914 3981
rect 9869 3911 9875 3947
rect 9909 3911 9914 3947
rect 9869 3877 9914 3911
rect 9869 3841 9875 3877
rect 9909 3841 9914 3877
rect 9730 3757 9746 3791
rect 9780 3757 9796 3791
rect 9869 3723 9914 3841
rect 10468 6526 10513 6570
rect 10468 6490 10474 6526
rect 10508 6490 10513 6526
rect 10468 6456 10513 6490
rect 10468 6420 10474 6456
rect 10508 6420 10513 6456
rect 10468 6386 10513 6420
rect 10468 6350 10474 6386
rect 10508 6350 10513 6386
rect 10468 6108 10513 6350
rect 10726 6526 10771 6570
rect 10726 6490 10732 6526
rect 10766 6490 10771 6526
rect 10726 6456 10771 6490
rect 10726 6420 10732 6456
rect 10766 6420 10771 6456
rect 10726 6386 10771 6420
rect 10726 6350 10732 6386
rect 10766 6350 10771 6386
rect 10587 6266 10603 6300
rect 10637 6266 10653 6300
rect 10587 6158 10603 6192
rect 10637 6158 10653 6192
rect 10468 6072 10474 6108
rect 10508 6072 10513 6108
rect 10468 6038 10513 6072
rect 10468 6002 10474 6038
rect 10508 6002 10513 6038
rect 10468 5968 10513 6002
rect 10468 5932 10474 5968
rect 10508 5932 10513 5968
rect 10468 5690 10513 5932
rect 10726 6108 10771 6350
rect 10983 6526 11028 6570
rect 10983 6490 10990 6526
rect 11024 6490 11028 6526
rect 10983 6456 11028 6490
rect 10983 6420 10990 6456
rect 11024 6420 11028 6456
rect 10983 6385 11028 6420
rect 10983 6349 10990 6385
rect 11024 6349 11028 6385
rect 10845 6266 10861 6300
rect 10895 6266 10911 6300
rect 10845 6158 10861 6192
rect 10895 6158 10911 6192
rect 10726 6072 10732 6108
rect 10766 6072 10771 6108
rect 10726 6038 10771 6072
rect 10726 6002 10732 6038
rect 10766 6002 10771 6038
rect 10726 5968 10771 6002
rect 10726 5932 10732 5968
rect 10766 5932 10771 5968
rect 10587 5848 10603 5882
rect 10637 5848 10653 5882
rect 10587 5740 10603 5774
rect 10637 5740 10653 5774
rect 10468 5654 10474 5690
rect 10508 5654 10513 5690
rect 10468 5620 10513 5654
rect 10468 5584 10474 5620
rect 10508 5584 10513 5620
rect 10468 5550 10513 5584
rect 10468 5514 10474 5550
rect 10508 5514 10513 5550
rect 10468 5272 10513 5514
rect 10726 5690 10771 5932
rect 10983 6108 11028 6349
rect 11243 6526 11288 6570
rect 11243 6490 11248 6526
rect 11282 6490 11288 6526
rect 11243 6456 11288 6490
rect 11243 6420 11248 6456
rect 11282 6420 11288 6456
rect 11243 6386 11288 6420
rect 11243 6350 11248 6386
rect 11282 6350 11288 6386
rect 11103 6266 11119 6300
rect 11153 6266 11169 6300
rect 11103 6158 11119 6192
rect 11153 6158 11169 6192
rect 10983 6072 10990 6108
rect 11024 6072 11028 6108
rect 10983 6038 11028 6072
rect 10983 6002 10990 6038
rect 11024 6002 11028 6038
rect 10983 5967 11028 6002
rect 10983 5931 10990 5967
rect 11024 5931 11028 5967
rect 10845 5848 10861 5882
rect 10895 5848 10911 5882
rect 10845 5740 10861 5774
rect 10895 5740 10911 5774
rect 10726 5654 10732 5690
rect 10766 5654 10771 5690
rect 10726 5620 10771 5654
rect 10726 5584 10732 5620
rect 10766 5584 10771 5620
rect 10726 5550 10771 5584
rect 10726 5514 10732 5550
rect 10766 5514 10771 5550
rect 10587 5430 10603 5464
rect 10637 5430 10653 5464
rect 10587 5322 10603 5356
rect 10637 5322 10653 5356
rect 10468 5236 10474 5272
rect 10508 5236 10513 5272
rect 10468 5202 10513 5236
rect 10468 5166 10474 5202
rect 10508 5166 10513 5202
rect 10468 5132 10513 5166
rect 10468 5096 10474 5132
rect 10508 5096 10513 5132
rect 10468 4854 10513 5096
rect 10726 5272 10771 5514
rect 10983 5690 11028 5931
rect 11243 6108 11288 6350
rect 11501 6526 11546 6570
rect 11501 6490 11506 6526
rect 11540 6490 11546 6526
rect 11501 6456 11546 6490
rect 11501 6420 11506 6456
rect 11540 6420 11546 6456
rect 11501 6386 11546 6420
rect 11501 6350 11506 6386
rect 11540 6350 11546 6386
rect 11361 6266 11377 6300
rect 11411 6266 11427 6300
rect 11361 6158 11377 6192
rect 11411 6158 11427 6192
rect 11243 6072 11248 6108
rect 11282 6072 11288 6108
rect 11243 6038 11288 6072
rect 11243 6002 11248 6038
rect 11282 6002 11288 6038
rect 11243 5968 11288 6002
rect 11243 5932 11248 5968
rect 11282 5932 11288 5968
rect 11103 5848 11119 5882
rect 11153 5848 11169 5882
rect 11103 5740 11119 5774
rect 11153 5740 11169 5774
rect 10983 5654 10990 5690
rect 11024 5654 11028 5690
rect 10983 5620 11028 5654
rect 10983 5584 10990 5620
rect 11024 5584 11028 5620
rect 10983 5549 11028 5584
rect 10983 5513 10990 5549
rect 11024 5513 11028 5549
rect 10845 5430 10861 5464
rect 10895 5430 10911 5464
rect 10845 5322 10861 5356
rect 10895 5322 10911 5356
rect 10726 5236 10732 5272
rect 10766 5236 10771 5272
rect 10726 5202 10771 5236
rect 10726 5166 10732 5202
rect 10766 5166 10771 5202
rect 10726 5132 10771 5166
rect 10726 5096 10732 5132
rect 10766 5096 10771 5132
rect 10587 5012 10603 5046
rect 10637 5012 10653 5046
rect 10587 4904 10603 4938
rect 10637 4904 10653 4938
rect 10468 4818 10474 4854
rect 10508 4818 10513 4854
rect 10468 4784 10513 4818
rect 10468 4748 10474 4784
rect 10508 4748 10513 4784
rect 10468 4714 10513 4748
rect 10468 4678 10474 4714
rect 10508 4678 10513 4714
rect 10468 4436 10513 4678
rect 10726 4854 10771 5096
rect 10983 5272 11028 5513
rect 11243 5690 11288 5932
rect 11501 6108 11546 6350
rect 11758 6526 11803 6570
rect 11758 6490 11764 6526
rect 11798 6490 11803 6526
rect 11758 6456 11803 6490
rect 11758 6420 11764 6456
rect 11798 6420 11803 6456
rect 11758 6386 11803 6420
rect 11758 6350 11764 6386
rect 11798 6350 11803 6386
rect 11619 6266 11635 6300
rect 11669 6266 11685 6300
rect 11619 6158 11635 6192
rect 11669 6158 11685 6192
rect 11501 6072 11506 6108
rect 11540 6072 11546 6108
rect 11501 6038 11546 6072
rect 11501 6002 11506 6038
rect 11540 6002 11546 6038
rect 11501 5968 11546 6002
rect 11501 5932 11506 5968
rect 11540 5932 11546 5968
rect 11361 5848 11377 5882
rect 11411 5848 11427 5882
rect 11361 5740 11377 5774
rect 11411 5740 11427 5774
rect 11243 5654 11248 5690
rect 11282 5654 11288 5690
rect 11243 5620 11288 5654
rect 11243 5584 11248 5620
rect 11282 5584 11288 5620
rect 11243 5550 11288 5584
rect 11243 5514 11248 5550
rect 11282 5514 11288 5550
rect 11103 5430 11119 5464
rect 11153 5430 11169 5464
rect 11103 5322 11119 5356
rect 11153 5322 11169 5356
rect 10983 5236 10990 5272
rect 11024 5236 11028 5272
rect 10983 5202 11028 5236
rect 10983 5166 10990 5202
rect 11024 5166 11028 5202
rect 10983 5131 11028 5166
rect 10983 5095 10990 5131
rect 11024 5095 11028 5131
rect 10845 5012 10861 5046
rect 10895 5012 10911 5046
rect 10845 4904 10861 4938
rect 10895 4904 10911 4938
rect 10726 4818 10732 4854
rect 10766 4818 10771 4854
rect 10726 4784 10771 4818
rect 10726 4748 10732 4784
rect 10766 4748 10771 4784
rect 10726 4714 10771 4748
rect 10726 4678 10732 4714
rect 10766 4678 10771 4714
rect 10587 4594 10603 4628
rect 10637 4594 10653 4628
rect 10587 4486 10603 4520
rect 10637 4486 10653 4520
rect 10468 4400 10474 4436
rect 10508 4400 10513 4436
rect 10468 4366 10513 4400
rect 10468 4330 10474 4366
rect 10508 4330 10513 4366
rect 10468 4296 10513 4330
rect 10468 4260 10474 4296
rect 10508 4260 10513 4296
rect 10468 4018 10513 4260
rect 10726 4436 10771 4678
rect 10983 4854 11028 5095
rect 11243 5272 11288 5514
rect 11501 5690 11546 5932
rect 11758 6108 11803 6350
rect 12015 6526 12060 6570
rect 12015 6490 12022 6526
rect 12056 6490 12060 6526
rect 12015 6456 12060 6490
rect 12015 6420 12022 6456
rect 12056 6420 12060 6456
rect 12015 6386 12060 6420
rect 12015 6350 12022 6386
rect 12056 6350 12060 6386
rect 11877 6266 11893 6300
rect 11927 6266 11943 6300
rect 11877 6158 11893 6192
rect 11927 6158 11943 6192
rect 11758 6072 11764 6108
rect 11798 6072 11803 6108
rect 11758 6038 11803 6072
rect 11758 6002 11764 6038
rect 11798 6002 11803 6038
rect 11758 5968 11803 6002
rect 11758 5932 11764 5968
rect 11798 5932 11803 5968
rect 11619 5848 11635 5882
rect 11669 5848 11685 5882
rect 11619 5740 11635 5774
rect 11669 5740 11685 5774
rect 11501 5654 11506 5690
rect 11540 5654 11546 5690
rect 11501 5620 11546 5654
rect 11501 5584 11506 5620
rect 11540 5584 11546 5620
rect 11501 5550 11546 5584
rect 11501 5514 11506 5550
rect 11540 5514 11546 5550
rect 11361 5430 11377 5464
rect 11411 5430 11427 5464
rect 11361 5322 11377 5356
rect 11411 5322 11427 5356
rect 11243 5236 11248 5272
rect 11282 5236 11288 5272
rect 11243 5202 11288 5236
rect 11243 5166 11248 5202
rect 11282 5166 11288 5202
rect 11243 5132 11288 5166
rect 11243 5096 11248 5132
rect 11282 5096 11288 5132
rect 11103 5012 11119 5046
rect 11153 5012 11169 5046
rect 11103 4904 11119 4938
rect 11153 4904 11169 4938
rect 10983 4818 10990 4854
rect 11024 4818 11028 4854
rect 10983 4784 11028 4818
rect 10983 4748 10990 4784
rect 11024 4748 11028 4784
rect 10983 4713 11028 4748
rect 10983 4677 10990 4713
rect 11024 4677 11028 4713
rect 10845 4594 10861 4628
rect 10895 4594 10911 4628
rect 10845 4486 10861 4520
rect 10895 4486 10911 4520
rect 10726 4400 10732 4436
rect 10766 4400 10771 4436
rect 10726 4366 10771 4400
rect 10726 4330 10732 4366
rect 10766 4330 10771 4366
rect 10726 4296 10771 4330
rect 10726 4260 10732 4296
rect 10766 4260 10771 4296
rect 10587 4176 10603 4210
rect 10637 4176 10653 4210
rect 10587 4068 10603 4102
rect 10637 4068 10653 4102
rect 10468 3982 10474 4018
rect 10508 3982 10513 4018
rect 10468 3948 10513 3982
rect 10468 3912 10474 3948
rect 10508 3912 10513 3948
rect 10468 3878 10513 3912
rect 10468 3842 10474 3878
rect 10508 3842 10513 3878
rect 10468 3600 10513 3842
rect 10726 4018 10771 4260
rect 10983 4436 11028 4677
rect 11243 4854 11288 5096
rect 11501 5272 11546 5514
rect 11758 5690 11803 5932
rect 12015 6108 12060 6350
rect 12274 6526 12319 6570
rect 12274 6490 12280 6526
rect 12314 6490 12319 6526
rect 12274 6456 12319 6490
rect 12274 6420 12280 6456
rect 12314 6420 12319 6456
rect 12274 6386 12319 6420
rect 12274 6350 12280 6386
rect 12314 6350 12319 6386
rect 12135 6266 12151 6300
rect 12185 6266 12201 6300
rect 12135 6158 12151 6192
rect 12185 6158 12201 6192
rect 12015 6072 12022 6108
rect 12056 6072 12060 6108
rect 12015 6038 12060 6072
rect 12015 6002 12022 6038
rect 12056 6002 12060 6038
rect 12015 5968 12060 6002
rect 12015 5932 12022 5968
rect 12056 5932 12060 5968
rect 11877 5848 11893 5882
rect 11927 5848 11943 5882
rect 11877 5740 11893 5774
rect 11927 5740 11943 5774
rect 11758 5654 11764 5690
rect 11798 5654 11803 5690
rect 11758 5620 11803 5654
rect 11758 5584 11764 5620
rect 11798 5584 11803 5620
rect 11758 5550 11803 5584
rect 11758 5514 11764 5550
rect 11798 5514 11803 5550
rect 11619 5430 11635 5464
rect 11669 5430 11685 5464
rect 11619 5322 11635 5356
rect 11669 5322 11685 5356
rect 11501 5236 11506 5272
rect 11540 5236 11546 5272
rect 11501 5202 11546 5236
rect 11501 5166 11506 5202
rect 11540 5166 11546 5202
rect 11501 5132 11546 5166
rect 11501 5096 11506 5132
rect 11540 5096 11546 5132
rect 11361 5012 11377 5046
rect 11411 5012 11427 5046
rect 11361 4904 11377 4938
rect 11411 4904 11427 4938
rect 11243 4818 11248 4854
rect 11282 4818 11288 4854
rect 11243 4784 11288 4818
rect 11243 4748 11248 4784
rect 11282 4748 11288 4784
rect 11243 4714 11288 4748
rect 11243 4678 11248 4714
rect 11282 4678 11288 4714
rect 11103 4594 11119 4628
rect 11153 4594 11169 4628
rect 11103 4486 11119 4520
rect 11153 4486 11169 4520
rect 10983 4400 10990 4436
rect 11024 4400 11028 4436
rect 10983 4366 11028 4400
rect 10983 4330 10990 4366
rect 11024 4330 11028 4366
rect 10983 4295 11028 4330
rect 10983 4259 10990 4295
rect 11024 4259 11028 4295
rect 10845 4176 10861 4210
rect 10895 4176 10911 4210
rect 10845 4068 10861 4102
rect 10895 4068 10911 4102
rect 10726 3982 10732 4018
rect 10766 3982 10771 4018
rect 10726 3948 10771 3982
rect 10726 3912 10732 3948
rect 10766 3912 10771 3948
rect 10726 3878 10771 3912
rect 10726 3842 10732 3878
rect 10766 3842 10771 3878
rect 10587 3758 10603 3792
rect 10637 3758 10653 3792
rect 10726 3724 10771 3842
rect 10983 4018 11028 4259
rect 11243 4436 11288 4678
rect 11501 4854 11546 5096
rect 11758 5272 11803 5514
rect 12015 5690 12060 5932
rect 12274 6108 12319 6350
rect 12532 6526 12577 6710
rect 13014 6684 13166 7050
rect 12532 6490 12538 6526
rect 12572 6490 12577 6526
rect 12532 6456 12577 6490
rect 12532 6420 12538 6456
rect 12572 6420 12577 6456
rect 12532 6386 12577 6420
rect 12532 6350 12538 6386
rect 12572 6350 12577 6386
rect 12393 6266 12409 6300
rect 12443 6266 12459 6300
rect 12393 6158 12409 6192
rect 12443 6158 12459 6192
rect 12274 6072 12280 6108
rect 12314 6072 12319 6108
rect 12274 6038 12319 6072
rect 12274 6002 12280 6038
rect 12314 6002 12319 6038
rect 12274 5968 12319 6002
rect 12274 5932 12280 5968
rect 12314 5932 12319 5968
rect 12135 5848 12151 5882
rect 12185 5848 12201 5882
rect 12135 5740 12151 5774
rect 12185 5740 12201 5774
rect 12015 5654 12022 5690
rect 12056 5654 12060 5690
rect 12015 5620 12060 5654
rect 12015 5584 12022 5620
rect 12056 5584 12060 5620
rect 12015 5550 12060 5584
rect 12015 5514 12022 5550
rect 12056 5514 12060 5550
rect 11877 5430 11893 5464
rect 11927 5430 11943 5464
rect 11877 5322 11893 5356
rect 11927 5322 11943 5356
rect 11758 5236 11764 5272
rect 11798 5236 11803 5272
rect 11758 5202 11803 5236
rect 11758 5166 11764 5202
rect 11798 5166 11803 5202
rect 11758 5132 11803 5166
rect 11758 5096 11764 5132
rect 11798 5096 11803 5132
rect 11619 5012 11635 5046
rect 11669 5012 11685 5046
rect 11619 4904 11635 4938
rect 11669 4904 11685 4938
rect 11501 4818 11506 4854
rect 11540 4818 11546 4854
rect 11501 4784 11546 4818
rect 11501 4748 11506 4784
rect 11540 4748 11546 4784
rect 11501 4714 11546 4748
rect 11501 4678 11506 4714
rect 11540 4678 11546 4714
rect 11361 4594 11377 4628
rect 11411 4594 11427 4628
rect 11361 4486 11377 4520
rect 11411 4486 11427 4520
rect 11243 4400 11248 4436
rect 11282 4400 11288 4436
rect 11243 4366 11288 4400
rect 11243 4330 11248 4366
rect 11282 4330 11288 4366
rect 11243 4296 11288 4330
rect 11243 4260 11248 4296
rect 11282 4260 11288 4296
rect 11103 4176 11119 4210
rect 11153 4176 11169 4210
rect 11103 4068 11119 4102
rect 11153 4068 11169 4102
rect 10983 3982 10990 4018
rect 11024 3982 11028 4018
rect 10983 3948 11028 3982
rect 10983 3912 10990 3948
rect 11024 3912 11028 3948
rect 10983 3877 11028 3912
rect 10983 3841 10990 3877
rect 11024 3841 11028 3877
rect 10845 3758 10861 3792
rect 10895 3758 10911 3792
rect 10983 3724 11028 3841
rect 11243 4018 11288 4260
rect 11501 4436 11546 4678
rect 11758 4854 11803 5096
rect 12015 5272 12060 5514
rect 12274 5690 12319 5932
rect 12532 6108 12577 6350
rect 12532 6072 12538 6108
rect 12572 6072 12577 6108
rect 12532 6038 12577 6072
rect 12532 6002 12538 6038
rect 12572 6002 12577 6038
rect 12532 5968 12577 6002
rect 12532 5932 12538 5968
rect 12572 5932 12577 5968
rect 12393 5848 12409 5882
rect 12443 5848 12459 5882
rect 12393 5740 12409 5774
rect 12443 5740 12459 5774
rect 12274 5654 12280 5690
rect 12314 5654 12319 5690
rect 12274 5620 12319 5654
rect 12274 5584 12280 5620
rect 12314 5584 12319 5620
rect 12274 5550 12319 5584
rect 12274 5514 12280 5550
rect 12314 5514 12319 5550
rect 12135 5430 12151 5464
rect 12185 5430 12201 5464
rect 12135 5322 12151 5356
rect 12185 5322 12201 5356
rect 12015 5236 12022 5272
rect 12056 5236 12060 5272
rect 12015 5202 12060 5236
rect 12015 5166 12022 5202
rect 12056 5166 12060 5202
rect 12015 5132 12060 5166
rect 12015 5096 12022 5132
rect 12056 5096 12060 5132
rect 11877 5012 11893 5046
rect 11927 5012 11943 5046
rect 11877 4904 11893 4938
rect 11927 4904 11943 4938
rect 11758 4818 11764 4854
rect 11798 4818 11803 4854
rect 11758 4784 11803 4818
rect 11758 4748 11764 4784
rect 11798 4748 11803 4784
rect 11758 4714 11803 4748
rect 11758 4678 11764 4714
rect 11798 4678 11803 4714
rect 11619 4594 11635 4628
rect 11669 4594 11685 4628
rect 11619 4486 11635 4520
rect 11669 4486 11685 4520
rect 11501 4400 11506 4436
rect 11540 4400 11546 4436
rect 11501 4366 11546 4400
rect 11501 4330 11506 4366
rect 11540 4330 11546 4366
rect 11501 4296 11546 4330
rect 11501 4260 11506 4296
rect 11540 4260 11546 4296
rect 11361 4176 11377 4210
rect 11411 4176 11427 4210
rect 11361 4068 11377 4102
rect 11411 4068 11427 4102
rect 11243 3982 11248 4018
rect 11282 3982 11288 4018
rect 11243 3948 11288 3982
rect 11243 3912 11248 3948
rect 11282 3912 11288 3948
rect 11243 3878 11288 3912
rect 11243 3842 11248 3878
rect 11282 3842 11288 3878
rect 11103 3758 11119 3792
rect 11153 3758 11169 3792
rect 11243 3724 11288 3842
rect 11501 4018 11546 4260
rect 11758 4436 11803 4678
rect 12015 4854 12060 5096
rect 12274 5272 12319 5514
rect 12532 5690 12577 5932
rect 12532 5654 12538 5690
rect 12572 5654 12577 5690
rect 12532 5620 12577 5654
rect 12532 5584 12538 5620
rect 12572 5584 12577 5620
rect 12532 5550 12577 5584
rect 12532 5514 12538 5550
rect 12572 5514 12577 5550
rect 12393 5430 12409 5464
rect 12443 5430 12459 5464
rect 12393 5322 12409 5356
rect 12443 5322 12459 5356
rect 12274 5236 12280 5272
rect 12314 5236 12319 5272
rect 12274 5202 12319 5236
rect 12274 5166 12280 5202
rect 12314 5166 12319 5202
rect 12274 5132 12319 5166
rect 12274 5096 12280 5132
rect 12314 5096 12319 5132
rect 12135 5012 12151 5046
rect 12185 5012 12201 5046
rect 12135 4904 12151 4938
rect 12185 4904 12201 4938
rect 12015 4818 12022 4854
rect 12056 4818 12060 4854
rect 12015 4784 12060 4818
rect 12015 4748 12022 4784
rect 12056 4748 12060 4784
rect 12015 4714 12060 4748
rect 12015 4678 12022 4714
rect 12056 4678 12060 4714
rect 11877 4594 11893 4628
rect 11927 4594 11943 4628
rect 11877 4486 11893 4520
rect 11927 4486 11943 4520
rect 11758 4400 11764 4436
rect 11798 4400 11803 4436
rect 11758 4366 11803 4400
rect 11758 4330 11764 4366
rect 11798 4330 11803 4366
rect 11758 4296 11803 4330
rect 11758 4260 11764 4296
rect 11798 4260 11803 4296
rect 11619 4176 11635 4210
rect 11669 4176 11685 4210
rect 11619 4068 11635 4102
rect 11669 4068 11685 4102
rect 11501 3982 11506 4018
rect 11540 3982 11546 4018
rect 11501 3948 11546 3982
rect 11501 3912 11506 3948
rect 11540 3912 11546 3948
rect 11501 3878 11546 3912
rect 11501 3842 11506 3878
rect 11540 3842 11546 3878
rect 11361 3758 11377 3792
rect 11411 3758 11427 3792
rect 11501 3724 11546 3842
rect 11758 4018 11803 4260
rect 12015 4436 12060 4678
rect 12274 4854 12319 5096
rect 12532 5272 12577 5514
rect 12532 5236 12538 5272
rect 12572 5236 12577 5272
rect 12532 5202 12577 5236
rect 12532 5166 12538 5202
rect 12572 5166 12577 5202
rect 12532 5132 12577 5166
rect 12532 5096 12538 5132
rect 12572 5096 12577 5132
rect 12393 5012 12409 5046
rect 12443 5012 12459 5046
rect 12393 4904 12409 4938
rect 12443 4904 12459 4938
rect 12274 4818 12280 4854
rect 12314 4818 12319 4854
rect 12274 4784 12319 4818
rect 12274 4748 12280 4784
rect 12314 4748 12319 4784
rect 12274 4714 12319 4748
rect 12274 4678 12280 4714
rect 12314 4678 12319 4714
rect 12135 4594 12151 4628
rect 12185 4594 12201 4628
rect 12135 4486 12151 4520
rect 12185 4486 12201 4520
rect 12015 4400 12022 4436
rect 12056 4400 12060 4436
rect 12015 4366 12060 4400
rect 12015 4330 12022 4366
rect 12056 4330 12060 4366
rect 12015 4296 12060 4330
rect 12015 4260 12022 4296
rect 12056 4260 12060 4296
rect 11877 4176 11893 4210
rect 11927 4176 11943 4210
rect 11877 4068 11893 4102
rect 11927 4068 11943 4102
rect 11758 3982 11764 4018
rect 11798 3982 11803 4018
rect 11758 3948 11803 3982
rect 11758 3912 11764 3948
rect 11798 3912 11803 3948
rect 11758 3878 11803 3912
rect 11758 3842 11764 3878
rect 11798 3842 11803 3878
rect 11619 3758 11635 3792
rect 11669 3758 11685 3792
rect 11758 3724 11803 3842
rect 12015 4018 12060 4260
rect 12274 4436 12319 4678
rect 12532 4854 12577 5096
rect 12532 4818 12538 4854
rect 12572 4818 12577 4854
rect 12532 4784 12577 4818
rect 12532 4748 12538 4784
rect 12572 4748 12577 4784
rect 12532 4714 12577 4748
rect 12532 4678 12538 4714
rect 12572 4678 12577 4714
rect 12393 4594 12409 4628
rect 12443 4594 12459 4628
rect 12393 4486 12409 4520
rect 12443 4486 12459 4520
rect 12274 4400 12280 4436
rect 12314 4400 12319 4436
rect 12274 4366 12319 4400
rect 12274 4330 12280 4366
rect 12314 4330 12319 4366
rect 12274 4296 12319 4330
rect 12274 4260 12280 4296
rect 12314 4260 12319 4296
rect 12135 4176 12151 4210
rect 12185 4176 12201 4210
rect 12135 4068 12151 4102
rect 12185 4068 12201 4102
rect 12015 3982 12022 4018
rect 12056 3982 12060 4018
rect 12015 3948 12060 3982
rect 12015 3912 12022 3948
rect 12056 3912 12060 3948
rect 12015 3878 12060 3912
rect 12015 3842 12022 3878
rect 12056 3842 12060 3878
rect 11877 3758 11893 3792
rect 11927 3758 11943 3792
rect 12015 3724 12060 3842
rect 12274 4018 12319 4260
rect 12532 4436 12577 4678
rect 12532 4400 12538 4436
rect 12572 4400 12577 4436
rect 12532 4366 12577 4400
rect 12532 4330 12538 4366
rect 12572 4330 12577 4366
rect 12532 4296 12577 4330
rect 12532 4260 12538 4296
rect 12572 4260 12577 4296
rect 12393 4176 12409 4210
rect 12443 4176 12459 4210
rect 12393 4068 12409 4102
rect 12443 4068 12459 4102
rect 12274 3982 12280 4018
rect 12314 3982 12319 4018
rect 12274 3948 12319 3982
rect 12274 3912 12280 3948
rect 12314 3912 12319 3948
rect 12274 3878 12319 3912
rect 12274 3842 12280 3878
rect 12314 3842 12319 3878
rect 12135 3758 12151 3792
rect 12185 3758 12201 3792
rect 12274 3724 12319 3842
rect 12532 4018 12577 4260
rect 12532 3982 12538 4018
rect 12572 3982 12577 4018
rect 12532 3948 12577 3982
rect 12532 3912 12538 3948
rect 12572 3912 12577 3948
rect 12532 3878 12577 3912
rect 12532 3842 12538 3878
rect 12572 3842 12577 3878
rect 12393 3758 12409 3792
rect 12443 3758 12459 3792
rect 12532 3724 12577 3842
rect 5135 3504 6361 3599
rect 7805 3504 9031 3599
rect 10468 3505 11694 3600
rect 5134 3415 5150 3449
rect 5184 3415 5200 3449
rect 5674 3415 5690 3449
rect 5724 3415 5740 3449
rect 6154 3415 6165 3449
rect 6215 3415 6220 3449
rect 4995 3363 5057 3385
rect 4995 3329 5021 3363
rect 5055 3329 5057 3363
rect 4995 3295 5057 3329
rect 4995 3259 5021 3295
rect 5055 3259 5057 3295
rect 4995 3225 5057 3259
rect 4995 3191 5021 3225
rect 5055 3191 5057 3225
rect 4995 3149 5057 3191
rect 5273 3363 5341 3383
rect 5273 3329 5279 3363
rect 5313 3329 5341 3363
rect 5273 3295 5341 3329
rect 5273 3259 5279 3295
rect 5313 3259 5341 3295
rect 5273 3225 5341 3259
rect 5273 3191 5279 3225
rect 5313 3191 5341 3225
rect 5273 3147 5341 3191
rect 5535 3363 5597 3385
rect 5535 3329 5561 3363
rect 5595 3329 5597 3363
rect 5535 3295 5597 3329
rect 5535 3259 5561 3295
rect 5595 3259 5597 3295
rect 5535 3225 5597 3259
rect 5535 3191 5561 3225
rect 5595 3191 5597 3225
rect 5535 3149 5597 3191
rect 5813 3363 5881 3383
rect 5813 3329 5819 3363
rect 5853 3329 5881 3363
rect 5813 3295 5881 3329
rect 5813 3259 5819 3295
rect 5853 3259 5881 3295
rect 5813 3225 5881 3259
rect 5813 3191 5819 3225
rect 5853 3191 5881 3225
rect 5813 3147 5881 3191
rect 6015 3363 6077 3385
rect 6015 3329 6041 3363
rect 6075 3329 6077 3363
rect 6015 3295 6077 3329
rect 6015 3259 6041 3295
rect 6075 3259 6077 3295
rect 6015 3225 6077 3259
rect 6015 3191 6041 3225
rect 6075 3191 6077 3225
rect 5134 3105 5150 3139
rect 5184 3105 5200 3139
rect 5674 3105 5690 3139
rect 5724 3105 5740 3139
rect 6015 3020 6077 3191
rect 6293 3363 6361 3504
rect 6657 3417 6673 3451
rect 6707 3417 6723 3451
rect 7167 3427 7183 3461
rect 7217 3427 7233 3461
rect 7804 3415 7820 3449
rect 7854 3415 7870 3449
rect 8344 3415 8360 3449
rect 8394 3415 8410 3449
rect 8824 3415 8835 3449
rect 8885 3415 8890 3449
rect 6293 3329 6299 3363
rect 6333 3329 6361 3363
rect 6293 3295 6361 3329
rect 6293 3259 6299 3295
rect 6333 3259 6361 3295
rect 6293 3225 6361 3259
rect 6293 3191 6299 3225
rect 6333 3191 6361 3225
rect 6293 3147 6361 3191
rect 6518 3365 6580 3387
rect 6518 3331 6544 3365
rect 6578 3331 6580 3365
rect 6518 3297 6580 3331
rect 6518 3261 6544 3297
rect 6578 3261 6580 3297
rect 6518 3227 6580 3261
rect 6518 3193 6544 3227
rect 6578 3193 6580 3227
rect 6518 3151 6580 3193
rect 6796 3365 6864 3385
rect 6796 3331 6802 3365
rect 6836 3331 6864 3365
rect 6796 3297 6864 3331
rect 6796 3261 6802 3297
rect 6836 3261 6864 3297
rect 6796 3227 6864 3261
rect 6796 3193 6802 3227
rect 6836 3193 6864 3227
rect 6796 3149 6864 3193
rect 7028 3375 7090 3397
rect 7028 3341 7054 3375
rect 7088 3341 7090 3375
rect 7028 3307 7090 3341
rect 7028 3271 7054 3307
rect 7088 3271 7090 3307
rect 7028 3237 7090 3271
rect 7028 3203 7054 3237
rect 7088 3203 7090 3237
rect 7028 3161 7090 3203
rect 7306 3375 7374 3395
rect 7306 3341 7312 3375
rect 7346 3341 7374 3375
rect 7306 3307 7374 3341
rect 7306 3271 7312 3307
rect 7346 3271 7374 3307
rect 7306 3237 7374 3271
rect 7306 3203 7312 3237
rect 7346 3203 7374 3237
rect 7306 3159 7374 3203
rect 7665 3363 7727 3385
rect 7665 3329 7691 3363
rect 7725 3329 7727 3363
rect 7665 3295 7727 3329
rect 7665 3259 7691 3295
rect 7725 3259 7727 3295
rect 7665 3225 7727 3259
rect 7665 3191 7691 3225
rect 7725 3191 7727 3225
rect 6154 3105 6168 3139
rect 6206 3105 6220 3139
rect 6657 3107 6673 3141
rect 6707 3107 6723 3141
rect 7167 3117 7183 3151
rect 7217 3117 7233 3151
rect 7665 3149 7727 3191
rect 7943 3363 8011 3383
rect 7943 3329 7949 3363
rect 7983 3329 8011 3363
rect 7943 3295 8011 3329
rect 7943 3259 7949 3295
rect 7983 3259 8011 3295
rect 7943 3225 8011 3259
rect 7943 3191 7949 3225
rect 7983 3191 8011 3225
rect 7943 3147 8011 3191
rect 8205 3363 8267 3385
rect 8205 3329 8231 3363
rect 8265 3329 8267 3363
rect 8205 3295 8267 3329
rect 8205 3259 8231 3295
rect 8265 3259 8267 3295
rect 8205 3225 8267 3259
rect 8205 3191 8231 3225
rect 8265 3191 8267 3225
rect 8205 3149 8267 3191
rect 8483 3363 8551 3383
rect 8483 3329 8489 3363
rect 8523 3329 8551 3363
rect 8483 3295 8551 3329
rect 8483 3259 8489 3295
rect 8523 3259 8551 3295
rect 8483 3225 8551 3259
rect 8483 3191 8489 3225
rect 8523 3191 8551 3225
rect 8483 3147 8551 3191
rect 8685 3363 8747 3385
rect 8685 3329 8711 3363
rect 8745 3329 8747 3363
rect 8685 3295 8747 3329
rect 8685 3259 8711 3295
rect 8745 3259 8747 3295
rect 8685 3225 8747 3259
rect 8685 3191 8711 3225
rect 8745 3191 8747 3225
rect 7804 3105 7820 3139
rect 7854 3105 7870 3139
rect 8344 3105 8360 3139
rect 8394 3105 8410 3139
rect 8685 3079 8747 3191
rect 8963 3363 9031 3504
rect 9327 3417 9343 3451
rect 9377 3417 9393 3451
rect 9837 3427 9853 3461
rect 9887 3427 9903 3461
rect 10467 3416 10483 3450
rect 10517 3416 10533 3450
rect 11007 3416 11023 3450
rect 11057 3416 11073 3450
rect 11487 3416 11498 3450
rect 11548 3416 11553 3450
rect 8963 3329 8969 3363
rect 9003 3329 9031 3363
rect 8963 3295 9031 3329
rect 8963 3259 8969 3295
rect 9003 3259 9031 3295
rect 8963 3225 9031 3259
rect 8963 3191 8969 3225
rect 9003 3191 9031 3225
rect 8963 3147 9031 3191
rect 9188 3365 9250 3387
rect 9188 3331 9214 3365
rect 9248 3331 9250 3365
rect 9188 3297 9250 3331
rect 9188 3261 9214 3297
rect 9248 3261 9250 3297
rect 9188 3227 9250 3261
rect 9188 3193 9214 3227
rect 9248 3193 9250 3227
rect 9188 3151 9250 3193
rect 9466 3365 9534 3385
rect 9466 3331 9472 3365
rect 9506 3331 9534 3365
rect 9466 3297 9534 3331
rect 9466 3261 9472 3297
rect 9506 3261 9534 3297
rect 9466 3227 9534 3261
rect 9466 3193 9472 3227
rect 9506 3193 9534 3227
rect 9466 3149 9534 3193
rect 9698 3375 9760 3397
rect 9698 3341 9724 3375
rect 9758 3341 9760 3375
rect 9698 3307 9760 3341
rect 9698 3271 9724 3307
rect 9758 3271 9760 3307
rect 9698 3237 9760 3271
rect 9698 3203 9724 3237
rect 9758 3203 9760 3237
rect 9698 3161 9760 3203
rect 9976 3375 10044 3395
rect 9976 3341 9982 3375
rect 10016 3341 10044 3375
rect 9976 3307 10044 3341
rect 9976 3271 9982 3307
rect 10016 3271 10044 3307
rect 9976 3237 10044 3271
rect 9976 3203 9982 3237
rect 10016 3203 10044 3237
rect 9976 3159 10044 3203
rect 10328 3364 10390 3386
rect 10328 3330 10354 3364
rect 10388 3330 10390 3364
rect 10328 3296 10390 3330
rect 10328 3260 10354 3296
rect 10388 3260 10390 3296
rect 10328 3226 10390 3260
rect 10328 3192 10354 3226
rect 10388 3192 10390 3226
rect 8824 3105 8838 3139
rect 8876 3105 8890 3139
rect 9327 3107 9343 3141
rect 9377 3107 9393 3141
rect 9837 3117 9853 3151
rect 9887 3117 9903 3151
rect 10328 3150 10390 3192
rect 10606 3364 10674 3384
rect 10606 3330 10612 3364
rect 10646 3330 10674 3364
rect 10606 3296 10674 3330
rect 10606 3260 10612 3296
rect 10646 3260 10674 3296
rect 10606 3226 10674 3260
rect 10606 3192 10612 3226
rect 10646 3192 10674 3226
rect 10606 3148 10674 3192
rect 10868 3364 10930 3386
rect 10868 3330 10894 3364
rect 10928 3330 10930 3364
rect 10868 3296 10930 3330
rect 10868 3260 10894 3296
rect 10928 3260 10930 3296
rect 10868 3226 10930 3260
rect 10868 3192 10894 3226
rect 10928 3192 10930 3226
rect 10868 3150 10930 3192
rect 11146 3364 11214 3384
rect 11146 3330 11152 3364
rect 11186 3330 11214 3364
rect 11146 3296 11214 3330
rect 11146 3260 11152 3296
rect 11186 3260 11214 3296
rect 11146 3226 11214 3260
rect 11146 3192 11152 3226
rect 11186 3192 11214 3226
rect 11146 3148 11214 3192
rect 11348 3364 11410 3386
rect 11348 3330 11374 3364
rect 11408 3330 11410 3364
rect 11348 3296 11410 3330
rect 11348 3260 11374 3296
rect 11408 3260 11410 3296
rect 11348 3226 11410 3260
rect 11348 3192 11374 3226
rect 11408 3192 11410 3226
rect 10467 3106 10483 3140
rect 10517 3106 10533 3140
rect 11007 3106 11023 3140
rect 11057 3106 11073 3140
rect 8684 3020 8747 3079
rect 11348 3020 11410 3192
rect 11626 3364 11694 3505
rect 11990 3418 12006 3452
rect 12040 3418 12056 3452
rect 12500 3428 12516 3462
rect 12550 3428 12566 3462
rect 11626 3330 11632 3364
rect 11666 3330 11694 3364
rect 11626 3296 11694 3330
rect 11626 3260 11632 3296
rect 11666 3260 11694 3296
rect 11626 3226 11694 3260
rect 11626 3192 11632 3226
rect 11666 3192 11694 3226
rect 11626 3148 11694 3192
rect 11851 3366 11913 3388
rect 11851 3332 11877 3366
rect 11911 3332 11913 3366
rect 11851 3298 11913 3332
rect 11851 3262 11877 3298
rect 11911 3262 11913 3298
rect 11851 3228 11913 3262
rect 11851 3194 11877 3228
rect 11911 3194 11913 3228
rect 11851 3152 11913 3194
rect 12129 3366 12197 3386
rect 12129 3332 12135 3366
rect 12169 3332 12197 3366
rect 12129 3298 12197 3332
rect 12129 3262 12135 3298
rect 12169 3262 12197 3298
rect 12129 3228 12197 3262
rect 12129 3194 12135 3228
rect 12169 3194 12197 3228
rect 12129 3150 12197 3194
rect 12361 3376 12423 3398
rect 12361 3342 12387 3376
rect 12421 3342 12423 3376
rect 12361 3308 12423 3342
rect 12361 3272 12387 3308
rect 12421 3272 12423 3308
rect 12361 3238 12423 3272
rect 12361 3204 12387 3238
rect 12421 3204 12423 3238
rect 12361 3162 12423 3204
rect 12639 3376 12707 3396
rect 12639 3342 12645 3376
rect 12679 3342 12707 3376
rect 12639 3308 12707 3342
rect 12639 3272 12645 3308
rect 12679 3272 12707 3308
rect 12639 3238 12707 3272
rect 12639 3204 12645 3238
rect 12679 3204 12707 3238
rect 12639 3160 12707 3204
rect 11487 3106 11500 3140
rect 11538 3106 11553 3140
rect 11990 3108 12006 3142
rect 12040 3108 12056 3142
rect 12500 3118 12516 3152
rect 12550 3118 12566 3152
rect 4833 3012 12841 3020
rect 4833 2906 5998 3012
rect 6104 2906 8662 3012
rect 8768 2906 11324 3012
rect 11430 2906 12841 3012
rect 4833 2900 12841 2906
rect 4512 2799 12841 2800
rect 13015 2799 13165 6684
rect 4512 2680 13165 2799
rect 4512 2374 4662 2680
rect 4512 2040 4664 2374
rect 4512 -2978 4662 2040
rect 5340 1930 5612 1960
rect 5340 1892 5436 1930
rect 5502 1892 5612 1930
rect 5340 1806 5612 1892
rect 5340 1804 5544 1806
rect 5340 1768 5358 1804
rect 5396 1770 5544 1804
rect 5582 1770 5612 1806
rect 5396 1768 5612 1770
rect 5340 1732 5612 1768
rect 5692 1888 5756 2680
rect 6726 1929 6998 1959
rect 6064 1889 6080 1923
rect 6234 1889 6250 1923
rect 6726 1891 6822 1929
rect 6888 1891 6998 1929
rect 5692 1804 5748 1888
rect 6572 1857 6636 1858
rect 5692 1770 5711 1804
rect 5745 1770 5748 1804
rect 5692 1732 5748 1770
rect 6567 1804 6636 1857
rect 6567 1770 6569 1804
rect 6603 1770 6636 1804
rect 6567 1738 6636 1770
rect 6064 1651 6080 1685
rect 6234 1651 6250 1685
rect 6564 1204 6636 1738
rect 6726 1805 6998 1891
rect 6726 1803 6930 1805
rect 6726 1767 6744 1803
rect 6782 1769 6930 1803
rect 6968 1769 6998 1805
rect 6782 1767 6998 1769
rect 6726 1731 6998 1767
rect 7096 1929 7368 1959
rect 7096 1891 7192 1929
rect 7258 1891 7368 1929
rect 7096 1805 7368 1891
rect 7096 1803 7300 1805
rect 7096 1767 7114 1803
rect 7152 1769 7300 1803
rect 7338 1769 7368 1805
rect 7152 1767 7368 1769
rect 7096 1731 7368 1767
rect 7518 1929 7790 1959
rect 7518 1891 7614 1929
rect 7680 1891 7790 1929
rect 7518 1805 7790 1891
rect 7518 1803 7722 1805
rect 7518 1767 7536 1803
rect 7574 1769 7722 1803
rect 7760 1769 7790 1805
rect 7574 1767 7790 1769
rect 7518 1731 7790 1767
rect 7940 1929 8212 1959
rect 7940 1891 8036 1929
rect 8102 1891 8212 1929
rect 7940 1805 8212 1891
rect 7940 1803 8144 1805
rect 7940 1767 7958 1803
rect 7996 1769 8144 1803
rect 8182 1769 8212 1805
rect 7996 1767 8212 1769
rect 7940 1731 8212 1767
rect 8362 1874 8426 2680
rect 9440 1933 9712 1961
rect 8741 1889 8757 1923
rect 8911 1889 8927 1923
rect 9440 1895 9536 1933
rect 9602 1895 9712 1933
rect 8362 1804 8424 1874
rect 8362 1770 8388 1804
rect 8422 1770 8424 1804
rect 8362 1728 8424 1770
rect 9244 1804 9317 1872
rect 9244 1770 9246 1804
rect 9280 1770 9317 1804
rect 9244 1726 9317 1770
rect 9440 1809 9712 1895
rect 9440 1807 9644 1809
rect 9440 1771 9458 1807
rect 9496 1773 9644 1807
rect 9682 1773 9712 1809
rect 9496 1771 9712 1773
rect 9440 1735 9712 1771
rect 9810 1933 10082 1961
rect 9810 1895 9906 1933
rect 9972 1895 10082 1933
rect 9810 1809 10082 1895
rect 9810 1807 10014 1809
rect 9810 1771 9828 1807
rect 9866 1773 10014 1807
rect 10052 1773 10082 1809
rect 9866 1771 10082 1773
rect 9810 1735 10082 1771
rect 10232 1933 10504 1961
rect 10232 1895 10328 1933
rect 10394 1895 10504 1933
rect 10232 1809 10504 1895
rect 10232 1807 10436 1809
rect 10232 1771 10250 1807
rect 10288 1773 10436 1807
rect 10474 1773 10504 1809
rect 10288 1771 10504 1773
rect 10232 1735 10504 1771
rect 10654 1933 10926 1961
rect 10654 1895 10750 1933
rect 10816 1895 10926 1933
rect 10654 1809 10926 1895
rect 11024 1826 11088 2680
rect 12568 2679 13165 2680
rect 13015 2390 13165 2679
rect 13014 2008 13166 2390
rect 12038 1930 12310 1960
rect 11405 1890 11421 1924
rect 11575 1890 11591 1924
rect 12038 1892 12134 1930
rect 12200 1892 12310 1930
rect 10654 1807 10858 1809
rect 10654 1771 10672 1807
rect 10710 1773 10858 1807
rect 10896 1773 10926 1809
rect 10710 1771 10926 1773
rect 10654 1735 10926 1771
rect 11025 1805 11088 1826
rect 11025 1771 11052 1805
rect 11086 1771 11088 1805
rect 11025 1748 11088 1771
rect 11908 1805 11962 1876
rect 11908 1771 11910 1805
rect 11944 1771 11962 1805
rect 8741 1651 8757 1685
rect 8911 1651 8927 1685
rect 4858 1168 7246 1204
rect 4852 1166 7246 1168
rect 4852 1085 4884 1166
rect 4851 1002 4884 1085
rect 5042 1002 7246 1166
rect 9244 1146 9316 1726
rect 11908 1712 11962 1771
rect 12038 1806 12310 1892
rect 12038 1804 12242 1806
rect 12038 1768 12056 1804
rect 12094 1770 12242 1804
rect 12280 1770 12310 1806
rect 12094 1768 12310 1770
rect 12038 1732 12310 1768
rect 12435 1925 12609 1946
rect 11405 1652 11421 1686
rect 11575 1652 11591 1686
rect 11907 1644 11962 1712
rect 12435 1663 12456 1925
rect 12593 1663 12609 1925
rect 12435 1647 12609 1663
rect 9244 1140 9916 1146
rect 11906 1140 11962 1644
rect 4851 994 7246 1002
rect 4852 986 7246 994
rect 4858 984 7246 986
rect 5066 972 7246 984
rect 7556 1116 9916 1140
rect 7556 982 7590 1116
rect 7708 982 9916 1116
rect 5254 858 5270 892
rect 5304 858 5320 892
rect 5512 858 5528 892
rect 5562 858 5578 892
rect 5770 858 5786 892
rect 5820 858 5836 892
rect 6028 858 6044 892
rect 6078 858 6094 892
rect 6286 858 6302 892
rect 6336 858 6352 892
rect 6544 858 6560 892
rect 6594 858 6610 892
rect 6802 858 6818 892
rect 6852 858 6868 892
rect 7060 858 7076 892
rect 7110 858 7126 892
rect 5135 808 5180 826
rect 5135 772 5141 808
rect 5175 772 5180 808
rect 5135 738 5180 772
rect 5135 702 5141 738
rect 5175 702 5180 738
rect 5135 668 5180 702
rect 5135 632 5141 668
rect 5175 632 5180 668
rect 5135 390 5180 632
rect 5393 808 5438 852
rect 5393 772 5399 808
rect 5433 772 5438 808
rect 5393 738 5438 772
rect 5393 702 5399 738
rect 5433 702 5438 738
rect 5393 668 5438 702
rect 5393 632 5399 668
rect 5433 632 5438 668
rect 5254 548 5270 582
rect 5304 548 5320 582
rect 5254 440 5270 474
rect 5304 440 5320 474
rect 5135 354 5141 390
rect 5175 354 5180 390
rect 5135 320 5180 354
rect 5135 284 5141 320
rect 5175 284 5180 320
rect 5135 250 5180 284
rect 5135 214 5141 250
rect 5175 214 5180 250
rect 5135 -28 5180 214
rect 5393 390 5438 632
rect 5650 808 5695 852
rect 5650 772 5657 808
rect 5691 772 5695 808
rect 5650 738 5695 772
rect 5650 702 5657 738
rect 5691 702 5695 738
rect 5650 667 5695 702
rect 5650 631 5657 667
rect 5691 631 5695 667
rect 5512 548 5528 582
rect 5562 548 5578 582
rect 5512 440 5528 474
rect 5562 440 5578 474
rect 5393 354 5399 390
rect 5433 354 5438 390
rect 5393 320 5438 354
rect 5393 284 5399 320
rect 5433 284 5438 320
rect 5393 250 5438 284
rect 5393 214 5399 250
rect 5433 214 5438 250
rect 5254 130 5270 164
rect 5304 130 5320 164
rect 5254 22 5270 56
rect 5304 22 5320 56
rect 5135 -64 5141 -28
rect 5175 -64 5180 -28
rect 5135 -98 5180 -64
rect 5135 -134 5141 -98
rect 5175 -134 5180 -98
rect 5135 -168 5180 -134
rect 5135 -204 5141 -168
rect 5175 -204 5180 -168
rect 5135 -446 5180 -204
rect 5393 -28 5438 214
rect 5650 390 5695 631
rect 5910 808 5955 852
rect 5910 772 5915 808
rect 5949 772 5955 808
rect 5910 738 5955 772
rect 5910 702 5915 738
rect 5949 702 5955 738
rect 5910 668 5955 702
rect 5910 632 5915 668
rect 5949 632 5955 668
rect 5770 548 5786 582
rect 5820 548 5836 582
rect 5770 440 5786 474
rect 5820 440 5836 474
rect 5650 354 5657 390
rect 5691 354 5695 390
rect 5650 320 5695 354
rect 5650 284 5657 320
rect 5691 284 5695 320
rect 5650 249 5695 284
rect 5650 213 5657 249
rect 5691 213 5695 249
rect 5512 130 5528 164
rect 5562 130 5578 164
rect 5512 22 5528 56
rect 5562 22 5578 56
rect 5393 -64 5399 -28
rect 5433 -64 5438 -28
rect 5393 -98 5438 -64
rect 5393 -134 5399 -98
rect 5433 -134 5438 -98
rect 5393 -168 5438 -134
rect 5393 -204 5399 -168
rect 5433 -204 5438 -168
rect 5254 -288 5270 -254
rect 5304 -288 5320 -254
rect 5254 -396 5270 -362
rect 5304 -396 5320 -362
rect 5135 -482 5141 -446
rect 5175 -482 5180 -446
rect 5135 -516 5180 -482
rect 5135 -552 5141 -516
rect 5175 -552 5180 -516
rect 5135 -586 5180 -552
rect 5135 -622 5141 -586
rect 5175 -622 5180 -586
rect 5135 -864 5180 -622
rect 5393 -446 5438 -204
rect 5650 -28 5695 213
rect 5910 390 5955 632
rect 6168 808 6213 852
rect 6168 772 6173 808
rect 6207 772 6213 808
rect 6168 738 6213 772
rect 6168 702 6173 738
rect 6207 702 6213 738
rect 6168 668 6213 702
rect 6168 632 6173 668
rect 6207 632 6213 668
rect 6028 548 6044 582
rect 6078 548 6094 582
rect 6028 440 6044 474
rect 6078 440 6094 474
rect 5910 354 5915 390
rect 5949 354 5955 390
rect 5910 320 5955 354
rect 5910 284 5915 320
rect 5949 284 5955 320
rect 5910 250 5955 284
rect 5910 214 5915 250
rect 5949 214 5955 250
rect 5770 130 5786 164
rect 5820 130 5836 164
rect 5770 22 5786 56
rect 5820 22 5836 56
rect 5650 -64 5657 -28
rect 5691 -64 5695 -28
rect 5650 -98 5695 -64
rect 5650 -134 5657 -98
rect 5691 -134 5695 -98
rect 5650 -169 5695 -134
rect 5650 -205 5657 -169
rect 5691 -205 5695 -169
rect 5512 -288 5528 -254
rect 5562 -288 5578 -254
rect 5512 -396 5528 -362
rect 5562 -396 5578 -362
rect 5393 -482 5399 -446
rect 5433 -482 5438 -446
rect 5393 -516 5438 -482
rect 5393 -552 5399 -516
rect 5433 -552 5438 -516
rect 5393 -586 5438 -552
rect 5393 -622 5399 -586
rect 5433 -622 5438 -586
rect 5254 -706 5270 -672
rect 5304 -706 5320 -672
rect 5254 -814 5270 -780
rect 5304 -814 5320 -780
rect 5135 -900 5141 -864
rect 5175 -900 5180 -864
rect 5135 -934 5180 -900
rect 5135 -970 5141 -934
rect 5175 -970 5180 -934
rect 5135 -1004 5180 -970
rect 5135 -1040 5141 -1004
rect 5175 -1040 5180 -1004
rect 5135 -1282 5180 -1040
rect 5393 -864 5438 -622
rect 5650 -446 5695 -205
rect 5910 -28 5955 214
rect 6168 390 6213 632
rect 6425 808 6470 852
rect 6425 772 6431 808
rect 6465 772 6470 808
rect 6425 738 6470 772
rect 6425 702 6431 738
rect 6465 702 6470 738
rect 6425 668 6470 702
rect 6425 632 6431 668
rect 6465 632 6470 668
rect 6286 548 6302 582
rect 6336 548 6352 582
rect 6286 440 6302 474
rect 6336 440 6352 474
rect 6168 354 6173 390
rect 6207 354 6213 390
rect 6168 320 6213 354
rect 6168 284 6173 320
rect 6207 284 6213 320
rect 6168 250 6213 284
rect 6168 214 6173 250
rect 6207 214 6213 250
rect 6028 130 6044 164
rect 6078 130 6094 164
rect 6028 22 6044 56
rect 6078 22 6094 56
rect 5910 -64 5915 -28
rect 5949 -64 5955 -28
rect 5910 -98 5955 -64
rect 5910 -134 5915 -98
rect 5949 -134 5955 -98
rect 5910 -168 5955 -134
rect 5910 -204 5915 -168
rect 5949 -204 5955 -168
rect 5770 -288 5786 -254
rect 5820 -288 5836 -254
rect 5770 -396 5786 -362
rect 5820 -396 5836 -362
rect 5650 -482 5657 -446
rect 5691 -482 5695 -446
rect 5650 -516 5695 -482
rect 5650 -552 5657 -516
rect 5691 -552 5695 -516
rect 5650 -587 5695 -552
rect 5650 -623 5657 -587
rect 5691 -623 5695 -587
rect 5512 -706 5528 -672
rect 5562 -706 5578 -672
rect 5512 -814 5528 -780
rect 5562 -814 5578 -780
rect 5393 -900 5399 -864
rect 5433 -900 5438 -864
rect 5393 -934 5438 -900
rect 5393 -970 5399 -934
rect 5433 -970 5438 -934
rect 5393 -1004 5438 -970
rect 5393 -1040 5399 -1004
rect 5433 -1040 5438 -1004
rect 5254 -1124 5270 -1090
rect 5304 -1124 5320 -1090
rect 5254 -1232 5270 -1198
rect 5304 -1232 5320 -1198
rect 5135 -1318 5141 -1282
rect 5175 -1318 5180 -1282
rect 5135 -1352 5180 -1318
rect 5135 -1388 5141 -1352
rect 5175 -1388 5180 -1352
rect 5135 -1422 5180 -1388
rect 5135 -1458 5141 -1422
rect 5175 -1458 5180 -1422
rect 5135 -1700 5180 -1458
rect 5393 -1282 5438 -1040
rect 5650 -864 5695 -623
rect 5910 -446 5955 -204
rect 6168 -28 6213 214
rect 6425 390 6470 632
rect 6682 808 6727 852
rect 6682 772 6689 808
rect 6723 772 6727 808
rect 6682 738 6727 772
rect 6682 702 6689 738
rect 6723 702 6727 738
rect 6682 668 6727 702
rect 6682 632 6689 668
rect 6723 632 6727 668
rect 6544 548 6560 582
rect 6594 548 6610 582
rect 6544 440 6560 474
rect 6594 440 6610 474
rect 6425 354 6431 390
rect 6465 354 6470 390
rect 6425 320 6470 354
rect 6425 284 6431 320
rect 6465 284 6470 320
rect 6425 250 6470 284
rect 6425 214 6431 250
rect 6465 214 6470 250
rect 6286 130 6302 164
rect 6336 130 6352 164
rect 6286 22 6302 56
rect 6336 22 6352 56
rect 6168 -64 6173 -28
rect 6207 -64 6213 -28
rect 6168 -98 6213 -64
rect 6168 -134 6173 -98
rect 6207 -134 6213 -98
rect 6168 -168 6213 -134
rect 6168 -204 6173 -168
rect 6207 -204 6213 -168
rect 6028 -288 6044 -254
rect 6078 -288 6094 -254
rect 6028 -396 6044 -362
rect 6078 -396 6094 -362
rect 5910 -482 5915 -446
rect 5949 -482 5955 -446
rect 5910 -516 5955 -482
rect 5910 -552 5915 -516
rect 5949 -552 5955 -516
rect 5910 -586 5955 -552
rect 5910 -622 5915 -586
rect 5949 -622 5955 -586
rect 5770 -706 5786 -672
rect 5820 -706 5836 -672
rect 5770 -814 5786 -780
rect 5820 -814 5836 -780
rect 5650 -900 5657 -864
rect 5691 -900 5695 -864
rect 5650 -934 5695 -900
rect 5650 -970 5657 -934
rect 5691 -970 5695 -934
rect 5650 -1005 5695 -970
rect 5650 -1041 5657 -1005
rect 5691 -1041 5695 -1005
rect 5512 -1124 5528 -1090
rect 5562 -1124 5578 -1090
rect 5512 -1232 5528 -1198
rect 5562 -1232 5578 -1198
rect 5393 -1318 5399 -1282
rect 5433 -1318 5438 -1282
rect 5393 -1352 5438 -1318
rect 5393 -1388 5399 -1352
rect 5433 -1388 5438 -1352
rect 5393 -1422 5438 -1388
rect 5393 -1458 5399 -1422
rect 5433 -1458 5438 -1422
rect 5254 -1542 5270 -1508
rect 5304 -1542 5320 -1508
rect 5254 -1650 5270 -1616
rect 5304 -1650 5320 -1616
rect 5135 -1736 5141 -1700
rect 5175 -1736 5180 -1700
rect 5135 -1770 5180 -1736
rect 5135 -1806 5141 -1770
rect 5175 -1806 5180 -1770
rect 5135 -1840 5180 -1806
rect 5135 -1876 5141 -1840
rect 5175 -1876 5180 -1840
rect 5135 -1900 5180 -1876
rect 5134 -2102 5180 -1900
rect 5393 -1700 5438 -1458
rect 5650 -1282 5695 -1041
rect 5910 -864 5955 -622
rect 6168 -446 6213 -204
rect 6425 -28 6470 214
rect 6682 390 6727 632
rect 6941 808 6986 852
rect 7198 816 7244 972
rect 7556 950 9916 982
rect 10162 1106 12696 1140
rect 10162 982 10196 1106
rect 10308 982 12696 1106
rect 10162 960 12696 982
rect 11906 954 12580 960
rect 7556 948 9914 950
rect 7924 858 7940 892
rect 7974 858 7990 892
rect 8182 858 8198 892
rect 8232 858 8248 892
rect 8440 858 8456 892
rect 8490 858 8506 892
rect 8698 858 8714 892
rect 8748 858 8764 892
rect 8956 858 8972 892
rect 9006 858 9022 892
rect 9214 858 9230 892
rect 9264 858 9280 892
rect 9472 858 9488 892
rect 9522 858 9538 892
rect 9730 858 9746 892
rect 9780 858 9796 892
rect 6941 772 6947 808
rect 6981 772 6986 808
rect 6941 738 6986 772
rect 6941 702 6947 738
rect 6981 702 6986 738
rect 6941 668 6986 702
rect 6941 632 6947 668
rect 6981 632 6986 668
rect 6802 548 6818 582
rect 6852 548 6868 582
rect 6802 440 6818 474
rect 6852 440 6868 474
rect 6682 354 6689 390
rect 6723 354 6727 390
rect 6682 320 6727 354
rect 6682 284 6689 320
rect 6723 284 6727 320
rect 6682 250 6727 284
rect 6682 214 6689 250
rect 6723 214 6727 250
rect 6544 130 6560 164
rect 6594 130 6610 164
rect 6544 22 6560 56
rect 6594 22 6610 56
rect 6425 -64 6431 -28
rect 6465 -64 6470 -28
rect 6425 -98 6470 -64
rect 6425 -134 6431 -98
rect 6465 -134 6470 -98
rect 6425 -168 6470 -134
rect 6425 -204 6431 -168
rect 6465 -204 6470 -168
rect 6286 -288 6302 -254
rect 6336 -288 6352 -254
rect 6286 -396 6302 -362
rect 6336 -396 6352 -362
rect 6168 -482 6173 -446
rect 6207 -482 6213 -446
rect 6168 -516 6213 -482
rect 6168 -552 6173 -516
rect 6207 -552 6213 -516
rect 6168 -586 6213 -552
rect 6168 -622 6173 -586
rect 6207 -622 6213 -586
rect 6028 -706 6044 -672
rect 6078 -706 6094 -672
rect 6028 -814 6044 -780
rect 6078 -814 6094 -780
rect 5910 -900 5915 -864
rect 5949 -900 5955 -864
rect 5910 -934 5955 -900
rect 5910 -970 5915 -934
rect 5949 -970 5955 -934
rect 5910 -1004 5955 -970
rect 5910 -1040 5915 -1004
rect 5949 -1040 5955 -1004
rect 5770 -1124 5786 -1090
rect 5820 -1124 5836 -1090
rect 5770 -1232 5786 -1198
rect 5820 -1232 5836 -1198
rect 5650 -1318 5657 -1282
rect 5691 -1318 5695 -1282
rect 5650 -1352 5695 -1318
rect 5650 -1388 5657 -1352
rect 5691 -1388 5695 -1352
rect 5650 -1423 5695 -1388
rect 5650 -1459 5657 -1423
rect 5691 -1459 5695 -1423
rect 5512 -1542 5528 -1508
rect 5562 -1542 5578 -1508
rect 5512 -1650 5528 -1616
rect 5562 -1650 5578 -1616
rect 5393 -1736 5399 -1700
rect 5433 -1736 5438 -1700
rect 5393 -1770 5438 -1736
rect 5393 -1806 5399 -1770
rect 5433 -1806 5438 -1770
rect 5393 -1840 5438 -1806
rect 5393 -1876 5399 -1840
rect 5433 -1876 5438 -1840
rect 5254 -1960 5270 -1926
rect 5304 -1960 5320 -1926
rect 5393 -1994 5438 -1876
rect 5650 -1700 5695 -1459
rect 5910 -1282 5955 -1040
rect 6168 -864 6213 -622
rect 6425 -446 6470 -204
rect 6682 -28 6727 214
rect 6941 390 6986 632
rect 7199 808 7244 816
rect 7199 772 7205 808
rect 7239 772 7244 808
rect 7199 738 7244 772
rect 7199 702 7205 738
rect 7239 702 7244 738
rect 7199 668 7244 702
rect 7199 632 7205 668
rect 7239 632 7244 668
rect 7060 548 7076 582
rect 7110 548 7126 582
rect 7060 440 7076 474
rect 7110 440 7126 474
rect 6941 354 6947 390
rect 6981 354 6986 390
rect 6941 320 6986 354
rect 6941 284 6947 320
rect 6981 284 6986 320
rect 6941 250 6986 284
rect 6941 214 6947 250
rect 6981 214 6986 250
rect 6802 130 6818 164
rect 6852 130 6868 164
rect 6802 22 6818 56
rect 6852 22 6868 56
rect 6682 -64 6689 -28
rect 6723 -64 6727 -28
rect 6682 -98 6727 -64
rect 6682 -134 6689 -98
rect 6723 -134 6727 -98
rect 6682 -168 6727 -134
rect 6682 -204 6689 -168
rect 6723 -204 6727 -168
rect 6544 -288 6560 -254
rect 6594 -288 6610 -254
rect 6544 -396 6560 -362
rect 6594 -396 6610 -362
rect 6425 -482 6431 -446
rect 6465 -482 6470 -446
rect 6425 -516 6470 -482
rect 6425 -552 6431 -516
rect 6465 -552 6470 -516
rect 6425 -586 6470 -552
rect 6425 -622 6431 -586
rect 6465 -622 6470 -586
rect 6286 -706 6302 -672
rect 6336 -706 6352 -672
rect 6286 -814 6302 -780
rect 6336 -814 6352 -780
rect 6168 -900 6173 -864
rect 6207 -900 6213 -864
rect 6168 -934 6213 -900
rect 6168 -970 6173 -934
rect 6207 -970 6213 -934
rect 6168 -1004 6213 -970
rect 6168 -1040 6173 -1004
rect 6207 -1040 6213 -1004
rect 6028 -1124 6044 -1090
rect 6078 -1124 6094 -1090
rect 6028 -1232 6044 -1198
rect 6078 -1232 6094 -1198
rect 5910 -1318 5915 -1282
rect 5949 -1318 5955 -1282
rect 5910 -1352 5955 -1318
rect 5910 -1388 5915 -1352
rect 5949 -1388 5955 -1352
rect 5910 -1422 5955 -1388
rect 5910 -1458 5915 -1422
rect 5949 -1458 5955 -1422
rect 5770 -1542 5786 -1508
rect 5820 -1542 5836 -1508
rect 5770 -1650 5786 -1616
rect 5820 -1650 5836 -1616
rect 5650 -1736 5657 -1700
rect 5691 -1736 5695 -1700
rect 5650 -1770 5695 -1736
rect 5650 -1806 5657 -1770
rect 5691 -1806 5695 -1770
rect 5650 -1841 5695 -1806
rect 5650 -1877 5657 -1841
rect 5691 -1877 5695 -1841
rect 5512 -1960 5528 -1926
rect 5562 -1960 5578 -1926
rect 5650 -1994 5695 -1877
rect 5910 -1700 5955 -1458
rect 6168 -1282 6213 -1040
rect 6425 -864 6470 -622
rect 6682 -446 6727 -204
rect 6941 -28 6986 214
rect 7199 390 7244 632
rect 7199 354 7205 390
rect 7239 354 7244 390
rect 7199 320 7244 354
rect 7199 284 7205 320
rect 7239 284 7244 320
rect 7199 250 7244 284
rect 7199 214 7205 250
rect 7239 214 7244 250
rect 7060 130 7076 164
rect 7110 130 7126 164
rect 7060 22 7076 56
rect 7110 22 7126 56
rect 6941 -64 6947 -28
rect 6981 -64 6986 -28
rect 6941 -98 6986 -64
rect 6941 -134 6947 -98
rect 6981 -134 6986 -98
rect 6941 -168 6986 -134
rect 6941 -204 6947 -168
rect 6981 -204 6986 -168
rect 6802 -288 6818 -254
rect 6852 -288 6868 -254
rect 6802 -396 6818 -362
rect 6852 -396 6868 -362
rect 6682 -482 6689 -446
rect 6723 -482 6727 -446
rect 6682 -516 6727 -482
rect 6682 -552 6689 -516
rect 6723 -552 6727 -516
rect 6682 -586 6727 -552
rect 6682 -622 6689 -586
rect 6723 -622 6727 -586
rect 6544 -706 6560 -672
rect 6594 -706 6610 -672
rect 6544 -814 6560 -780
rect 6594 -814 6610 -780
rect 6425 -900 6431 -864
rect 6465 -900 6470 -864
rect 6425 -934 6470 -900
rect 6425 -970 6431 -934
rect 6465 -970 6470 -934
rect 6425 -1004 6470 -970
rect 6425 -1040 6431 -1004
rect 6465 -1040 6470 -1004
rect 6286 -1124 6302 -1090
rect 6336 -1124 6352 -1090
rect 6286 -1232 6302 -1198
rect 6336 -1232 6352 -1198
rect 6168 -1318 6173 -1282
rect 6207 -1318 6213 -1282
rect 6168 -1352 6213 -1318
rect 6168 -1388 6173 -1352
rect 6207 -1388 6213 -1352
rect 6168 -1422 6213 -1388
rect 6168 -1458 6173 -1422
rect 6207 -1458 6213 -1422
rect 6028 -1542 6044 -1508
rect 6078 -1542 6094 -1508
rect 6028 -1650 6044 -1616
rect 6078 -1650 6094 -1616
rect 5910 -1736 5915 -1700
rect 5949 -1736 5955 -1700
rect 5910 -1770 5955 -1736
rect 5910 -1806 5915 -1770
rect 5949 -1806 5955 -1770
rect 5910 -1840 5955 -1806
rect 5910 -1876 5915 -1840
rect 5949 -1876 5955 -1840
rect 5770 -1960 5786 -1926
rect 5820 -1960 5836 -1926
rect 5910 -1994 5955 -1876
rect 6168 -1700 6213 -1458
rect 6425 -1282 6470 -1040
rect 6682 -864 6727 -622
rect 6941 -446 6986 -204
rect 7199 -28 7244 214
rect 7199 -64 7205 -28
rect 7239 -64 7244 -28
rect 7199 -98 7244 -64
rect 7199 -134 7205 -98
rect 7239 -134 7244 -98
rect 7199 -168 7244 -134
rect 7199 -204 7205 -168
rect 7239 -204 7244 -168
rect 7060 -288 7076 -254
rect 7110 -288 7126 -254
rect 7060 -396 7076 -362
rect 7110 -396 7126 -362
rect 6941 -482 6947 -446
rect 6981 -482 6986 -446
rect 6941 -516 6986 -482
rect 6941 -552 6947 -516
rect 6981 -552 6986 -516
rect 6941 -586 6986 -552
rect 6941 -622 6947 -586
rect 6981 -622 6986 -586
rect 6802 -706 6818 -672
rect 6852 -706 6868 -672
rect 6802 -814 6818 -780
rect 6852 -814 6868 -780
rect 6682 -900 6689 -864
rect 6723 -900 6727 -864
rect 6682 -934 6727 -900
rect 6682 -970 6689 -934
rect 6723 -970 6727 -934
rect 6682 -1004 6727 -970
rect 6682 -1040 6689 -1004
rect 6723 -1040 6727 -1004
rect 6544 -1124 6560 -1090
rect 6594 -1124 6610 -1090
rect 6544 -1232 6560 -1198
rect 6594 -1232 6610 -1198
rect 6425 -1318 6431 -1282
rect 6465 -1318 6470 -1282
rect 6425 -1352 6470 -1318
rect 6425 -1388 6431 -1352
rect 6465 -1388 6470 -1352
rect 6425 -1422 6470 -1388
rect 6425 -1458 6431 -1422
rect 6465 -1458 6470 -1422
rect 6286 -1542 6302 -1508
rect 6336 -1542 6352 -1508
rect 6286 -1650 6302 -1616
rect 6336 -1650 6352 -1616
rect 6168 -1736 6173 -1700
rect 6207 -1736 6213 -1700
rect 6168 -1770 6213 -1736
rect 6168 -1806 6173 -1770
rect 6207 -1806 6213 -1770
rect 6168 -1840 6213 -1806
rect 6168 -1876 6173 -1840
rect 6207 -1876 6213 -1840
rect 6028 -1960 6044 -1926
rect 6078 -1960 6094 -1926
rect 6168 -1994 6213 -1876
rect 6425 -1700 6470 -1458
rect 6682 -1282 6727 -1040
rect 6941 -864 6986 -622
rect 7199 -446 7244 -204
rect 7199 -482 7205 -446
rect 7239 -482 7244 -446
rect 7199 -516 7244 -482
rect 7199 -552 7205 -516
rect 7239 -552 7244 -516
rect 7199 -586 7244 -552
rect 7199 -622 7205 -586
rect 7239 -622 7244 -586
rect 7060 -706 7076 -672
rect 7110 -706 7126 -672
rect 7060 -814 7076 -780
rect 7110 -814 7126 -780
rect 6941 -900 6947 -864
rect 6981 -900 6986 -864
rect 6941 -934 6986 -900
rect 6941 -970 6947 -934
rect 6981 -970 6986 -934
rect 6941 -1004 6986 -970
rect 6941 -1040 6947 -1004
rect 6981 -1040 6986 -1004
rect 6802 -1124 6818 -1090
rect 6852 -1124 6868 -1090
rect 6802 -1232 6818 -1198
rect 6852 -1232 6868 -1198
rect 6682 -1318 6689 -1282
rect 6723 -1318 6727 -1282
rect 6682 -1352 6727 -1318
rect 6682 -1388 6689 -1352
rect 6723 -1388 6727 -1352
rect 6682 -1422 6727 -1388
rect 6682 -1458 6689 -1422
rect 6723 -1458 6727 -1422
rect 6544 -1542 6560 -1508
rect 6594 -1542 6610 -1508
rect 6544 -1650 6560 -1616
rect 6594 -1650 6610 -1616
rect 6425 -1736 6431 -1700
rect 6465 -1736 6470 -1700
rect 6425 -1770 6470 -1736
rect 6425 -1806 6431 -1770
rect 6465 -1806 6470 -1770
rect 6425 -1840 6470 -1806
rect 6425 -1876 6431 -1840
rect 6465 -1876 6470 -1840
rect 6286 -1960 6302 -1926
rect 6336 -1960 6352 -1926
rect 6425 -1994 6470 -1876
rect 6682 -1700 6727 -1458
rect 6941 -1282 6986 -1040
rect 7199 -864 7244 -622
rect 7199 -900 7205 -864
rect 7239 -900 7244 -864
rect 7199 -934 7244 -900
rect 7199 -970 7205 -934
rect 7239 -970 7244 -934
rect 7199 -1004 7244 -970
rect 7199 -1040 7205 -1004
rect 7239 -1040 7244 -1004
rect 7060 -1124 7076 -1090
rect 7110 -1124 7126 -1090
rect 7060 -1232 7076 -1198
rect 7110 -1232 7126 -1198
rect 6941 -1318 6947 -1282
rect 6981 -1318 6986 -1282
rect 6941 -1352 6986 -1318
rect 6941 -1388 6947 -1352
rect 6981 -1388 6986 -1352
rect 6941 -1422 6986 -1388
rect 6941 -1458 6947 -1422
rect 6981 -1458 6986 -1422
rect 6802 -1542 6818 -1508
rect 6852 -1542 6868 -1508
rect 6802 -1650 6818 -1616
rect 6852 -1650 6868 -1616
rect 6682 -1736 6689 -1700
rect 6723 -1736 6727 -1700
rect 6682 -1770 6727 -1736
rect 6682 -1806 6689 -1770
rect 6723 -1806 6727 -1770
rect 6682 -1840 6727 -1806
rect 6682 -1876 6689 -1840
rect 6723 -1876 6727 -1840
rect 6544 -1960 6560 -1926
rect 6594 -1960 6610 -1926
rect 6682 -1994 6727 -1876
rect 6941 -1700 6986 -1458
rect 7199 -1282 7244 -1040
rect 7199 -1318 7205 -1282
rect 7239 -1318 7244 -1282
rect 7199 -1352 7244 -1318
rect 7199 -1388 7205 -1352
rect 7239 -1388 7244 -1352
rect 7199 -1422 7244 -1388
rect 7199 -1458 7205 -1422
rect 7239 -1458 7244 -1422
rect 7060 -1542 7076 -1508
rect 7110 -1542 7126 -1508
rect 7060 -1650 7076 -1616
rect 7110 -1650 7126 -1616
rect 6941 -1736 6947 -1700
rect 6981 -1736 6986 -1700
rect 6941 -1770 6986 -1736
rect 6941 -1806 6947 -1770
rect 6981 -1806 6986 -1770
rect 6941 -1840 6986 -1806
rect 6941 -1876 6947 -1840
rect 6981 -1876 6986 -1840
rect 6802 -1960 6818 -1926
rect 6852 -1960 6868 -1926
rect 6941 -1994 6986 -1876
rect 7199 -1700 7244 -1458
rect 7199 -1736 7205 -1700
rect 7239 -1736 7244 -1700
rect 7199 -1770 7244 -1736
rect 7199 -1806 7205 -1770
rect 7239 -1806 7244 -1770
rect 7199 -1840 7244 -1806
rect 7199 -1876 7205 -1840
rect 7239 -1876 7244 -1840
rect 7199 -1924 7244 -1876
rect 7805 808 7850 826
rect 7805 772 7811 808
rect 7845 772 7850 808
rect 7805 738 7850 772
rect 7805 702 7811 738
rect 7845 702 7850 738
rect 7805 668 7850 702
rect 7805 632 7811 668
rect 7845 632 7850 668
rect 7805 390 7850 632
rect 8063 808 8108 852
rect 8063 772 8069 808
rect 8103 772 8108 808
rect 8063 738 8108 772
rect 8063 702 8069 738
rect 8103 702 8108 738
rect 8063 668 8108 702
rect 8063 632 8069 668
rect 8103 632 8108 668
rect 7924 548 7940 582
rect 7974 548 7990 582
rect 7924 440 7940 474
rect 7974 440 7990 474
rect 7805 354 7811 390
rect 7845 354 7850 390
rect 7805 320 7850 354
rect 7805 284 7811 320
rect 7845 284 7850 320
rect 7805 250 7850 284
rect 7805 214 7811 250
rect 7845 214 7850 250
rect 7805 -28 7850 214
rect 8063 390 8108 632
rect 8320 808 8365 852
rect 8320 772 8327 808
rect 8361 772 8365 808
rect 8320 738 8365 772
rect 8320 702 8327 738
rect 8361 702 8365 738
rect 8320 667 8365 702
rect 8320 631 8327 667
rect 8361 631 8365 667
rect 8182 548 8198 582
rect 8232 548 8248 582
rect 8182 440 8198 474
rect 8232 440 8248 474
rect 8063 354 8069 390
rect 8103 354 8108 390
rect 8063 320 8108 354
rect 8063 284 8069 320
rect 8103 284 8108 320
rect 8063 250 8108 284
rect 8063 214 8069 250
rect 8103 214 8108 250
rect 7924 130 7940 164
rect 7974 130 7990 164
rect 7924 22 7940 56
rect 7974 22 7990 56
rect 7805 -64 7811 -28
rect 7845 -64 7850 -28
rect 7805 -98 7850 -64
rect 7805 -134 7811 -98
rect 7845 -134 7850 -98
rect 7805 -168 7850 -134
rect 7805 -204 7811 -168
rect 7845 -204 7850 -168
rect 7805 -446 7850 -204
rect 8063 -28 8108 214
rect 8320 390 8365 631
rect 8580 808 8625 852
rect 8580 772 8585 808
rect 8619 772 8625 808
rect 8580 738 8625 772
rect 8580 702 8585 738
rect 8619 702 8625 738
rect 8580 668 8625 702
rect 8580 632 8585 668
rect 8619 632 8625 668
rect 8440 548 8456 582
rect 8490 548 8506 582
rect 8440 440 8456 474
rect 8490 440 8506 474
rect 8320 354 8327 390
rect 8361 354 8365 390
rect 8320 320 8365 354
rect 8320 284 8327 320
rect 8361 284 8365 320
rect 8320 249 8365 284
rect 8320 213 8327 249
rect 8361 213 8365 249
rect 8182 130 8198 164
rect 8232 130 8248 164
rect 8182 22 8198 56
rect 8232 22 8248 56
rect 8063 -64 8069 -28
rect 8103 -64 8108 -28
rect 8063 -98 8108 -64
rect 8063 -134 8069 -98
rect 8103 -134 8108 -98
rect 8063 -168 8108 -134
rect 8063 -204 8069 -168
rect 8103 -204 8108 -168
rect 7924 -288 7940 -254
rect 7974 -288 7990 -254
rect 7924 -396 7940 -362
rect 7974 -396 7990 -362
rect 7805 -482 7811 -446
rect 7845 -482 7850 -446
rect 7805 -516 7850 -482
rect 7805 -552 7811 -516
rect 7845 -552 7850 -516
rect 7805 -586 7850 -552
rect 7805 -622 7811 -586
rect 7845 -622 7850 -586
rect 7805 -864 7850 -622
rect 8063 -446 8108 -204
rect 8320 -28 8365 213
rect 8580 390 8625 632
rect 8838 808 8883 852
rect 8838 772 8843 808
rect 8877 772 8883 808
rect 8838 738 8883 772
rect 8838 702 8843 738
rect 8877 702 8883 738
rect 8838 668 8883 702
rect 8838 632 8843 668
rect 8877 632 8883 668
rect 8698 548 8714 582
rect 8748 548 8764 582
rect 8698 440 8714 474
rect 8748 440 8764 474
rect 8580 354 8585 390
rect 8619 354 8625 390
rect 8580 320 8625 354
rect 8580 284 8585 320
rect 8619 284 8625 320
rect 8580 250 8625 284
rect 8580 214 8585 250
rect 8619 214 8625 250
rect 8440 130 8456 164
rect 8490 130 8506 164
rect 8440 22 8456 56
rect 8490 22 8506 56
rect 8320 -64 8327 -28
rect 8361 -64 8365 -28
rect 8320 -98 8365 -64
rect 8320 -134 8327 -98
rect 8361 -134 8365 -98
rect 8320 -169 8365 -134
rect 8320 -205 8327 -169
rect 8361 -205 8365 -169
rect 8182 -288 8198 -254
rect 8232 -288 8248 -254
rect 8182 -396 8198 -362
rect 8232 -396 8248 -362
rect 8063 -482 8069 -446
rect 8103 -482 8108 -446
rect 8063 -516 8108 -482
rect 8063 -552 8069 -516
rect 8103 -552 8108 -516
rect 8063 -586 8108 -552
rect 8063 -622 8069 -586
rect 8103 -622 8108 -586
rect 7924 -706 7940 -672
rect 7974 -706 7990 -672
rect 7924 -814 7940 -780
rect 7974 -814 7990 -780
rect 7805 -900 7811 -864
rect 7845 -900 7850 -864
rect 7805 -934 7850 -900
rect 7805 -970 7811 -934
rect 7845 -970 7850 -934
rect 7805 -1004 7850 -970
rect 7805 -1040 7811 -1004
rect 7845 -1040 7850 -1004
rect 7805 -1282 7850 -1040
rect 8063 -864 8108 -622
rect 8320 -446 8365 -205
rect 8580 -28 8625 214
rect 8838 390 8883 632
rect 9095 808 9140 852
rect 9095 772 9101 808
rect 9135 772 9140 808
rect 9095 738 9140 772
rect 9095 702 9101 738
rect 9135 702 9140 738
rect 9095 668 9140 702
rect 9095 632 9101 668
rect 9135 632 9140 668
rect 8956 548 8972 582
rect 9006 548 9022 582
rect 8956 440 8972 474
rect 9006 440 9022 474
rect 8838 354 8843 390
rect 8877 354 8883 390
rect 8838 320 8883 354
rect 8838 284 8843 320
rect 8877 284 8883 320
rect 8838 250 8883 284
rect 8838 214 8843 250
rect 8877 214 8883 250
rect 8698 130 8714 164
rect 8748 130 8764 164
rect 8698 22 8714 56
rect 8748 22 8764 56
rect 8580 -64 8585 -28
rect 8619 -64 8625 -28
rect 8580 -98 8625 -64
rect 8580 -134 8585 -98
rect 8619 -134 8625 -98
rect 8580 -168 8625 -134
rect 8580 -204 8585 -168
rect 8619 -204 8625 -168
rect 8440 -288 8456 -254
rect 8490 -288 8506 -254
rect 8440 -396 8456 -362
rect 8490 -396 8506 -362
rect 8320 -482 8327 -446
rect 8361 -482 8365 -446
rect 8320 -516 8365 -482
rect 8320 -552 8327 -516
rect 8361 -552 8365 -516
rect 8320 -587 8365 -552
rect 8320 -623 8327 -587
rect 8361 -623 8365 -587
rect 8182 -706 8198 -672
rect 8232 -706 8248 -672
rect 8182 -814 8198 -780
rect 8232 -814 8248 -780
rect 8063 -900 8069 -864
rect 8103 -900 8108 -864
rect 8063 -934 8108 -900
rect 8063 -970 8069 -934
rect 8103 -970 8108 -934
rect 8063 -1004 8108 -970
rect 8063 -1040 8069 -1004
rect 8103 -1040 8108 -1004
rect 7924 -1124 7940 -1090
rect 7974 -1124 7990 -1090
rect 7924 -1232 7940 -1198
rect 7974 -1232 7990 -1198
rect 7805 -1318 7811 -1282
rect 7845 -1318 7850 -1282
rect 7805 -1352 7850 -1318
rect 7805 -1388 7811 -1352
rect 7845 -1388 7850 -1352
rect 7805 -1422 7850 -1388
rect 7805 -1458 7811 -1422
rect 7845 -1458 7850 -1422
rect 7805 -1700 7850 -1458
rect 8063 -1282 8108 -1040
rect 8320 -864 8365 -623
rect 8580 -446 8625 -204
rect 8838 -28 8883 214
rect 9095 390 9140 632
rect 9352 808 9397 852
rect 9352 772 9359 808
rect 9393 772 9397 808
rect 9352 738 9397 772
rect 9352 702 9359 738
rect 9393 702 9397 738
rect 9352 668 9397 702
rect 9352 632 9359 668
rect 9393 632 9397 668
rect 9214 548 9230 582
rect 9264 548 9280 582
rect 9214 440 9230 474
rect 9264 440 9280 474
rect 9095 354 9101 390
rect 9135 354 9140 390
rect 9095 320 9140 354
rect 9095 284 9101 320
rect 9135 284 9140 320
rect 9095 250 9140 284
rect 9095 214 9101 250
rect 9135 214 9140 250
rect 8956 130 8972 164
rect 9006 130 9022 164
rect 8956 22 8972 56
rect 9006 22 9022 56
rect 8838 -64 8843 -28
rect 8877 -64 8883 -28
rect 8838 -98 8883 -64
rect 8838 -134 8843 -98
rect 8877 -134 8883 -98
rect 8838 -168 8883 -134
rect 8838 -204 8843 -168
rect 8877 -204 8883 -168
rect 8698 -288 8714 -254
rect 8748 -288 8764 -254
rect 8698 -396 8714 -362
rect 8748 -396 8764 -362
rect 8580 -482 8585 -446
rect 8619 -482 8625 -446
rect 8580 -516 8625 -482
rect 8580 -552 8585 -516
rect 8619 -552 8625 -516
rect 8580 -586 8625 -552
rect 8580 -622 8585 -586
rect 8619 -622 8625 -586
rect 8440 -706 8456 -672
rect 8490 -706 8506 -672
rect 8440 -814 8456 -780
rect 8490 -814 8506 -780
rect 8320 -900 8327 -864
rect 8361 -900 8365 -864
rect 8320 -934 8365 -900
rect 8320 -970 8327 -934
rect 8361 -970 8365 -934
rect 8320 -1005 8365 -970
rect 8320 -1041 8327 -1005
rect 8361 -1041 8365 -1005
rect 8182 -1124 8198 -1090
rect 8232 -1124 8248 -1090
rect 8182 -1232 8198 -1198
rect 8232 -1232 8248 -1198
rect 8063 -1318 8069 -1282
rect 8103 -1318 8108 -1282
rect 8063 -1352 8108 -1318
rect 8063 -1388 8069 -1352
rect 8103 -1388 8108 -1352
rect 8063 -1422 8108 -1388
rect 8063 -1458 8069 -1422
rect 8103 -1458 8108 -1422
rect 7924 -1542 7940 -1508
rect 7974 -1542 7990 -1508
rect 7924 -1650 7940 -1616
rect 7974 -1650 7990 -1616
rect 7805 -1736 7811 -1700
rect 7845 -1736 7850 -1700
rect 7805 -1770 7850 -1736
rect 7805 -1806 7811 -1770
rect 7845 -1806 7850 -1770
rect 7805 -1840 7850 -1806
rect 7805 -1876 7811 -1840
rect 7845 -1876 7850 -1840
rect 7060 -1960 7076 -1926
rect 7110 -1960 7126 -1926
rect 7805 -1944 7850 -1876
rect 8063 -1700 8108 -1458
rect 8320 -1282 8365 -1041
rect 8580 -864 8625 -622
rect 8838 -446 8883 -204
rect 9095 -28 9140 214
rect 9352 390 9397 632
rect 9611 808 9656 852
rect 9870 828 9914 948
rect 10587 859 10603 893
rect 10637 859 10653 893
rect 10845 859 10861 893
rect 10895 859 10911 893
rect 11103 859 11119 893
rect 11153 859 11169 893
rect 11361 859 11377 893
rect 11411 859 11427 893
rect 11619 859 11635 893
rect 11669 859 11685 893
rect 11877 859 11893 893
rect 11927 859 11943 893
rect 12135 859 12151 893
rect 12185 859 12201 893
rect 12393 859 12409 893
rect 12443 859 12459 893
rect 9611 772 9617 808
rect 9651 772 9656 808
rect 9611 738 9656 772
rect 9611 702 9617 738
rect 9651 702 9656 738
rect 9611 668 9656 702
rect 9611 632 9617 668
rect 9651 632 9656 668
rect 9472 548 9488 582
rect 9522 548 9538 582
rect 9472 440 9488 474
rect 9522 440 9538 474
rect 9352 354 9359 390
rect 9393 354 9397 390
rect 9352 320 9397 354
rect 9352 284 9359 320
rect 9393 284 9397 320
rect 9352 250 9397 284
rect 9352 214 9359 250
rect 9393 214 9397 250
rect 9214 130 9230 164
rect 9264 130 9280 164
rect 9214 22 9230 56
rect 9264 22 9280 56
rect 9095 -64 9101 -28
rect 9135 -64 9140 -28
rect 9095 -98 9140 -64
rect 9095 -134 9101 -98
rect 9135 -134 9140 -98
rect 9095 -168 9140 -134
rect 9095 -204 9101 -168
rect 9135 -204 9140 -168
rect 8956 -288 8972 -254
rect 9006 -288 9022 -254
rect 8956 -396 8972 -362
rect 9006 -396 9022 -362
rect 8838 -482 8843 -446
rect 8877 -482 8883 -446
rect 8838 -516 8883 -482
rect 8838 -552 8843 -516
rect 8877 -552 8883 -516
rect 8838 -586 8883 -552
rect 8838 -622 8843 -586
rect 8877 -622 8883 -586
rect 8698 -706 8714 -672
rect 8748 -706 8764 -672
rect 8698 -814 8714 -780
rect 8748 -814 8764 -780
rect 8580 -900 8585 -864
rect 8619 -900 8625 -864
rect 8580 -934 8625 -900
rect 8580 -970 8585 -934
rect 8619 -970 8625 -934
rect 8580 -1004 8625 -970
rect 8580 -1040 8585 -1004
rect 8619 -1040 8625 -1004
rect 8440 -1124 8456 -1090
rect 8490 -1124 8506 -1090
rect 8440 -1232 8456 -1198
rect 8490 -1232 8506 -1198
rect 8320 -1318 8327 -1282
rect 8361 -1318 8365 -1282
rect 8320 -1352 8365 -1318
rect 8320 -1388 8327 -1352
rect 8361 -1388 8365 -1352
rect 8320 -1423 8365 -1388
rect 8320 -1459 8327 -1423
rect 8361 -1459 8365 -1423
rect 8182 -1542 8198 -1508
rect 8232 -1542 8248 -1508
rect 8182 -1650 8198 -1616
rect 8232 -1650 8248 -1616
rect 8063 -1736 8069 -1700
rect 8103 -1736 8108 -1700
rect 8063 -1770 8108 -1736
rect 8063 -1806 8069 -1770
rect 8103 -1806 8108 -1770
rect 8063 -1840 8108 -1806
rect 8063 -1876 8069 -1840
rect 8103 -1876 8108 -1840
rect 5134 -2184 6364 -2102
rect 7802 -2126 7850 -1944
rect 7924 -1960 7940 -1926
rect 7974 -1960 7990 -1926
rect 8063 -1994 8108 -1876
rect 8320 -1700 8365 -1459
rect 8580 -1282 8625 -1040
rect 8838 -864 8883 -622
rect 9095 -446 9140 -204
rect 9352 -28 9397 214
rect 9611 390 9656 632
rect 9869 808 9914 828
rect 9869 772 9875 808
rect 9909 772 9914 808
rect 9869 738 9914 772
rect 9869 702 9875 738
rect 9909 702 9914 738
rect 9869 668 9914 702
rect 9869 632 9875 668
rect 9909 632 9914 668
rect 9730 548 9746 582
rect 9780 548 9796 582
rect 9730 440 9746 474
rect 9780 440 9796 474
rect 9611 354 9617 390
rect 9651 354 9656 390
rect 9611 320 9656 354
rect 9611 284 9617 320
rect 9651 284 9656 320
rect 9611 250 9656 284
rect 9611 214 9617 250
rect 9651 214 9656 250
rect 9472 130 9488 164
rect 9522 130 9538 164
rect 9472 22 9488 56
rect 9522 22 9538 56
rect 9352 -64 9359 -28
rect 9393 -64 9397 -28
rect 9352 -98 9397 -64
rect 9352 -134 9359 -98
rect 9393 -134 9397 -98
rect 9352 -168 9397 -134
rect 9352 -204 9359 -168
rect 9393 -204 9397 -168
rect 9214 -288 9230 -254
rect 9264 -288 9280 -254
rect 9214 -396 9230 -362
rect 9264 -396 9280 -362
rect 9095 -482 9101 -446
rect 9135 -482 9140 -446
rect 9095 -516 9140 -482
rect 9095 -552 9101 -516
rect 9135 -552 9140 -516
rect 9095 -586 9140 -552
rect 9095 -622 9101 -586
rect 9135 -622 9140 -586
rect 8956 -706 8972 -672
rect 9006 -706 9022 -672
rect 8956 -814 8972 -780
rect 9006 -814 9022 -780
rect 8838 -900 8843 -864
rect 8877 -900 8883 -864
rect 8838 -934 8883 -900
rect 8838 -970 8843 -934
rect 8877 -970 8883 -934
rect 8838 -1004 8883 -970
rect 8838 -1040 8843 -1004
rect 8877 -1040 8883 -1004
rect 8698 -1124 8714 -1090
rect 8748 -1124 8764 -1090
rect 8698 -1232 8714 -1198
rect 8748 -1232 8764 -1198
rect 8580 -1318 8585 -1282
rect 8619 -1318 8625 -1282
rect 8580 -1352 8625 -1318
rect 8580 -1388 8585 -1352
rect 8619 -1388 8625 -1352
rect 8580 -1422 8625 -1388
rect 8580 -1458 8585 -1422
rect 8619 -1458 8625 -1422
rect 8440 -1542 8456 -1508
rect 8490 -1542 8506 -1508
rect 8440 -1650 8456 -1616
rect 8490 -1650 8506 -1616
rect 8320 -1736 8327 -1700
rect 8361 -1736 8365 -1700
rect 8320 -1770 8365 -1736
rect 8320 -1806 8327 -1770
rect 8361 -1806 8365 -1770
rect 8320 -1841 8365 -1806
rect 8320 -1877 8327 -1841
rect 8361 -1877 8365 -1841
rect 8182 -1960 8198 -1926
rect 8232 -1960 8248 -1926
rect 8320 -1994 8365 -1877
rect 8580 -1700 8625 -1458
rect 8838 -1282 8883 -1040
rect 9095 -864 9140 -622
rect 9352 -446 9397 -204
rect 9611 -28 9656 214
rect 9869 390 9914 632
rect 9869 354 9875 390
rect 9909 354 9914 390
rect 9869 320 9914 354
rect 9869 284 9875 320
rect 9909 284 9914 320
rect 9869 250 9914 284
rect 9869 214 9875 250
rect 9909 214 9914 250
rect 9730 130 9746 164
rect 9780 130 9796 164
rect 9730 22 9746 56
rect 9780 22 9796 56
rect 9611 -64 9617 -28
rect 9651 -64 9656 -28
rect 9611 -98 9656 -64
rect 9611 -134 9617 -98
rect 9651 -134 9656 -98
rect 9611 -168 9656 -134
rect 9611 -204 9617 -168
rect 9651 -204 9656 -168
rect 9472 -288 9488 -254
rect 9522 -288 9538 -254
rect 9472 -396 9488 -362
rect 9522 -396 9538 -362
rect 9352 -482 9359 -446
rect 9393 -482 9397 -446
rect 9352 -516 9397 -482
rect 9352 -552 9359 -516
rect 9393 -552 9397 -516
rect 9352 -586 9397 -552
rect 9352 -622 9359 -586
rect 9393 -622 9397 -586
rect 9214 -706 9230 -672
rect 9264 -706 9280 -672
rect 9214 -814 9230 -780
rect 9264 -814 9280 -780
rect 9095 -900 9101 -864
rect 9135 -900 9140 -864
rect 9095 -934 9140 -900
rect 9095 -970 9101 -934
rect 9135 -970 9140 -934
rect 9095 -1004 9140 -970
rect 9095 -1040 9101 -1004
rect 9135 -1040 9140 -1004
rect 8956 -1124 8972 -1090
rect 9006 -1124 9022 -1090
rect 8956 -1232 8972 -1198
rect 9006 -1232 9022 -1198
rect 8838 -1318 8843 -1282
rect 8877 -1318 8883 -1282
rect 8838 -1352 8883 -1318
rect 8838 -1388 8843 -1352
rect 8877 -1388 8883 -1352
rect 8838 -1422 8883 -1388
rect 8838 -1458 8843 -1422
rect 8877 -1458 8883 -1422
rect 8698 -1542 8714 -1508
rect 8748 -1542 8764 -1508
rect 8698 -1650 8714 -1616
rect 8748 -1650 8764 -1616
rect 8580 -1736 8585 -1700
rect 8619 -1736 8625 -1700
rect 8580 -1770 8625 -1736
rect 8580 -1806 8585 -1770
rect 8619 -1806 8625 -1770
rect 8580 -1840 8625 -1806
rect 8580 -1876 8585 -1840
rect 8619 -1876 8625 -1840
rect 8440 -1960 8456 -1926
rect 8490 -1960 8506 -1926
rect 8580 -1994 8625 -1876
rect 8838 -1700 8883 -1458
rect 9095 -1282 9140 -1040
rect 9352 -864 9397 -622
rect 9611 -446 9656 -204
rect 9869 -28 9914 214
rect 9869 -64 9875 -28
rect 9909 -64 9914 -28
rect 9869 -98 9914 -64
rect 9869 -134 9875 -98
rect 9909 -134 9914 -98
rect 9869 -168 9914 -134
rect 9869 -204 9875 -168
rect 9909 -204 9914 -168
rect 9730 -288 9746 -254
rect 9780 -288 9796 -254
rect 9730 -396 9746 -362
rect 9780 -396 9796 -362
rect 9611 -482 9617 -446
rect 9651 -482 9656 -446
rect 9611 -516 9656 -482
rect 9611 -552 9617 -516
rect 9651 -552 9656 -516
rect 9611 -586 9656 -552
rect 9611 -622 9617 -586
rect 9651 -622 9656 -586
rect 9472 -706 9488 -672
rect 9522 -706 9538 -672
rect 9472 -814 9488 -780
rect 9522 -814 9538 -780
rect 9352 -900 9359 -864
rect 9393 -900 9397 -864
rect 9352 -934 9397 -900
rect 9352 -970 9359 -934
rect 9393 -970 9397 -934
rect 9352 -1004 9397 -970
rect 9352 -1040 9359 -1004
rect 9393 -1040 9397 -1004
rect 9214 -1124 9230 -1090
rect 9264 -1124 9280 -1090
rect 9214 -1232 9230 -1198
rect 9264 -1232 9280 -1198
rect 9095 -1318 9101 -1282
rect 9135 -1318 9140 -1282
rect 9095 -1352 9140 -1318
rect 9095 -1388 9101 -1352
rect 9135 -1388 9140 -1352
rect 9095 -1422 9140 -1388
rect 9095 -1458 9101 -1422
rect 9135 -1458 9140 -1422
rect 8956 -1542 8972 -1508
rect 9006 -1542 9022 -1508
rect 8956 -1650 8972 -1616
rect 9006 -1650 9022 -1616
rect 8838 -1736 8843 -1700
rect 8877 -1736 8883 -1700
rect 8838 -1770 8883 -1736
rect 8838 -1806 8843 -1770
rect 8877 -1806 8883 -1770
rect 8838 -1840 8883 -1806
rect 8838 -1876 8843 -1840
rect 8877 -1876 8883 -1840
rect 8698 -1960 8714 -1926
rect 8748 -1960 8764 -1926
rect 8838 -1994 8883 -1876
rect 9095 -1700 9140 -1458
rect 9352 -1282 9397 -1040
rect 9611 -864 9656 -622
rect 9869 -446 9914 -204
rect 9869 -482 9875 -446
rect 9909 -482 9914 -446
rect 9869 -516 9914 -482
rect 9869 -552 9875 -516
rect 9909 -552 9914 -516
rect 9869 -586 9914 -552
rect 9869 -622 9875 -586
rect 9909 -622 9914 -586
rect 9730 -706 9746 -672
rect 9780 -706 9796 -672
rect 9730 -814 9746 -780
rect 9780 -814 9796 -780
rect 9611 -900 9617 -864
rect 9651 -900 9656 -864
rect 9611 -934 9656 -900
rect 9611 -970 9617 -934
rect 9651 -970 9656 -934
rect 9611 -1004 9656 -970
rect 9611 -1040 9617 -1004
rect 9651 -1040 9656 -1004
rect 9472 -1124 9488 -1090
rect 9522 -1124 9538 -1090
rect 9472 -1232 9488 -1198
rect 9522 -1232 9538 -1198
rect 9352 -1318 9359 -1282
rect 9393 -1318 9397 -1282
rect 9352 -1352 9397 -1318
rect 9352 -1388 9359 -1352
rect 9393 -1388 9397 -1352
rect 9352 -1422 9397 -1388
rect 9352 -1458 9359 -1422
rect 9393 -1458 9397 -1422
rect 9214 -1542 9230 -1508
rect 9264 -1542 9280 -1508
rect 9214 -1650 9230 -1616
rect 9264 -1650 9280 -1616
rect 9095 -1736 9101 -1700
rect 9135 -1736 9140 -1700
rect 9095 -1770 9140 -1736
rect 9095 -1806 9101 -1770
rect 9135 -1806 9140 -1770
rect 9095 -1840 9140 -1806
rect 9095 -1876 9101 -1840
rect 9135 -1876 9140 -1840
rect 8956 -1960 8972 -1926
rect 9006 -1960 9022 -1926
rect 9095 -1994 9140 -1876
rect 9352 -1700 9397 -1458
rect 9611 -1282 9656 -1040
rect 9869 -864 9914 -622
rect 9869 -900 9875 -864
rect 9909 -900 9914 -864
rect 9869 -934 9914 -900
rect 9869 -970 9875 -934
rect 9909 -970 9914 -934
rect 9869 -1004 9914 -970
rect 9869 -1040 9875 -1004
rect 9909 -1040 9914 -1004
rect 9730 -1124 9746 -1090
rect 9780 -1124 9796 -1090
rect 9730 -1232 9746 -1198
rect 9780 -1232 9796 -1198
rect 9611 -1318 9617 -1282
rect 9651 -1318 9656 -1282
rect 9611 -1352 9656 -1318
rect 9611 -1388 9617 -1352
rect 9651 -1388 9656 -1352
rect 9611 -1422 9656 -1388
rect 9611 -1458 9617 -1422
rect 9651 -1458 9656 -1422
rect 9472 -1542 9488 -1508
rect 9522 -1542 9538 -1508
rect 9472 -1650 9488 -1616
rect 9522 -1650 9538 -1616
rect 9352 -1736 9359 -1700
rect 9393 -1736 9397 -1700
rect 9352 -1770 9397 -1736
rect 9352 -1806 9359 -1770
rect 9393 -1806 9397 -1770
rect 9352 -1840 9397 -1806
rect 9352 -1876 9359 -1840
rect 9393 -1876 9397 -1840
rect 9214 -1960 9230 -1926
rect 9264 -1960 9280 -1926
rect 9352 -1994 9397 -1876
rect 9611 -1700 9656 -1458
rect 9869 -1282 9914 -1040
rect 9869 -1318 9875 -1282
rect 9909 -1318 9914 -1282
rect 9869 -1352 9914 -1318
rect 9869 -1388 9875 -1352
rect 9909 -1388 9914 -1352
rect 9869 -1422 9914 -1388
rect 9869 -1458 9875 -1422
rect 9909 -1458 9914 -1422
rect 9730 -1542 9746 -1508
rect 9780 -1542 9796 -1508
rect 9730 -1650 9746 -1616
rect 9780 -1650 9796 -1616
rect 9611 -1736 9617 -1700
rect 9651 -1736 9656 -1700
rect 9611 -1770 9656 -1736
rect 9611 -1806 9617 -1770
rect 9651 -1806 9656 -1770
rect 9611 -1840 9656 -1806
rect 9611 -1876 9617 -1840
rect 9651 -1876 9656 -1840
rect 9472 -1960 9488 -1926
rect 9522 -1960 9538 -1926
rect 9611 -1994 9656 -1876
rect 9869 -1700 9914 -1458
rect 9869 -1736 9875 -1700
rect 9909 -1736 9914 -1700
rect 9869 -1770 9914 -1736
rect 9869 -1806 9875 -1770
rect 9909 -1806 9914 -1770
rect 9869 -1840 9914 -1806
rect 9869 -1876 9875 -1840
rect 9909 -1876 9914 -1840
rect 9869 -1906 9914 -1876
rect 10468 809 10513 826
rect 10468 773 10474 809
rect 10508 773 10513 809
rect 10468 739 10513 773
rect 10468 703 10474 739
rect 10508 703 10513 739
rect 10468 669 10513 703
rect 10468 633 10474 669
rect 10508 633 10513 669
rect 10468 391 10513 633
rect 10726 809 10771 853
rect 10726 773 10732 809
rect 10766 773 10771 809
rect 10726 739 10771 773
rect 10726 703 10732 739
rect 10766 703 10771 739
rect 10726 669 10771 703
rect 10726 633 10732 669
rect 10766 633 10771 669
rect 10587 549 10603 583
rect 10637 549 10653 583
rect 10587 441 10603 475
rect 10637 441 10653 475
rect 10468 355 10474 391
rect 10508 355 10513 391
rect 10468 321 10513 355
rect 10468 285 10474 321
rect 10508 285 10513 321
rect 10468 251 10513 285
rect 10468 215 10474 251
rect 10508 215 10513 251
rect 10468 -27 10513 215
rect 10726 391 10771 633
rect 10983 809 11028 853
rect 10983 773 10990 809
rect 11024 773 11028 809
rect 10983 739 11028 773
rect 10983 703 10990 739
rect 11024 703 11028 739
rect 10983 668 11028 703
rect 10983 632 10990 668
rect 11024 632 11028 668
rect 10845 549 10861 583
rect 10895 549 10911 583
rect 10845 441 10861 475
rect 10895 441 10911 475
rect 10726 355 10732 391
rect 10766 355 10771 391
rect 10726 321 10771 355
rect 10726 285 10732 321
rect 10766 285 10771 321
rect 10726 251 10771 285
rect 10726 215 10732 251
rect 10766 215 10771 251
rect 10587 131 10603 165
rect 10637 131 10653 165
rect 10587 23 10603 57
rect 10637 23 10653 57
rect 10468 -63 10474 -27
rect 10508 -63 10513 -27
rect 10468 -97 10513 -63
rect 10468 -133 10474 -97
rect 10508 -133 10513 -97
rect 10468 -167 10513 -133
rect 10468 -203 10474 -167
rect 10508 -203 10513 -167
rect 10468 -445 10513 -203
rect 10726 -27 10771 215
rect 10983 391 11028 632
rect 11243 809 11288 853
rect 11243 773 11248 809
rect 11282 773 11288 809
rect 11243 739 11288 773
rect 11243 703 11248 739
rect 11282 703 11288 739
rect 11243 669 11288 703
rect 11243 633 11248 669
rect 11282 633 11288 669
rect 11103 549 11119 583
rect 11153 549 11169 583
rect 11103 441 11119 475
rect 11153 441 11169 475
rect 10983 355 10990 391
rect 11024 355 11028 391
rect 10983 321 11028 355
rect 10983 285 10990 321
rect 11024 285 11028 321
rect 10983 250 11028 285
rect 10983 214 10990 250
rect 11024 214 11028 250
rect 10845 131 10861 165
rect 10895 131 10911 165
rect 10845 23 10861 57
rect 10895 23 10911 57
rect 10726 -63 10732 -27
rect 10766 -63 10771 -27
rect 10726 -97 10771 -63
rect 10726 -133 10732 -97
rect 10766 -133 10771 -97
rect 10726 -167 10771 -133
rect 10726 -203 10732 -167
rect 10766 -203 10771 -167
rect 10587 -287 10603 -253
rect 10637 -287 10653 -253
rect 10587 -395 10603 -361
rect 10637 -395 10653 -361
rect 10468 -481 10474 -445
rect 10508 -481 10513 -445
rect 10468 -515 10513 -481
rect 10468 -551 10474 -515
rect 10508 -551 10513 -515
rect 10468 -585 10513 -551
rect 10468 -621 10474 -585
rect 10508 -621 10513 -585
rect 10468 -863 10513 -621
rect 10726 -445 10771 -203
rect 10983 -27 11028 214
rect 11243 391 11288 633
rect 11501 809 11546 853
rect 11501 773 11506 809
rect 11540 773 11546 809
rect 11501 739 11546 773
rect 11501 703 11506 739
rect 11540 703 11546 739
rect 11501 669 11546 703
rect 11501 633 11506 669
rect 11540 633 11546 669
rect 11361 549 11377 583
rect 11411 549 11427 583
rect 11361 441 11377 475
rect 11411 441 11427 475
rect 11243 355 11248 391
rect 11282 355 11288 391
rect 11243 321 11288 355
rect 11243 285 11248 321
rect 11282 285 11288 321
rect 11243 251 11288 285
rect 11243 215 11248 251
rect 11282 215 11288 251
rect 11103 131 11119 165
rect 11153 131 11169 165
rect 11103 23 11119 57
rect 11153 23 11169 57
rect 10983 -63 10990 -27
rect 11024 -63 11028 -27
rect 10983 -97 11028 -63
rect 10983 -133 10990 -97
rect 11024 -133 11028 -97
rect 10983 -168 11028 -133
rect 10983 -204 10990 -168
rect 11024 -204 11028 -168
rect 10845 -287 10861 -253
rect 10895 -287 10911 -253
rect 10845 -395 10861 -361
rect 10895 -395 10911 -361
rect 10726 -481 10732 -445
rect 10766 -481 10771 -445
rect 10726 -515 10771 -481
rect 10726 -551 10732 -515
rect 10766 -551 10771 -515
rect 10726 -585 10771 -551
rect 10726 -621 10732 -585
rect 10766 -621 10771 -585
rect 10587 -705 10603 -671
rect 10637 -705 10653 -671
rect 10587 -813 10603 -779
rect 10637 -813 10653 -779
rect 10468 -899 10474 -863
rect 10508 -899 10513 -863
rect 10468 -933 10513 -899
rect 10468 -969 10474 -933
rect 10508 -969 10513 -933
rect 10468 -1003 10513 -969
rect 10468 -1039 10474 -1003
rect 10508 -1039 10513 -1003
rect 10468 -1281 10513 -1039
rect 10726 -863 10771 -621
rect 10983 -445 11028 -204
rect 11243 -27 11288 215
rect 11501 391 11546 633
rect 11758 809 11803 853
rect 11758 773 11764 809
rect 11798 773 11803 809
rect 11758 739 11803 773
rect 11758 703 11764 739
rect 11798 703 11803 739
rect 11758 669 11803 703
rect 11758 633 11764 669
rect 11798 633 11803 669
rect 11619 549 11635 583
rect 11669 549 11685 583
rect 11619 441 11635 475
rect 11669 441 11685 475
rect 11501 355 11506 391
rect 11540 355 11546 391
rect 11501 321 11546 355
rect 11501 285 11506 321
rect 11540 285 11546 321
rect 11501 251 11546 285
rect 11501 215 11506 251
rect 11540 215 11546 251
rect 11361 131 11377 165
rect 11411 131 11427 165
rect 11361 23 11377 57
rect 11411 23 11427 57
rect 11243 -63 11248 -27
rect 11282 -63 11288 -27
rect 11243 -97 11288 -63
rect 11243 -133 11248 -97
rect 11282 -133 11288 -97
rect 11243 -167 11288 -133
rect 11243 -203 11248 -167
rect 11282 -203 11288 -167
rect 11103 -287 11119 -253
rect 11153 -287 11169 -253
rect 11103 -395 11119 -361
rect 11153 -395 11169 -361
rect 10983 -481 10990 -445
rect 11024 -481 11028 -445
rect 10983 -515 11028 -481
rect 10983 -551 10990 -515
rect 11024 -551 11028 -515
rect 10983 -586 11028 -551
rect 10983 -622 10990 -586
rect 11024 -622 11028 -586
rect 10845 -705 10861 -671
rect 10895 -705 10911 -671
rect 10845 -813 10861 -779
rect 10895 -813 10911 -779
rect 10726 -899 10732 -863
rect 10766 -899 10771 -863
rect 10726 -933 10771 -899
rect 10726 -969 10732 -933
rect 10766 -969 10771 -933
rect 10726 -1003 10771 -969
rect 10726 -1039 10732 -1003
rect 10766 -1039 10771 -1003
rect 10587 -1123 10603 -1089
rect 10637 -1123 10653 -1089
rect 10587 -1231 10603 -1197
rect 10637 -1231 10653 -1197
rect 10468 -1317 10474 -1281
rect 10508 -1317 10513 -1281
rect 10468 -1351 10513 -1317
rect 10468 -1387 10474 -1351
rect 10508 -1387 10513 -1351
rect 10468 -1421 10513 -1387
rect 10468 -1457 10474 -1421
rect 10508 -1457 10513 -1421
rect 10468 -1699 10513 -1457
rect 10726 -1281 10771 -1039
rect 10983 -863 11028 -622
rect 11243 -445 11288 -203
rect 11501 -27 11546 215
rect 11758 391 11803 633
rect 12015 809 12060 853
rect 12015 773 12022 809
rect 12056 773 12060 809
rect 12015 739 12060 773
rect 12015 703 12022 739
rect 12056 703 12060 739
rect 12015 669 12060 703
rect 12015 633 12022 669
rect 12056 633 12060 669
rect 11877 549 11893 583
rect 11927 549 11943 583
rect 11877 441 11893 475
rect 11927 441 11943 475
rect 11758 355 11764 391
rect 11798 355 11803 391
rect 11758 321 11803 355
rect 11758 285 11764 321
rect 11798 285 11803 321
rect 11758 251 11803 285
rect 11758 215 11764 251
rect 11798 215 11803 251
rect 11619 131 11635 165
rect 11669 131 11685 165
rect 11619 23 11635 57
rect 11669 23 11685 57
rect 11501 -63 11506 -27
rect 11540 -63 11546 -27
rect 11501 -97 11546 -63
rect 11501 -133 11506 -97
rect 11540 -133 11546 -97
rect 11501 -167 11546 -133
rect 11501 -203 11506 -167
rect 11540 -203 11546 -167
rect 11361 -287 11377 -253
rect 11411 -287 11427 -253
rect 11361 -395 11377 -361
rect 11411 -395 11427 -361
rect 11243 -481 11248 -445
rect 11282 -481 11288 -445
rect 11243 -515 11288 -481
rect 11243 -551 11248 -515
rect 11282 -551 11288 -515
rect 11243 -585 11288 -551
rect 11243 -621 11248 -585
rect 11282 -621 11288 -585
rect 11103 -705 11119 -671
rect 11153 -705 11169 -671
rect 11103 -813 11119 -779
rect 11153 -813 11169 -779
rect 10983 -899 10990 -863
rect 11024 -899 11028 -863
rect 10983 -933 11028 -899
rect 10983 -969 10990 -933
rect 11024 -969 11028 -933
rect 10983 -1004 11028 -969
rect 10983 -1040 10990 -1004
rect 11024 -1040 11028 -1004
rect 10845 -1123 10861 -1089
rect 10895 -1123 10911 -1089
rect 10845 -1231 10861 -1197
rect 10895 -1231 10911 -1197
rect 10726 -1317 10732 -1281
rect 10766 -1317 10771 -1281
rect 10726 -1351 10771 -1317
rect 10726 -1387 10732 -1351
rect 10766 -1387 10771 -1351
rect 10726 -1421 10771 -1387
rect 10726 -1457 10732 -1421
rect 10766 -1457 10771 -1421
rect 10587 -1541 10603 -1507
rect 10637 -1541 10653 -1507
rect 10587 -1649 10603 -1615
rect 10637 -1649 10653 -1615
rect 10468 -1735 10474 -1699
rect 10508 -1735 10513 -1699
rect 10468 -1769 10513 -1735
rect 10468 -1805 10474 -1769
rect 10508 -1805 10513 -1769
rect 10468 -1839 10513 -1805
rect 10468 -1875 10474 -1839
rect 10508 -1875 10513 -1839
rect 9730 -1960 9746 -1926
rect 9780 -1960 9796 -1926
rect 10468 -2032 10513 -1875
rect 10726 -1699 10771 -1457
rect 10983 -1281 11028 -1040
rect 11243 -863 11288 -621
rect 11501 -445 11546 -203
rect 11758 -27 11803 215
rect 12015 391 12060 633
rect 12274 809 12319 853
rect 12274 773 12280 809
rect 12314 773 12319 809
rect 12274 739 12319 773
rect 12274 703 12280 739
rect 12314 703 12319 739
rect 12274 669 12319 703
rect 12274 633 12280 669
rect 12314 633 12319 669
rect 12135 549 12151 583
rect 12185 549 12201 583
rect 12135 441 12151 475
rect 12185 441 12201 475
rect 12015 355 12022 391
rect 12056 355 12060 391
rect 12015 321 12060 355
rect 12015 285 12022 321
rect 12056 285 12060 321
rect 12015 251 12060 285
rect 12015 215 12022 251
rect 12056 215 12060 251
rect 11877 131 11893 165
rect 11927 131 11943 165
rect 11877 23 11893 57
rect 11927 23 11943 57
rect 11758 -63 11764 -27
rect 11798 -63 11803 -27
rect 11758 -97 11803 -63
rect 11758 -133 11764 -97
rect 11798 -133 11803 -97
rect 11758 -167 11803 -133
rect 11758 -203 11764 -167
rect 11798 -203 11803 -167
rect 11619 -287 11635 -253
rect 11669 -287 11685 -253
rect 11619 -395 11635 -361
rect 11669 -395 11685 -361
rect 11501 -481 11506 -445
rect 11540 -481 11546 -445
rect 11501 -515 11546 -481
rect 11501 -551 11506 -515
rect 11540 -551 11546 -515
rect 11501 -585 11546 -551
rect 11501 -621 11506 -585
rect 11540 -621 11546 -585
rect 11361 -705 11377 -671
rect 11411 -705 11427 -671
rect 11361 -813 11377 -779
rect 11411 -813 11427 -779
rect 11243 -899 11248 -863
rect 11282 -899 11288 -863
rect 11243 -933 11288 -899
rect 11243 -969 11248 -933
rect 11282 -969 11288 -933
rect 11243 -1003 11288 -969
rect 11243 -1039 11248 -1003
rect 11282 -1039 11288 -1003
rect 11103 -1123 11119 -1089
rect 11153 -1123 11169 -1089
rect 11103 -1231 11119 -1197
rect 11153 -1231 11169 -1197
rect 10983 -1317 10990 -1281
rect 11024 -1317 11028 -1281
rect 10983 -1351 11028 -1317
rect 10983 -1387 10990 -1351
rect 11024 -1387 11028 -1351
rect 10983 -1422 11028 -1387
rect 10983 -1458 10990 -1422
rect 11024 -1458 11028 -1422
rect 10845 -1541 10861 -1507
rect 10895 -1541 10911 -1507
rect 10845 -1649 10861 -1615
rect 10895 -1649 10911 -1615
rect 10726 -1735 10732 -1699
rect 10766 -1735 10771 -1699
rect 10726 -1769 10771 -1735
rect 10726 -1805 10732 -1769
rect 10766 -1805 10771 -1769
rect 10726 -1839 10771 -1805
rect 10726 -1875 10732 -1839
rect 10766 -1875 10771 -1839
rect 10587 -1959 10603 -1925
rect 10637 -1959 10653 -1925
rect 10726 -1993 10771 -1875
rect 10983 -1699 11028 -1458
rect 11243 -1281 11288 -1039
rect 11501 -863 11546 -621
rect 11758 -445 11803 -203
rect 12015 -27 12060 215
rect 12274 391 12319 633
rect 12532 824 12578 954
rect 12532 809 12577 824
rect 12532 773 12538 809
rect 12572 773 12577 809
rect 12532 739 12577 773
rect 12532 703 12538 739
rect 12572 703 12577 739
rect 12532 669 12577 703
rect 12532 633 12538 669
rect 12572 633 12577 669
rect 12393 549 12409 583
rect 12443 549 12459 583
rect 12393 441 12409 475
rect 12443 441 12459 475
rect 12274 355 12280 391
rect 12314 355 12319 391
rect 12274 321 12319 355
rect 12274 285 12280 321
rect 12314 285 12319 321
rect 12274 251 12319 285
rect 12274 215 12280 251
rect 12314 215 12319 251
rect 12135 131 12151 165
rect 12185 131 12201 165
rect 12135 23 12151 57
rect 12185 23 12201 57
rect 12015 -63 12022 -27
rect 12056 -63 12060 -27
rect 12015 -97 12060 -63
rect 12015 -133 12022 -97
rect 12056 -133 12060 -97
rect 12015 -167 12060 -133
rect 12015 -203 12022 -167
rect 12056 -203 12060 -167
rect 11877 -287 11893 -253
rect 11927 -287 11943 -253
rect 11877 -395 11893 -361
rect 11927 -395 11943 -361
rect 11758 -481 11764 -445
rect 11798 -481 11803 -445
rect 11758 -515 11803 -481
rect 11758 -551 11764 -515
rect 11798 -551 11803 -515
rect 11758 -585 11803 -551
rect 11758 -621 11764 -585
rect 11798 -621 11803 -585
rect 11619 -705 11635 -671
rect 11669 -705 11685 -671
rect 11619 -813 11635 -779
rect 11669 -813 11685 -779
rect 11501 -899 11506 -863
rect 11540 -899 11546 -863
rect 11501 -933 11546 -899
rect 11501 -969 11506 -933
rect 11540 -969 11546 -933
rect 11501 -1003 11546 -969
rect 11501 -1039 11506 -1003
rect 11540 -1039 11546 -1003
rect 11361 -1123 11377 -1089
rect 11411 -1123 11427 -1089
rect 11361 -1231 11377 -1197
rect 11411 -1231 11427 -1197
rect 11243 -1317 11248 -1281
rect 11282 -1317 11288 -1281
rect 11243 -1351 11288 -1317
rect 11243 -1387 11248 -1351
rect 11282 -1387 11288 -1351
rect 11243 -1421 11288 -1387
rect 11243 -1457 11248 -1421
rect 11282 -1457 11288 -1421
rect 11103 -1541 11119 -1507
rect 11153 -1541 11169 -1507
rect 11103 -1649 11119 -1615
rect 11153 -1649 11169 -1615
rect 10983 -1735 10990 -1699
rect 11024 -1735 11028 -1699
rect 10983 -1769 11028 -1735
rect 10983 -1805 10990 -1769
rect 11024 -1805 11028 -1769
rect 10983 -1840 11028 -1805
rect 10983 -1876 10990 -1840
rect 11024 -1876 11028 -1840
rect 10845 -1959 10861 -1925
rect 10895 -1959 10911 -1925
rect 10983 -1993 11028 -1876
rect 11243 -1699 11288 -1457
rect 11501 -1281 11546 -1039
rect 11758 -863 11803 -621
rect 12015 -445 12060 -203
rect 12274 -27 12319 215
rect 12532 391 12577 633
rect 12532 355 12538 391
rect 12572 355 12577 391
rect 12532 321 12577 355
rect 12532 285 12538 321
rect 12572 285 12577 321
rect 12532 251 12577 285
rect 12532 215 12538 251
rect 12572 215 12577 251
rect 12393 131 12409 165
rect 12443 131 12459 165
rect 12393 23 12409 57
rect 12443 23 12459 57
rect 12274 -63 12280 -27
rect 12314 -63 12319 -27
rect 12274 -97 12319 -63
rect 12274 -133 12280 -97
rect 12314 -133 12319 -97
rect 12274 -167 12319 -133
rect 12274 -203 12280 -167
rect 12314 -203 12319 -167
rect 12135 -287 12151 -253
rect 12185 -287 12201 -253
rect 12135 -395 12151 -361
rect 12185 -395 12201 -361
rect 12015 -481 12022 -445
rect 12056 -481 12060 -445
rect 12015 -515 12060 -481
rect 12015 -551 12022 -515
rect 12056 -551 12060 -515
rect 12015 -585 12060 -551
rect 12015 -621 12022 -585
rect 12056 -621 12060 -585
rect 11877 -705 11893 -671
rect 11927 -705 11943 -671
rect 11877 -813 11893 -779
rect 11927 -813 11943 -779
rect 11758 -899 11764 -863
rect 11798 -899 11803 -863
rect 11758 -933 11803 -899
rect 11758 -969 11764 -933
rect 11798 -969 11803 -933
rect 11758 -1003 11803 -969
rect 11758 -1039 11764 -1003
rect 11798 -1039 11803 -1003
rect 11619 -1123 11635 -1089
rect 11669 -1123 11685 -1089
rect 11619 -1231 11635 -1197
rect 11669 -1231 11685 -1197
rect 11501 -1317 11506 -1281
rect 11540 -1317 11546 -1281
rect 11501 -1351 11546 -1317
rect 11501 -1387 11506 -1351
rect 11540 -1387 11546 -1351
rect 11501 -1421 11546 -1387
rect 11501 -1457 11506 -1421
rect 11540 -1457 11546 -1421
rect 11361 -1541 11377 -1507
rect 11411 -1541 11427 -1507
rect 11361 -1649 11377 -1615
rect 11411 -1649 11427 -1615
rect 11243 -1735 11248 -1699
rect 11282 -1735 11288 -1699
rect 11243 -1769 11288 -1735
rect 11243 -1805 11248 -1769
rect 11282 -1805 11288 -1769
rect 11243 -1839 11288 -1805
rect 11243 -1875 11248 -1839
rect 11282 -1875 11288 -1839
rect 11103 -1959 11119 -1925
rect 11153 -1959 11169 -1925
rect 11243 -1993 11288 -1875
rect 11501 -1699 11546 -1457
rect 11758 -1281 11803 -1039
rect 12015 -863 12060 -621
rect 12274 -445 12319 -203
rect 12532 -27 12577 215
rect 12532 -63 12538 -27
rect 12572 -63 12577 -27
rect 12532 -97 12577 -63
rect 12532 -133 12538 -97
rect 12572 -133 12577 -97
rect 12532 -167 12577 -133
rect 12532 -203 12538 -167
rect 12572 -203 12577 -167
rect 12393 -287 12409 -253
rect 12443 -287 12459 -253
rect 12393 -395 12409 -361
rect 12443 -395 12459 -361
rect 12274 -481 12280 -445
rect 12314 -481 12319 -445
rect 12274 -515 12319 -481
rect 12274 -551 12280 -515
rect 12314 -551 12319 -515
rect 12274 -585 12319 -551
rect 12274 -621 12280 -585
rect 12314 -621 12319 -585
rect 12135 -705 12151 -671
rect 12185 -705 12201 -671
rect 12135 -813 12151 -779
rect 12185 -813 12201 -779
rect 12015 -899 12022 -863
rect 12056 -899 12060 -863
rect 12015 -933 12060 -899
rect 12015 -969 12022 -933
rect 12056 -969 12060 -933
rect 12015 -1003 12060 -969
rect 12015 -1039 12022 -1003
rect 12056 -1039 12060 -1003
rect 11877 -1123 11893 -1089
rect 11927 -1123 11943 -1089
rect 11877 -1231 11893 -1197
rect 11927 -1231 11943 -1197
rect 11758 -1317 11764 -1281
rect 11798 -1317 11803 -1281
rect 11758 -1351 11803 -1317
rect 11758 -1387 11764 -1351
rect 11798 -1387 11803 -1351
rect 11758 -1421 11803 -1387
rect 11758 -1457 11764 -1421
rect 11798 -1457 11803 -1421
rect 11619 -1541 11635 -1507
rect 11669 -1541 11685 -1507
rect 11619 -1649 11635 -1615
rect 11669 -1649 11685 -1615
rect 11501 -1735 11506 -1699
rect 11540 -1735 11546 -1699
rect 11501 -1769 11546 -1735
rect 11501 -1805 11506 -1769
rect 11540 -1805 11546 -1769
rect 11501 -1839 11546 -1805
rect 11501 -1875 11506 -1839
rect 11540 -1875 11546 -1839
rect 11361 -1959 11377 -1925
rect 11411 -1959 11427 -1925
rect 11501 -1993 11546 -1875
rect 11758 -1699 11803 -1457
rect 12015 -1281 12060 -1039
rect 12274 -863 12319 -621
rect 12532 -445 12577 -203
rect 12532 -481 12538 -445
rect 12572 -481 12577 -445
rect 12532 -515 12577 -481
rect 12532 -551 12538 -515
rect 12572 -551 12577 -515
rect 12532 -585 12577 -551
rect 12532 -621 12538 -585
rect 12572 -621 12577 -585
rect 12393 -705 12409 -671
rect 12443 -705 12459 -671
rect 12393 -813 12409 -779
rect 12443 -813 12459 -779
rect 12274 -899 12280 -863
rect 12314 -899 12319 -863
rect 12274 -933 12319 -899
rect 12274 -969 12280 -933
rect 12314 -969 12319 -933
rect 12274 -1003 12319 -969
rect 12274 -1039 12280 -1003
rect 12314 -1039 12319 -1003
rect 12135 -1123 12151 -1089
rect 12185 -1123 12201 -1089
rect 12135 -1231 12151 -1197
rect 12185 -1231 12201 -1197
rect 12015 -1317 12022 -1281
rect 12056 -1317 12060 -1281
rect 12015 -1351 12060 -1317
rect 12015 -1387 12022 -1351
rect 12056 -1387 12060 -1351
rect 12015 -1421 12060 -1387
rect 12015 -1457 12022 -1421
rect 12056 -1457 12060 -1421
rect 11877 -1541 11893 -1507
rect 11927 -1541 11943 -1507
rect 11877 -1649 11893 -1615
rect 11927 -1649 11943 -1615
rect 11758 -1735 11764 -1699
rect 11798 -1735 11803 -1699
rect 11758 -1769 11803 -1735
rect 11758 -1805 11764 -1769
rect 11798 -1805 11803 -1769
rect 11758 -1839 11803 -1805
rect 11758 -1875 11764 -1839
rect 11798 -1875 11803 -1839
rect 11619 -1959 11635 -1925
rect 11669 -1959 11685 -1925
rect 11758 -1993 11803 -1875
rect 12015 -1699 12060 -1457
rect 12274 -1281 12319 -1039
rect 12532 -863 12577 -621
rect 12532 -899 12538 -863
rect 12572 -899 12577 -863
rect 12532 -933 12577 -899
rect 12532 -969 12538 -933
rect 12572 -969 12577 -933
rect 12532 -1003 12577 -969
rect 12532 -1039 12538 -1003
rect 12572 -1039 12577 -1003
rect 12393 -1123 12409 -1089
rect 12443 -1123 12459 -1089
rect 12393 -1231 12409 -1197
rect 12443 -1231 12459 -1197
rect 12274 -1317 12280 -1281
rect 12314 -1317 12319 -1281
rect 12274 -1351 12319 -1317
rect 12274 -1387 12280 -1351
rect 12314 -1387 12319 -1351
rect 12274 -1421 12319 -1387
rect 12274 -1457 12280 -1421
rect 12314 -1457 12319 -1421
rect 12135 -1541 12151 -1507
rect 12185 -1541 12201 -1507
rect 12135 -1649 12151 -1615
rect 12185 -1649 12201 -1615
rect 12015 -1735 12022 -1699
rect 12056 -1735 12060 -1699
rect 12015 -1769 12060 -1735
rect 12015 -1805 12022 -1769
rect 12056 -1805 12060 -1769
rect 12015 -1839 12060 -1805
rect 12015 -1875 12022 -1839
rect 12056 -1875 12060 -1839
rect 11877 -1959 11893 -1925
rect 11927 -1959 11943 -1925
rect 12015 -1993 12060 -1875
rect 12274 -1699 12319 -1457
rect 12532 -1281 12577 -1039
rect 12532 -1317 12538 -1281
rect 12572 -1317 12577 -1281
rect 12532 -1351 12577 -1317
rect 12532 -1387 12538 -1351
rect 12572 -1387 12577 -1351
rect 12532 -1421 12577 -1387
rect 12532 -1457 12538 -1421
rect 12572 -1457 12577 -1421
rect 12393 -1541 12409 -1507
rect 12443 -1541 12459 -1507
rect 12393 -1649 12409 -1615
rect 12443 -1649 12459 -1615
rect 12274 -1735 12280 -1699
rect 12314 -1735 12319 -1699
rect 12274 -1769 12319 -1735
rect 12274 -1805 12280 -1769
rect 12314 -1805 12319 -1769
rect 12274 -1839 12319 -1805
rect 12274 -1875 12280 -1839
rect 12314 -1875 12319 -1839
rect 12135 -1959 12151 -1925
rect 12185 -1959 12201 -1925
rect 12274 -1993 12319 -1875
rect 12532 -1699 12577 -1457
rect 12532 -1735 12538 -1699
rect 12572 -1735 12577 -1699
rect 12532 -1769 12577 -1735
rect 12532 -1805 12538 -1769
rect 12572 -1805 12577 -1769
rect 12532 -1839 12577 -1805
rect 12532 -1875 12538 -1839
rect 12572 -1875 12577 -1839
rect 13015 -1856 13165 2008
rect 12532 -1896 12577 -1875
rect 12393 -1959 12409 -1925
rect 12443 -1959 12459 -1925
rect 10462 -2116 10514 -2032
rect 10462 -2117 11692 -2116
rect 6292 -2244 6362 -2184
rect 7802 -2214 9030 -2126
rect 10462 -2178 11694 -2117
rect 7802 -2222 9031 -2214
rect 5134 -2302 5150 -2268
rect 5184 -2302 5200 -2268
rect 5674 -2302 5690 -2268
rect 5724 -2302 5740 -2268
rect 6154 -2302 6165 -2268
rect 6215 -2302 6220 -2268
rect 4995 -2354 5057 -2332
rect 4995 -2388 5021 -2354
rect 5055 -2388 5057 -2354
rect 4995 -2422 5057 -2388
rect 4995 -2458 5021 -2422
rect 5055 -2458 5057 -2422
rect 4995 -2492 5057 -2458
rect 4995 -2526 5021 -2492
rect 5055 -2526 5057 -2492
rect 4995 -2568 5057 -2526
rect 5273 -2354 5341 -2334
rect 5273 -2388 5279 -2354
rect 5313 -2388 5341 -2354
rect 5273 -2422 5341 -2388
rect 5273 -2458 5279 -2422
rect 5313 -2458 5341 -2422
rect 5273 -2492 5341 -2458
rect 5273 -2526 5279 -2492
rect 5313 -2526 5341 -2492
rect 5273 -2570 5341 -2526
rect 5535 -2354 5597 -2332
rect 5535 -2388 5561 -2354
rect 5595 -2388 5597 -2354
rect 5535 -2422 5597 -2388
rect 5535 -2458 5561 -2422
rect 5595 -2458 5597 -2422
rect 5535 -2492 5597 -2458
rect 5535 -2526 5561 -2492
rect 5595 -2526 5597 -2492
rect 5535 -2568 5597 -2526
rect 5813 -2354 5881 -2334
rect 5813 -2388 5819 -2354
rect 5853 -2388 5881 -2354
rect 5813 -2422 5881 -2388
rect 5813 -2458 5819 -2422
rect 5853 -2458 5881 -2422
rect 5813 -2492 5881 -2458
rect 5813 -2526 5819 -2492
rect 5853 -2526 5881 -2492
rect 5813 -2570 5881 -2526
rect 6015 -2354 6077 -2332
rect 6015 -2388 6041 -2354
rect 6075 -2388 6077 -2354
rect 6015 -2422 6077 -2388
rect 6015 -2458 6041 -2422
rect 6075 -2458 6077 -2422
rect 6015 -2492 6077 -2458
rect 6015 -2526 6041 -2492
rect 6075 -2526 6077 -2492
rect 5134 -2612 5150 -2578
rect 5184 -2612 5200 -2578
rect 5674 -2612 5690 -2578
rect 5724 -2612 5740 -2578
rect 6015 -2697 6077 -2526
rect 6293 -2354 6361 -2244
rect 6657 -2300 6673 -2266
rect 6707 -2300 6723 -2266
rect 7167 -2290 7183 -2256
rect 7217 -2290 7233 -2256
rect 7804 -2302 7820 -2268
rect 7854 -2302 7870 -2268
rect 8344 -2302 8360 -2268
rect 8394 -2302 8410 -2268
rect 8824 -2302 8835 -2268
rect 8885 -2302 8890 -2268
rect 6293 -2388 6299 -2354
rect 6333 -2388 6361 -2354
rect 6293 -2422 6361 -2388
rect 6293 -2458 6299 -2422
rect 6333 -2458 6361 -2422
rect 6293 -2492 6361 -2458
rect 6293 -2526 6299 -2492
rect 6333 -2526 6361 -2492
rect 6293 -2570 6361 -2526
rect 6518 -2352 6580 -2330
rect 6518 -2386 6544 -2352
rect 6578 -2386 6580 -2352
rect 6518 -2420 6580 -2386
rect 6518 -2456 6544 -2420
rect 6578 -2456 6580 -2420
rect 6518 -2490 6580 -2456
rect 6518 -2524 6544 -2490
rect 6578 -2524 6580 -2490
rect 6518 -2566 6580 -2524
rect 6796 -2352 6864 -2332
rect 6796 -2386 6802 -2352
rect 6836 -2386 6864 -2352
rect 6796 -2420 6864 -2386
rect 6796 -2456 6802 -2420
rect 6836 -2456 6864 -2420
rect 6796 -2490 6864 -2456
rect 6796 -2524 6802 -2490
rect 6836 -2524 6864 -2490
rect 6796 -2568 6864 -2524
rect 7028 -2342 7090 -2320
rect 7028 -2376 7054 -2342
rect 7088 -2376 7090 -2342
rect 7028 -2410 7090 -2376
rect 7028 -2446 7054 -2410
rect 7088 -2446 7090 -2410
rect 7028 -2480 7090 -2446
rect 7028 -2514 7054 -2480
rect 7088 -2514 7090 -2480
rect 7028 -2556 7090 -2514
rect 7306 -2342 7374 -2322
rect 7306 -2376 7312 -2342
rect 7346 -2376 7374 -2342
rect 7306 -2410 7374 -2376
rect 7306 -2446 7312 -2410
rect 7346 -2446 7374 -2410
rect 7306 -2480 7374 -2446
rect 7306 -2514 7312 -2480
rect 7346 -2514 7374 -2480
rect 7306 -2558 7374 -2514
rect 7665 -2354 7727 -2332
rect 7665 -2388 7691 -2354
rect 7725 -2388 7727 -2354
rect 7665 -2422 7727 -2388
rect 7665 -2458 7691 -2422
rect 7725 -2458 7727 -2422
rect 7665 -2492 7727 -2458
rect 7665 -2526 7691 -2492
rect 7725 -2526 7727 -2492
rect 6154 -2612 6168 -2578
rect 6208 -2612 6220 -2578
rect 6657 -2610 6673 -2576
rect 6707 -2610 6723 -2576
rect 7167 -2600 7183 -2566
rect 7217 -2600 7233 -2566
rect 7665 -2568 7727 -2526
rect 7943 -2354 8011 -2334
rect 7943 -2388 7949 -2354
rect 7983 -2388 8011 -2354
rect 7943 -2422 8011 -2388
rect 7943 -2458 7949 -2422
rect 7983 -2458 8011 -2422
rect 7943 -2492 8011 -2458
rect 7943 -2526 7949 -2492
rect 7983 -2526 8011 -2492
rect 7943 -2570 8011 -2526
rect 8205 -2354 8267 -2332
rect 8205 -2388 8231 -2354
rect 8265 -2388 8267 -2354
rect 8205 -2422 8267 -2388
rect 8205 -2458 8231 -2422
rect 8265 -2458 8267 -2422
rect 8205 -2492 8267 -2458
rect 8205 -2526 8231 -2492
rect 8265 -2526 8267 -2492
rect 8205 -2568 8267 -2526
rect 8483 -2354 8551 -2334
rect 8483 -2388 8489 -2354
rect 8523 -2388 8551 -2354
rect 8483 -2422 8551 -2388
rect 8483 -2458 8489 -2422
rect 8523 -2458 8551 -2422
rect 8483 -2492 8551 -2458
rect 8483 -2526 8489 -2492
rect 8523 -2526 8551 -2492
rect 8483 -2570 8551 -2526
rect 8685 -2354 8747 -2332
rect 8685 -2388 8711 -2354
rect 8745 -2388 8747 -2354
rect 8685 -2422 8747 -2388
rect 8685 -2458 8711 -2422
rect 8745 -2458 8747 -2422
rect 8685 -2492 8747 -2458
rect 8685 -2526 8711 -2492
rect 8745 -2526 8747 -2492
rect 7804 -2612 7820 -2578
rect 7854 -2612 7870 -2578
rect 8344 -2612 8360 -2578
rect 8394 -2612 8410 -2578
rect 8685 -2638 8747 -2526
rect 8963 -2354 9031 -2222
rect 9327 -2300 9343 -2266
rect 9377 -2300 9393 -2266
rect 9837 -2290 9853 -2256
rect 9887 -2290 9903 -2256
rect 10467 -2301 10483 -2267
rect 10517 -2301 10533 -2267
rect 11007 -2301 11023 -2267
rect 11057 -2301 11073 -2267
rect 11487 -2301 11498 -2267
rect 11548 -2301 11553 -2267
rect 8963 -2388 8969 -2354
rect 9003 -2388 9031 -2354
rect 8963 -2422 9031 -2388
rect 8963 -2458 8969 -2422
rect 9003 -2458 9031 -2422
rect 8963 -2492 9031 -2458
rect 8963 -2526 8969 -2492
rect 9003 -2526 9031 -2492
rect 8963 -2570 9031 -2526
rect 9188 -2352 9250 -2330
rect 9188 -2386 9214 -2352
rect 9248 -2386 9250 -2352
rect 9188 -2420 9250 -2386
rect 9188 -2456 9214 -2420
rect 9248 -2456 9250 -2420
rect 9188 -2490 9250 -2456
rect 9188 -2524 9214 -2490
rect 9248 -2524 9250 -2490
rect 9188 -2566 9250 -2524
rect 9466 -2352 9534 -2332
rect 9466 -2386 9472 -2352
rect 9506 -2386 9534 -2352
rect 9466 -2420 9534 -2386
rect 9466 -2456 9472 -2420
rect 9506 -2456 9534 -2420
rect 9466 -2490 9534 -2456
rect 9466 -2524 9472 -2490
rect 9506 -2524 9534 -2490
rect 9466 -2568 9534 -2524
rect 9698 -2342 9760 -2320
rect 9698 -2376 9724 -2342
rect 9758 -2376 9760 -2342
rect 9698 -2410 9760 -2376
rect 9698 -2446 9724 -2410
rect 9758 -2446 9760 -2410
rect 9698 -2480 9760 -2446
rect 9698 -2514 9724 -2480
rect 9758 -2514 9760 -2480
rect 9698 -2556 9760 -2514
rect 9976 -2342 10044 -2322
rect 9976 -2376 9982 -2342
rect 10016 -2376 10044 -2342
rect 9976 -2410 10044 -2376
rect 9976 -2446 9982 -2410
rect 10016 -2446 10044 -2410
rect 9976 -2480 10044 -2446
rect 9976 -2514 9982 -2480
rect 10016 -2514 10044 -2480
rect 9976 -2558 10044 -2514
rect 10328 -2353 10390 -2331
rect 10328 -2387 10354 -2353
rect 10388 -2387 10390 -2353
rect 10328 -2421 10390 -2387
rect 10328 -2457 10354 -2421
rect 10388 -2457 10390 -2421
rect 10328 -2491 10390 -2457
rect 10328 -2525 10354 -2491
rect 10388 -2525 10390 -2491
rect 8824 -2612 8838 -2578
rect 8878 -2612 8890 -2578
rect 9327 -2610 9343 -2576
rect 9377 -2610 9393 -2576
rect 9837 -2600 9853 -2566
rect 9887 -2600 9903 -2566
rect 10328 -2567 10390 -2525
rect 10606 -2353 10674 -2333
rect 10606 -2387 10612 -2353
rect 10646 -2387 10674 -2353
rect 10606 -2421 10674 -2387
rect 10606 -2457 10612 -2421
rect 10646 -2457 10674 -2421
rect 10606 -2491 10674 -2457
rect 10606 -2525 10612 -2491
rect 10646 -2525 10674 -2491
rect 10606 -2569 10674 -2525
rect 10868 -2353 10930 -2331
rect 10868 -2387 10894 -2353
rect 10928 -2387 10930 -2353
rect 10868 -2421 10930 -2387
rect 10868 -2457 10894 -2421
rect 10928 -2457 10930 -2421
rect 10868 -2491 10930 -2457
rect 10868 -2525 10894 -2491
rect 10928 -2525 10930 -2491
rect 10868 -2567 10930 -2525
rect 11146 -2353 11214 -2333
rect 11146 -2387 11152 -2353
rect 11186 -2387 11214 -2353
rect 11146 -2421 11214 -2387
rect 11146 -2457 11152 -2421
rect 11186 -2457 11214 -2421
rect 11146 -2491 11214 -2457
rect 11146 -2525 11152 -2491
rect 11186 -2525 11214 -2491
rect 11146 -2569 11214 -2525
rect 11348 -2353 11410 -2331
rect 11348 -2387 11374 -2353
rect 11408 -2387 11410 -2353
rect 11348 -2421 11410 -2387
rect 11348 -2457 11374 -2421
rect 11408 -2457 11410 -2421
rect 11348 -2491 11410 -2457
rect 11348 -2525 11374 -2491
rect 11408 -2525 11410 -2491
rect 10467 -2611 10483 -2577
rect 10517 -2611 10533 -2577
rect 11007 -2611 11023 -2577
rect 11057 -2611 11073 -2577
rect 8684 -2697 8747 -2638
rect 11348 -2697 11410 -2525
rect 11626 -2353 11694 -2178
rect 11990 -2299 12006 -2265
rect 12040 -2299 12056 -2265
rect 12500 -2289 12516 -2255
rect 12550 -2289 12566 -2255
rect 11626 -2387 11632 -2353
rect 11666 -2387 11694 -2353
rect 11626 -2421 11694 -2387
rect 11626 -2457 11632 -2421
rect 11666 -2457 11694 -2421
rect 11626 -2491 11694 -2457
rect 11626 -2525 11632 -2491
rect 11666 -2525 11694 -2491
rect 11626 -2569 11694 -2525
rect 11851 -2351 11913 -2329
rect 11851 -2385 11877 -2351
rect 11911 -2385 11913 -2351
rect 11851 -2419 11913 -2385
rect 11851 -2455 11877 -2419
rect 11911 -2455 11913 -2419
rect 11851 -2489 11913 -2455
rect 11851 -2523 11877 -2489
rect 11911 -2523 11913 -2489
rect 11851 -2565 11913 -2523
rect 12129 -2351 12197 -2331
rect 12129 -2385 12135 -2351
rect 12169 -2385 12197 -2351
rect 12129 -2419 12197 -2385
rect 12129 -2455 12135 -2419
rect 12169 -2455 12197 -2419
rect 12129 -2489 12197 -2455
rect 12129 -2523 12135 -2489
rect 12169 -2523 12197 -2489
rect 12129 -2567 12197 -2523
rect 12361 -2341 12423 -2319
rect 12361 -2375 12387 -2341
rect 12421 -2375 12423 -2341
rect 12361 -2409 12423 -2375
rect 12361 -2445 12387 -2409
rect 12421 -2445 12423 -2409
rect 12361 -2479 12423 -2445
rect 12361 -2513 12387 -2479
rect 12421 -2513 12423 -2479
rect 12361 -2555 12423 -2513
rect 12639 -2341 12707 -2321
rect 12639 -2375 12645 -2341
rect 12679 -2375 12707 -2341
rect 12639 -2409 12707 -2375
rect 12639 -2445 12645 -2409
rect 12679 -2445 12707 -2409
rect 12639 -2479 12707 -2445
rect 12639 -2513 12645 -2479
rect 12679 -2513 12707 -2479
rect 12639 -2557 12707 -2513
rect 11487 -2611 11498 -2577
rect 11540 -2611 11553 -2577
rect 11990 -2609 12006 -2575
rect 12040 -2609 12056 -2575
rect 12500 -2599 12516 -2565
rect 12550 -2599 12566 -2565
rect 4851 -2707 12841 -2697
rect 4851 -2813 5992 -2707
rect 6098 -2712 12841 -2707
rect 6098 -2806 8668 -2712
rect 8760 -2806 11334 -2712
rect 11426 -2806 12841 -2712
rect 6098 -2813 12841 -2806
rect 4851 -2817 12841 -2813
rect 8684 -2818 8746 -2817
rect 13014 -2978 13166 -1856
rect 4512 -3102 13166 -2978
rect 4979 -3950 5163 -3931
rect 4979 -4214 4998 -3950
rect 5141 -4214 5163 -3950
rect 5385 -3994 5647 -3964
rect 5692 -3994 5756 -3102
rect 8360 -3958 8424 -3102
rect 5385 -4032 5481 -3994
rect 5547 -4032 5647 -3994
rect 5385 -4118 5647 -4032
rect 5385 -4120 5589 -4118
rect 5385 -4156 5403 -4120
rect 5441 -4154 5589 -4120
rect 5627 -4154 5647 -4118
rect 5441 -4156 5647 -4154
rect 5385 -4192 5647 -4156
rect 5693 -4121 5755 -3994
rect 6726 -3996 6998 -3966
rect 6072 -4036 6088 -4002
rect 6242 -4036 6258 -4002
rect 6726 -4034 6822 -3996
rect 6888 -4034 6998 -3996
rect 5693 -4155 5719 -4121
rect 5753 -4155 5755 -4121
rect 4979 -4247 5163 -4214
rect 5693 -4226 5755 -4155
rect 6577 -4121 6622 -4105
rect 6611 -4155 6622 -4121
rect 6072 -4274 6088 -4240
rect 6242 -4274 6258 -4240
rect 6577 -4362 6622 -4155
rect 6726 -4120 6998 -4034
rect 6726 -4122 6930 -4120
rect 6726 -4158 6744 -4122
rect 6782 -4156 6930 -4122
rect 6968 -4156 6998 -4120
rect 6782 -4158 6998 -4156
rect 6726 -4194 6998 -4158
rect 7096 -3996 7368 -3966
rect 7096 -4034 7192 -3996
rect 7258 -4034 7368 -3996
rect 7096 -4120 7368 -4034
rect 7096 -4122 7300 -4120
rect 7096 -4158 7114 -4122
rect 7152 -4156 7300 -4122
rect 7338 -4156 7368 -4120
rect 7152 -4158 7368 -4156
rect 7096 -4194 7368 -4158
rect 7518 -3996 7790 -3966
rect 7518 -4034 7614 -3996
rect 7680 -4034 7790 -3996
rect 7518 -4120 7790 -4034
rect 7518 -4122 7722 -4120
rect 7518 -4158 7536 -4122
rect 7574 -4156 7722 -4122
rect 7760 -4156 7790 -4120
rect 7574 -4158 7790 -4156
rect 7518 -4194 7790 -4158
rect 7940 -3996 8212 -3966
rect 8360 -3974 8425 -3958
rect 7940 -4034 8036 -3996
rect 8102 -4034 8212 -3996
rect 7940 -4120 8212 -4034
rect 7940 -4122 8144 -4120
rect 7940 -4158 7958 -4122
rect 7996 -4156 8144 -4122
rect 8182 -4156 8212 -4120
rect 7996 -4158 8212 -4156
rect 7940 -4194 8212 -4158
rect 8363 -4121 8425 -3974
rect 9427 -3996 9699 -3966
rect 8742 -4036 8758 -4002
rect 8912 -4036 8928 -4002
rect 9427 -4034 9523 -3996
rect 9589 -4034 9699 -3996
rect 8363 -4155 8389 -4121
rect 8423 -4155 8425 -4121
rect 8363 -4226 8425 -4155
rect 9247 -4121 9292 -4105
rect 9281 -4155 9292 -4121
rect 8742 -4274 8758 -4240
rect 8912 -4274 8928 -4240
rect 9247 -4349 9292 -4155
rect 9427 -4120 9699 -4034
rect 9427 -4122 9631 -4120
rect 9427 -4158 9445 -4122
rect 9483 -4156 9631 -4122
rect 9669 -4156 9699 -4120
rect 9483 -4158 9699 -4156
rect 9427 -4194 9699 -4158
rect 9797 -3996 10069 -3966
rect 9797 -4034 9893 -3996
rect 9959 -4034 10069 -3996
rect 9797 -4120 10069 -4034
rect 9797 -4122 10001 -4120
rect 9797 -4158 9815 -4122
rect 9853 -4156 10001 -4122
rect 10039 -4156 10069 -4120
rect 9853 -4158 10069 -4156
rect 9797 -4194 10069 -4158
rect 10219 -3996 10491 -3966
rect 10219 -4034 10315 -3996
rect 10381 -4034 10491 -3996
rect 10219 -4120 10491 -4034
rect 10219 -4122 10423 -4120
rect 10219 -4158 10237 -4122
rect 10275 -4156 10423 -4122
rect 10461 -4156 10491 -4120
rect 10275 -4158 10491 -4156
rect 10219 -4194 10491 -4158
rect 10641 -3996 10913 -3966
rect 10641 -4034 10737 -3996
rect 10803 -4034 10913 -3996
rect 10641 -4120 10913 -4034
rect 10641 -4122 10845 -4120
rect 10641 -4158 10659 -4122
rect 10697 -4156 10845 -4122
rect 10883 -4156 10913 -4120
rect 10697 -4158 10913 -4156
rect 10641 -4194 10913 -4158
rect 11026 -4006 11090 -3102
rect 12261 -3404 12495 -3390
rect 12710 -3402 12726 -3368
rect 12760 -3402 12776 -3368
rect 13100 -3404 13116 -3370
rect 13150 -3404 13166 -3370
rect 12261 -3719 12275 -3404
rect 12477 -3406 12495 -3404
rect 12478 -3557 12495 -3406
rect 12682 -3461 12716 -3445
rect 12478 -3558 12540 -3557
rect 12478 -3576 12682 -3558
rect 12478 -3638 12538 -3576
rect 12594 -3638 12682 -3576
rect 12478 -3652 12682 -3638
rect 12478 -3654 12626 -3652
rect 12478 -3657 12540 -3654
rect 12261 -3720 12276 -3719
rect 12478 -3720 12495 -3657
rect 12261 -3737 12495 -3720
rect 12670 -3773 12682 -3652
rect 12670 -3789 12716 -3773
rect 12770 -3461 12804 -3445
rect 13072 -3463 13106 -3447
rect 12912 -3574 13072 -3560
rect 12912 -3646 12915 -3574
rect 12986 -3646 13072 -3574
rect 12912 -3654 13072 -3646
rect 12804 -3773 12864 -3654
rect 12912 -3656 13016 -3654
rect 12670 -3790 12704 -3789
rect 12770 -3790 12864 -3773
rect 12710 -3866 12726 -3832
rect 12760 -3866 12776 -3832
rect 12820 -3996 12864 -3790
rect 13060 -3775 13072 -3654
rect 13060 -3791 13106 -3775
rect 13160 -3463 13194 -3447
rect 13194 -3775 13254 -3656
rect 13060 -3792 13094 -3791
rect 13160 -3792 13254 -3775
rect 13100 -3868 13116 -3834
rect 13150 -3868 13166 -3834
rect 13210 -3990 13254 -3792
rect 11026 -4120 11088 -4006
rect 11405 -4035 11421 -4001
rect 11575 -4035 11591 -4001
rect 12820 -4008 12950 -3996
rect 12820 -4046 12876 -4008
rect 12930 -4046 12950 -4008
rect 12820 -4054 12950 -4046
rect 13210 -4010 13326 -3990
rect 13210 -4054 13264 -4010
rect 13312 -4054 13326 -4010
rect 11026 -4154 11052 -4120
rect 11086 -4154 11088 -4120
rect 11026 -4225 11088 -4154
rect 11910 -4120 11955 -4104
rect 11944 -4154 11955 -4120
rect 11405 -4273 11421 -4239
rect 11575 -4273 11591 -4239
rect 6577 -4741 6621 -4362
rect 6576 -4803 6621 -4741
rect 9246 -4766 9292 -4349
rect 11910 -4741 11955 -4154
rect 12714 -4198 12730 -4164
rect 12764 -4198 12780 -4164
rect 12538 -4232 12610 -4226
rect 12820 -4232 12864 -4054
rect 13210 -4070 13326 -4054
rect 13104 -4198 13120 -4164
rect 13154 -4198 13170 -4164
rect 12538 -4242 12722 -4232
rect 12538 -4315 12551 -4242
rect 12607 -4248 12722 -4242
rect 12607 -4308 12686 -4248
rect 12720 -4308 12722 -4248
rect 12607 -4315 12722 -4308
rect 12538 -4324 12722 -4315
rect 12774 -4248 12864 -4232
rect 12808 -4308 12864 -4248
rect 12774 -4324 12864 -4308
rect 12928 -4232 13000 -4226
rect 13210 -4232 13254 -4070
rect 12928 -4242 13112 -4232
rect 12928 -4315 12943 -4242
rect 12989 -4248 13112 -4242
rect 12989 -4308 13076 -4248
rect 13110 -4308 13112 -4248
rect 12989 -4315 13112 -4308
rect 12928 -4324 13112 -4315
rect 13164 -4248 13254 -4232
rect 13198 -4308 13254 -4248
rect 13164 -4324 13254 -4308
rect 12538 -4330 12610 -4324
rect 12928 -4330 13000 -4324
rect 12714 -4392 12730 -4358
rect 12764 -4392 12780 -4358
rect 13104 -4392 13120 -4358
rect 13154 -4392 13170 -4358
rect 9246 -4803 9291 -4766
rect 6576 -4814 8917 -4803
rect 6576 -4893 8783 -4814
rect 8878 -4893 8917 -4814
rect 6576 -4908 8917 -4893
rect 6576 -4910 7247 -4908
rect 8654 -4909 8917 -4908
rect 9246 -4814 11575 -4803
rect 11909 -4804 11955 -4741
rect 12524 -4526 12818 -4524
rect 12524 -4568 12870 -4526
rect 12524 -4804 12570 -4568
rect 9246 -4893 11456 -4814
rect 11551 -4893 11575 -4814
rect 9246 -4908 11575 -4893
rect 11906 -4858 12570 -4804
rect 12820 -4858 12870 -4568
rect 11906 -4894 12870 -4858
rect 9246 -4910 9922 -4908
rect 11327 -4909 11575 -4908
rect 11909 -4908 12870 -4894
rect 11909 -4909 12841 -4908
rect 5254 -5046 5270 -5012
rect 5304 -5046 5320 -5012
rect 5512 -5046 5528 -5012
rect 5562 -5046 5578 -5012
rect 5770 -5046 5786 -5012
rect 5820 -5046 5836 -5012
rect 6028 -5046 6044 -5012
rect 6078 -5046 6094 -5012
rect 6286 -5046 6302 -5012
rect 6336 -5046 6352 -5012
rect 6544 -5046 6560 -5012
rect 6594 -5046 6610 -5012
rect 6802 -5046 6818 -5012
rect 6852 -5046 6868 -5012
rect 7060 -5046 7076 -5012
rect 7110 -5046 7126 -5012
rect 5135 -5096 5180 -5052
rect 5135 -5132 5141 -5096
rect 5175 -5132 5180 -5096
rect 5135 -5166 5180 -5132
rect 5135 -5202 5141 -5166
rect 5175 -5202 5180 -5166
rect 5135 -5236 5180 -5202
rect 5135 -5272 5141 -5236
rect 5175 -5272 5180 -5236
rect 5135 -5514 5180 -5272
rect 5393 -5096 5438 -5052
rect 5393 -5132 5399 -5096
rect 5433 -5132 5438 -5096
rect 5393 -5166 5438 -5132
rect 5393 -5202 5399 -5166
rect 5433 -5202 5438 -5166
rect 5393 -5236 5438 -5202
rect 5393 -5272 5399 -5236
rect 5433 -5272 5438 -5236
rect 5254 -5356 5270 -5322
rect 5304 -5356 5320 -5322
rect 5254 -5464 5270 -5430
rect 5304 -5464 5320 -5430
rect 5135 -5550 5141 -5514
rect 5175 -5550 5180 -5514
rect 5135 -5584 5180 -5550
rect 5135 -5620 5141 -5584
rect 5175 -5620 5180 -5584
rect 5135 -5654 5180 -5620
rect 5135 -5690 5141 -5654
rect 5175 -5690 5180 -5654
rect 5135 -5932 5180 -5690
rect 5393 -5514 5438 -5272
rect 5650 -5096 5695 -5052
rect 5650 -5132 5657 -5096
rect 5691 -5132 5695 -5096
rect 5650 -5166 5695 -5132
rect 5650 -5202 5657 -5166
rect 5691 -5202 5695 -5166
rect 5650 -5237 5695 -5202
rect 5650 -5273 5657 -5237
rect 5691 -5273 5695 -5237
rect 5512 -5356 5528 -5322
rect 5562 -5356 5578 -5322
rect 5512 -5464 5528 -5430
rect 5562 -5464 5578 -5430
rect 5393 -5550 5399 -5514
rect 5433 -5550 5438 -5514
rect 5393 -5584 5438 -5550
rect 5393 -5620 5399 -5584
rect 5433 -5620 5438 -5584
rect 5393 -5654 5438 -5620
rect 5393 -5690 5399 -5654
rect 5433 -5690 5438 -5654
rect 5254 -5774 5270 -5740
rect 5304 -5774 5320 -5740
rect 5254 -5882 5270 -5848
rect 5304 -5882 5320 -5848
rect 5135 -5968 5141 -5932
rect 5175 -5968 5180 -5932
rect 5135 -6002 5180 -5968
rect 5135 -6038 5141 -6002
rect 5175 -6038 5180 -6002
rect 5135 -6072 5180 -6038
rect 5135 -6108 5141 -6072
rect 5175 -6108 5180 -6072
rect 5135 -6350 5180 -6108
rect 5393 -5932 5438 -5690
rect 5650 -5514 5695 -5273
rect 5910 -5096 5955 -5052
rect 5910 -5132 5915 -5096
rect 5949 -5132 5955 -5096
rect 5910 -5166 5955 -5132
rect 5910 -5202 5915 -5166
rect 5949 -5202 5955 -5166
rect 5910 -5236 5955 -5202
rect 5910 -5272 5915 -5236
rect 5949 -5272 5955 -5236
rect 5770 -5356 5786 -5322
rect 5820 -5356 5836 -5322
rect 5770 -5464 5786 -5430
rect 5820 -5464 5836 -5430
rect 5650 -5550 5657 -5514
rect 5691 -5550 5695 -5514
rect 5650 -5584 5695 -5550
rect 5650 -5620 5657 -5584
rect 5691 -5620 5695 -5584
rect 5650 -5655 5695 -5620
rect 5650 -5691 5657 -5655
rect 5691 -5691 5695 -5655
rect 5512 -5774 5528 -5740
rect 5562 -5774 5578 -5740
rect 5512 -5882 5528 -5848
rect 5562 -5882 5578 -5848
rect 5393 -5968 5399 -5932
rect 5433 -5968 5438 -5932
rect 5393 -6002 5438 -5968
rect 5393 -6038 5399 -6002
rect 5433 -6038 5438 -6002
rect 5393 -6072 5438 -6038
rect 5393 -6108 5399 -6072
rect 5433 -6108 5438 -6072
rect 5254 -6192 5270 -6158
rect 5304 -6192 5320 -6158
rect 5254 -6300 5270 -6266
rect 5304 -6300 5320 -6266
rect 5135 -6386 5141 -6350
rect 5175 -6386 5180 -6350
rect 5135 -6420 5180 -6386
rect 5135 -6456 5141 -6420
rect 5175 -6456 5180 -6420
rect 5135 -6490 5180 -6456
rect 5135 -6526 5141 -6490
rect 5175 -6526 5180 -6490
rect 5135 -6768 5180 -6526
rect 5393 -6350 5438 -6108
rect 5650 -5932 5695 -5691
rect 5910 -5514 5955 -5272
rect 6168 -5096 6213 -5052
rect 6168 -5132 6173 -5096
rect 6207 -5132 6213 -5096
rect 6168 -5166 6213 -5132
rect 6168 -5202 6173 -5166
rect 6207 -5202 6213 -5166
rect 6168 -5236 6213 -5202
rect 6168 -5272 6173 -5236
rect 6207 -5272 6213 -5236
rect 6028 -5356 6044 -5322
rect 6078 -5356 6094 -5322
rect 6028 -5464 6044 -5430
rect 6078 -5464 6094 -5430
rect 5910 -5550 5915 -5514
rect 5949 -5550 5955 -5514
rect 5910 -5584 5955 -5550
rect 5910 -5620 5915 -5584
rect 5949 -5620 5955 -5584
rect 5910 -5654 5955 -5620
rect 5910 -5690 5915 -5654
rect 5949 -5690 5955 -5654
rect 5770 -5774 5786 -5740
rect 5820 -5774 5836 -5740
rect 5770 -5882 5786 -5848
rect 5820 -5882 5836 -5848
rect 5650 -5968 5657 -5932
rect 5691 -5968 5695 -5932
rect 5650 -6002 5695 -5968
rect 5650 -6038 5657 -6002
rect 5691 -6038 5695 -6002
rect 5650 -6073 5695 -6038
rect 5650 -6109 5657 -6073
rect 5691 -6109 5695 -6073
rect 5512 -6192 5528 -6158
rect 5562 -6192 5578 -6158
rect 5512 -6300 5528 -6266
rect 5562 -6300 5578 -6266
rect 5393 -6386 5399 -6350
rect 5433 -6386 5438 -6350
rect 5393 -6420 5438 -6386
rect 5393 -6456 5399 -6420
rect 5433 -6456 5438 -6420
rect 5393 -6490 5438 -6456
rect 5393 -6526 5399 -6490
rect 5433 -6526 5438 -6490
rect 5254 -6610 5270 -6576
rect 5304 -6610 5320 -6576
rect 5254 -6718 5270 -6684
rect 5304 -6718 5320 -6684
rect 5135 -6804 5141 -6768
rect 5175 -6804 5180 -6768
rect 5135 -6838 5180 -6804
rect 5135 -6874 5141 -6838
rect 5175 -6874 5180 -6838
rect 5135 -6908 5180 -6874
rect 5135 -6944 5141 -6908
rect 5175 -6944 5180 -6908
rect 5135 -7186 5180 -6944
rect 5393 -6768 5438 -6526
rect 5650 -6350 5695 -6109
rect 5910 -5932 5955 -5690
rect 6168 -5514 6213 -5272
rect 6425 -5096 6470 -5052
rect 6425 -5132 6431 -5096
rect 6465 -5132 6470 -5096
rect 6425 -5166 6470 -5132
rect 6425 -5202 6431 -5166
rect 6465 -5202 6470 -5166
rect 6425 -5236 6470 -5202
rect 6425 -5272 6431 -5236
rect 6465 -5272 6470 -5236
rect 6286 -5356 6302 -5322
rect 6336 -5356 6352 -5322
rect 6286 -5464 6302 -5430
rect 6336 -5464 6352 -5430
rect 6168 -5550 6173 -5514
rect 6207 -5550 6213 -5514
rect 6168 -5584 6213 -5550
rect 6168 -5620 6173 -5584
rect 6207 -5620 6213 -5584
rect 6168 -5654 6213 -5620
rect 6168 -5690 6173 -5654
rect 6207 -5690 6213 -5654
rect 6028 -5774 6044 -5740
rect 6078 -5774 6094 -5740
rect 6028 -5882 6044 -5848
rect 6078 -5882 6094 -5848
rect 5910 -5968 5915 -5932
rect 5949 -5968 5955 -5932
rect 5910 -6002 5955 -5968
rect 5910 -6038 5915 -6002
rect 5949 -6038 5955 -6002
rect 5910 -6072 5955 -6038
rect 5910 -6108 5915 -6072
rect 5949 -6108 5955 -6072
rect 5770 -6192 5786 -6158
rect 5820 -6192 5836 -6158
rect 5770 -6300 5786 -6266
rect 5820 -6300 5836 -6266
rect 5650 -6386 5657 -6350
rect 5691 -6386 5695 -6350
rect 5650 -6420 5695 -6386
rect 5650 -6456 5657 -6420
rect 5691 -6456 5695 -6420
rect 5650 -6491 5695 -6456
rect 5650 -6527 5657 -6491
rect 5691 -6527 5695 -6491
rect 5512 -6610 5528 -6576
rect 5562 -6610 5578 -6576
rect 5512 -6718 5528 -6684
rect 5562 -6718 5578 -6684
rect 5393 -6804 5399 -6768
rect 5433 -6804 5438 -6768
rect 5393 -6838 5438 -6804
rect 5393 -6874 5399 -6838
rect 5433 -6874 5438 -6838
rect 5393 -6908 5438 -6874
rect 5393 -6944 5399 -6908
rect 5433 -6944 5438 -6908
rect 5254 -7028 5270 -6994
rect 5304 -7028 5320 -6994
rect 5254 -7136 5270 -7102
rect 5304 -7136 5320 -7102
rect 5135 -7222 5141 -7186
rect 5175 -7222 5180 -7186
rect 5135 -7256 5180 -7222
rect 5135 -7292 5141 -7256
rect 5175 -7292 5180 -7256
rect 5135 -7326 5180 -7292
rect 5135 -7362 5141 -7326
rect 5175 -7362 5180 -7326
rect 5135 -7604 5180 -7362
rect 5393 -7186 5438 -6944
rect 5650 -6768 5695 -6527
rect 5910 -6350 5955 -6108
rect 6168 -5932 6213 -5690
rect 6425 -5514 6470 -5272
rect 6682 -5096 6727 -5052
rect 6682 -5132 6689 -5096
rect 6723 -5132 6727 -5096
rect 6682 -5166 6727 -5132
rect 6682 -5202 6689 -5166
rect 6723 -5202 6727 -5166
rect 6682 -5236 6727 -5202
rect 6682 -5272 6689 -5236
rect 6723 -5272 6727 -5236
rect 6544 -5356 6560 -5322
rect 6594 -5356 6610 -5322
rect 6544 -5464 6560 -5430
rect 6594 -5464 6610 -5430
rect 6425 -5550 6431 -5514
rect 6465 -5550 6470 -5514
rect 6425 -5584 6470 -5550
rect 6425 -5620 6431 -5584
rect 6465 -5620 6470 -5584
rect 6425 -5654 6470 -5620
rect 6425 -5690 6431 -5654
rect 6465 -5690 6470 -5654
rect 6286 -5774 6302 -5740
rect 6336 -5774 6352 -5740
rect 6286 -5882 6302 -5848
rect 6336 -5882 6352 -5848
rect 6168 -5968 6173 -5932
rect 6207 -5968 6213 -5932
rect 6168 -6002 6213 -5968
rect 6168 -6038 6173 -6002
rect 6207 -6038 6213 -6002
rect 6168 -6072 6213 -6038
rect 6168 -6108 6173 -6072
rect 6207 -6108 6213 -6072
rect 6028 -6192 6044 -6158
rect 6078 -6192 6094 -6158
rect 6028 -6300 6044 -6266
rect 6078 -6300 6094 -6266
rect 5910 -6386 5915 -6350
rect 5949 -6386 5955 -6350
rect 5910 -6420 5955 -6386
rect 5910 -6456 5915 -6420
rect 5949 -6456 5955 -6420
rect 5910 -6490 5955 -6456
rect 5910 -6526 5915 -6490
rect 5949 -6526 5955 -6490
rect 5770 -6610 5786 -6576
rect 5820 -6610 5836 -6576
rect 5770 -6718 5786 -6684
rect 5820 -6718 5836 -6684
rect 5650 -6804 5657 -6768
rect 5691 -6804 5695 -6768
rect 5650 -6838 5695 -6804
rect 5650 -6874 5657 -6838
rect 5691 -6874 5695 -6838
rect 5650 -6909 5695 -6874
rect 5650 -6945 5657 -6909
rect 5691 -6945 5695 -6909
rect 5512 -7028 5528 -6994
rect 5562 -7028 5578 -6994
rect 5512 -7136 5528 -7102
rect 5562 -7136 5578 -7102
rect 5393 -7222 5399 -7186
rect 5433 -7222 5438 -7186
rect 5393 -7256 5438 -7222
rect 5393 -7292 5399 -7256
rect 5433 -7292 5438 -7256
rect 5393 -7326 5438 -7292
rect 5393 -7362 5399 -7326
rect 5433 -7362 5438 -7326
rect 5254 -7446 5270 -7412
rect 5304 -7446 5320 -7412
rect 5254 -7554 5270 -7520
rect 5304 -7554 5320 -7520
rect 5135 -7640 5141 -7604
rect 5175 -7640 5180 -7604
rect 5135 -7674 5180 -7640
rect 5135 -7710 5141 -7674
rect 5175 -7710 5180 -7674
rect 5135 -7744 5180 -7710
rect 5135 -7780 5141 -7744
rect 5175 -7780 5180 -7744
rect 5135 -8022 5180 -7780
rect 5393 -7604 5438 -7362
rect 5650 -7186 5695 -6945
rect 5910 -6768 5955 -6526
rect 6168 -6350 6213 -6108
rect 6425 -5932 6470 -5690
rect 6682 -5514 6727 -5272
rect 6941 -5096 6986 -5052
rect 6941 -5132 6947 -5096
rect 6981 -5132 6986 -5096
rect 6941 -5166 6986 -5132
rect 6941 -5202 6947 -5166
rect 6981 -5202 6986 -5166
rect 6941 -5236 6986 -5202
rect 6941 -5272 6947 -5236
rect 6981 -5272 6986 -5236
rect 6802 -5356 6818 -5322
rect 6852 -5356 6868 -5322
rect 6802 -5464 6818 -5430
rect 6852 -5464 6868 -5430
rect 6682 -5550 6689 -5514
rect 6723 -5550 6727 -5514
rect 6682 -5584 6727 -5550
rect 6682 -5620 6689 -5584
rect 6723 -5620 6727 -5584
rect 6682 -5654 6727 -5620
rect 6682 -5690 6689 -5654
rect 6723 -5690 6727 -5654
rect 6544 -5774 6560 -5740
rect 6594 -5774 6610 -5740
rect 6544 -5882 6560 -5848
rect 6594 -5882 6610 -5848
rect 6425 -5968 6431 -5932
rect 6465 -5968 6470 -5932
rect 6425 -6002 6470 -5968
rect 6425 -6038 6431 -6002
rect 6465 -6038 6470 -6002
rect 6425 -6072 6470 -6038
rect 6425 -6108 6431 -6072
rect 6465 -6108 6470 -6072
rect 6286 -6192 6302 -6158
rect 6336 -6192 6352 -6158
rect 6286 -6300 6302 -6266
rect 6336 -6300 6352 -6266
rect 6168 -6386 6173 -6350
rect 6207 -6386 6213 -6350
rect 6168 -6420 6213 -6386
rect 6168 -6456 6173 -6420
rect 6207 -6456 6213 -6420
rect 6168 -6490 6213 -6456
rect 6168 -6526 6173 -6490
rect 6207 -6526 6213 -6490
rect 6028 -6610 6044 -6576
rect 6078 -6610 6094 -6576
rect 6028 -6718 6044 -6684
rect 6078 -6718 6094 -6684
rect 5910 -6804 5915 -6768
rect 5949 -6804 5955 -6768
rect 5910 -6838 5955 -6804
rect 5910 -6874 5915 -6838
rect 5949 -6874 5955 -6838
rect 5910 -6908 5955 -6874
rect 5910 -6944 5915 -6908
rect 5949 -6944 5955 -6908
rect 5770 -7028 5786 -6994
rect 5820 -7028 5836 -6994
rect 5770 -7136 5786 -7102
rect 5820 -7136 5836 -7102
rect 5650 -7222 5657 -7186
rect 5691 -7222 5695 -7186
rect 5650 -7256 5695 -7222
rect 5650 -7292 5657 -7256
rect 5691 -7292 5695 -7256
rect 5650 -7327 5695 -7292
rect 5650 -7363 5657 -7327
rect 5691 -7363 5695 -7327
rect 5512 -7446 5528 -7412
rect 5562 -7446 5578 -7412
rect 5512 -7554 5528 -7520
rect 5562 -7554 5578 -7520
rect 5393 -7640 5399 -7604
rect 5433 -7640 5438 -7604
rect 5393 -7674 5438 -7640
rect 5393 -7710 5399 -7674
rect 5433 -7710 5438 -7674
rect 5393 -7744 5438 -7710
rect 5393 -7780 5399 -7744
rect 5433 -7780 5438 -7744
rect 5254 -7864 5270 -7830
rect 5304 -7864 5320 -7830
rect 5393 -7898 5438 -7780
rect 5650 -7604 5695 -7363
rect 5910 -7186 5955 -6944
rect 6168 -6768 6213 -6526
rect 6425 -6350 6470 -6108
rect 6682 -5932 6727 -5690
rect 6941 -5514 6986 -5272
rect 7199 -5096 7244 -4910
rect 7924 -5046 7940 -5012
rect 7974 -5046 7990 -5012
rect 8182 -5046 8198 -5012
rect 8232 -5046 8248 -5012
rect 8440 -5046 8456 -5012
rect 8490 -5046 8506 -5012
rect 8698 -5046 8714 -5012
rect 8748 -5046 8764 -5012
rect 8956 -5046 8972 -5012
rect 9006 -5046 9022 -5012
rect 9214 -5046 9230 -5012
rect 9264 -5046 9280 -5012
rect 9472 -5046 9488 -5012
rect 9522 -5046 9538 -5012
rect 9730 -5046 9746 -5012
rect 9780 -5046 9796 -5012
rect 7199 -5132 7205 -5096
rect 7239 -5132 7244 -5096
rect 7199 -5166 7244 -5132
rect 7199 -5202 7205 -5166
rect 7239 -5202 7244 -5166
rect 7199 -5236 7244 -5202
rect 7199 -5272 7205 -5236
rect 7239 -5272 7244 -5236
rect 7060 -5356 7076 -5322
rect 7110 -5356 7126 -5322
rect 7060 -5464 7076 -5430
rect 7110 -5464 7126 -5430
rect 6941 -5550 6947 -5514
rect 6981 -5550 6986 -5514
rect 6941 -5584 6986 -5550
rect 6941 -5620 6947 -5584
rect 6981 -5620 6986 -5584
rect 6941 -5654 6986 -5620
rect 6941 -5690 6947 -5654
rect 6981 -5690 6986 -5654
rect 6802 -5774 6818 -5740
rect 6852 -5774 6868 -5740
rect 6802 -5882 6818 -5848
rect 6852 -5882 6868 -5848
rect 6682 -5968 6689 -5932
rect 6723 -5968 6727 -5932
rect 6682 -6002 6727 -5968
rect 6682 -6038 6689 -6002
rect 6723 -6038 6727 -6002
rect 6682 -6072 6727 -6038
rect 6682 -6108 6689 -6072
rect 6723 -6108 6727 -6072
rect 6544 -6192 6560 -6158
rect 6594 -6192 6610 -6158
rect 6544 -6300 6560 -6266
rect 6594 -6300 6610 -6266
rect 6425 -6386 6431 -6350
rect 6465 -6386 6470 -6350
rect 6425 -6420 6470 -6386
rect 6425 -6456 6431 -6420
rect 6465 -6456 6470 -6420
rect 6425 -6490 6470 -6456
rect 6425 -6526 6431 -6490
rect 6465 -6526 6470 -6490
rect 6286 -6610 6302 -6576
rect 6336 -6610 6352 -6576
rect 6286 -6718 6302 -6684
rect 6336 -6718 6352 -6684
rect 6168 -6804 6173 -6768
rect 6207 -6804 6213 -6768
rect 6168 -6838 6213 -6804
rect 6168 -6874 6173 -6838
rect 6207 -6874 6213 -6838
rect 6168 -6908 6213 -6874
rect 6168 -6944 6173 -6908
rect 6207 -6944 6213 -6908
rect 6028 -7028 6044 -6994
rect 6078 -7028 6094 -6994
rect 6028 -7136 6044 -7102
rect 6078 -7136 6094 -7102
rect 5910 -7222 5915 -7186
rect 5949 -7222 5955 -7186
rect 5910 -7256 5955 -7222
rect 5910 -7292 5915 -7256
rect 5949 -7292 5955 -7256
rect 5910 -7326 5955 -7292
rect 5910 -7362 5915 -7326
rect 5949 -7362 5955 -7326
rect 5770 -7446 5786 -7412
rect 5820 -7446 5836 -7412
rect 5770 -7554 5786 -7520
rect 5820 -7554 5836 -7520
rect 5650 -7640 5657 -7604
rect 5691 -7640 5695 -7604
rect 5650 -7674 5695 -7640
rect 5650 -7710 5657 -7674
rect 5691 -7710 5695 -7674
rect 5650 -7745 5695 -7710
rect 5650 -7781 5657 -7745
rect 5691 -7781 5695 -7745
rect 5512 -7864 5528 -7830
rect 5562 -7864 5578 -7830
rect 5650 -7898 5695 -7781
rect 5910 -7604 5955 -7362
rect 6168 -7186 6213 -6944
rect 6425 -6768 6470 -6526
rect 6682 -6350 6727 -6108
rect 6941 -5932 6986 -5690
rect 7199 -5514 7244 -5272
rect 7199 -5550 7205 -5514
rect 7239 -5550 7244 -5514
rect 7199 -5584 7244 -5550
rect 7199 -5620 7205 -5584
rect 7239 -5620 7244 -5584
rect 7199 -5654 7244 -5620
rect 7199 -5690 7205 -5654
rect 7239 -5690 7244 -5654
rect 7060 -5774 7076 -5740
rect 7110 -5774 7126 -5740
rect 7060 -5882 7076 -5848
rect 7110 -5882 7126 -5848
rect 6941 -5968 6947 -5932
rect 6981 -5968 6986 -5932
rect 6941 -6002 6986 -5968
rect 6941 -6038 6947 -6002
rect 6981 -6038 6986 -6002
rect 6941 -6072 6986 -6038
rect 6941 -6108 6947 -6072
rect 6981 -6108 6986 -6072
rect 6802 -6192 6818 -6158
rect 6852 -6192 6868 -6158
rect 6802 -6300 6818 -6266
rect 6852 -6300 6868 -6266
rect 6682 -6386 6689 -6350
rect 6723 -6386 6727 -6350
rect 6682 -6420 6727 -6386
rect 6682 -6456 6689 -6420
rect 6723 -6456 6727 -6420
rect 6682 -6490 6727 -6456
rect 6682 -6526 6689 -6490
rect 6723 -6526 6727 -6490
rect 6544 -6610 6560 -6576
rect 6594 -6610 6610 -6576
rect 6544 -6718 6560 -6684
rect 6594 -6718 6610 -6684
rect 6425 -6804 6431 -6768
rect 6465 -6804 6470 -6768
rect 6425 -6838 6470 -6804
rect 6425 -6874 6431 -6838
rect 6465 -6874 6470 -6838
rect 6425 -6908 6470 -6874
rect 6425 -6944 6431 -6908
rect 6465 -6944 6470 -6908
rect 6286 -7028 6302 -6994
rect 6336 -7028 6352 -6994
rect 6286 -7136 6302 -7102
rect 6336 -7136 6352 -7102
rect 6168 -7222 6173 -7186
rect 6207 -7222 6213 -7186
rect 6168 -7256 6213 -7222
rect 6168 -7292 6173 -7256
rect 6207 -7292 6213 -7256
rect 6168 -7326 6213 -7292
rect 6168 -7362 6173 -7326
rect 6207 -7362 6213 -7326
rect 6028 -7446 6044 -7412
rect 6078 -7446 6094 -7412
rect 6028 -7554 6044 -7520
rect 6078 -7554 6094 -7520
rect 5910 -7640 5915 -7604
rect 5949 -7640 5955 -7604
rect 5910 -7674 5955 -7640
rect 5910 -7710 5915 -7674
rect 5949 -7710 5955 -7674
rect 5910 -7744 5955 -7710
rect 5910 -7780 5915 -7744
rect 5949 -7780 5955 -7744
rect 5770 -7864 5786 -7830
rect 5820 -7864 5836 -7830
rect 5910 -7898 5955 -7780
rect 6168 -7604 6213 -7362
rect 6425 -7186 6470 -6944
rect 6682 -6768 6727 -6526
rect 6941 -6350 6986 -6108
rect 7199 -5932 7244 -5690
rect 7199 -5968 7205 -5932
rect 7239 -5968 7244 -5932
rect 7199 -6002 7244 -5968
rect 7199 -6038 7205 -6002
rect 7239 -6038 7244 -6002
rect 7199 -6072 7244 -6038
rect 7199 -6108 7205 -6072
rect 7239 -6108 7244 -6072
rect 7060 -6192 7076 -6158
rect 7110 -6192 7126 -6158
rect 7060 -6300 7076 -6266
rect 7110 -6300 7126 -6266
rect 6941 -6386 6947 -6350
rect 6981 -6386 6986 -6350
rect 6941 -6420 6986 -6386
rect 6941 -6456 6947 -6420
rect 6981 -6456 6986 -6420
rect 6941 -6490 6986 -6456
rect 6941 -6526 6947 -6490
rect 6981 -6526 6986 -6490
rect 6802 -6610 6818 -6576
rect 6852 -6610 6868 -6576
rect 6802 -6718 6818 -6684
rect 6852 -6718 6868 -6684
rect 6682 -6804 6689 -6768
rect 6723 -6804 6727 -6768
rect 6682 -6838 6727 -6804
rect 6682 -6874 6689 -6838
rect 6723 -6874 6727 -6838
rect 6682 -6908 6727 -6874
rect 6682 -6944 6689 -6908
rect 6723 -6944 6727 -6908
rect 6544 -7028 6560 -6994
rect 6594 -7028 6610 -6994
rect 6544 -7136 6560 -7102
rect 6594 -7136 6610 -7102
rect 6425 -7222 6431 -7186
rect 6465 -7222 6470 -7186
rect 6425 -7256 6470 -7222
rect 6425 -7292 6431 -7256
rect 6465 -7292 6470 -7256
rect 6425 -7326 6470 -7292
rect 6425 -7362 6431 -7326
rect 6465 -7362 6470 -7326
rect 6286 -7446 6302 -7412
rect 6336 -7446 6352 -7412
rect 6286 -7554 6302 -7520
rect 6336 -7554 6352 -7520
rect 6168 -7640 6173 -7604
rect 6207 -7640 6213 -7604
rect 6168 -7674 6213 -7640
rect 6168 -7710 6173 -7674
rect 6207 -7710 6213 -7674
rect 6168 -7744 6213 -7710
rect 6168 -7780 6173 -7744
rect 6207 -7780 6213 -7744
rect 6028 -7864 6044 -7830
rect 6078 -7864 6094 -7830
rect 6168 -7898 6213 -7780
rect 6425 -7604 6470 -7362
rect 6682 -7186 6727 -6944
rect 6941 -6768 6986 -6526
rect 7199 -6350 7244 -6108
rect 7199 -6386 7205 -6350
rect 7239 -6386 7244 -6350
rect 7199 -6420 7244 -6386
rect 7199 -6456 7205 -6420
rect 7239 -6456 7244 -6420
rect 7199 -6490 7244 -6456
rect 7199 -6526 7205 -6490
rect 7239 -6526 7244 -6490
rect 7060 -6610 7076 -6576
rect 7110 -6610 7126 -6576
rect 7060 -6718 7076 -6684
rect 7110 -6718 7126 -6684
rect 6941 -6804 6947 -6768
rect 6981 -6804 6986 -6768
rect 6941 -6838 6986 -6804
rect 6941 -6874 6947 -6838
rect 6981 -6874 6986 -6838
rect 6941 -6908 6986 -6874
rect 6941 -6944 6947 -6908
rect 6981 -6944 6986 -6908
rect 6802 -7028 6818 -6994
rect 6852 -7028 6868 -6994
rect 6802 -7136 6818 -7102
rect 6852 -7136 6868 -7102
rect 6682 -7222 6689 -7186
rect 6723 -7222 6727 -7186
rect 6682 -7256 6727 -7222
rect 6682 -7292 6689 -7256
rect 6723 -7292 6727 -7256
rect 6682 -7326 6727 -7292
rect 6682 -7362 6689 -7326
rect 6723 -7362 6727 -7326
rect 6544 -7446 6560 -7412
rect 6594 -7446 6610 -7412
rect 6544 -7554 6560 -7520
rect 6594 -7554 6610 -7520
rect 6425 -7640 6431 -7604
rect 6465 -7640 6470 -7604
rect 6425 -7674 6470 -7640
rect 6425 -7710 6431 -7674
rect 6465 -7710 6470 -7674
rect 6425 -7744 6470 -7710
rect 6425 -7780 6431 -7744
rect 6465 -7780 6470 -7744
rect 6286 -7864 6302 -7830
rect 6336 -7864 6352 -7830
rect 6425 -7898 6470 -7780
rect 6682 -7604 6727 -7362
rect 6941 -7186 6986 -6944
rect 7199 -6768 7244 -6526
rect 7199 -6804 7205 -6768
rect 7239 -6804 7244 -6768
rect 7199 -6838 7244 -6804
rect 7199 -6874 7205 -6838
rect 7239 -6874 7244 -6838
rect 7199 -6908 7244 -6874
rect 7199 -6944 7205 -6908
rect 7239 -6944 7244 -6908
rect 7060 -7028 7076 -6994
rect 7110 -7028 7126 -6994
rect 7060 -7136 7076 -7102
rect 7110 -7136 7126 -7102
rect 6941 -7222 6947 -7186
rect 6981 -7222 6986 -7186
rect 6941 -7256 6986 -7222
rect 6941 -7292 6947 -7256
rect 6981 -7292 6986 -7256
rect 6941 -7326 6986 -7292
rect 6941 -7362 6947 -7326
rect 6981 -7362 6986 -7326
rect 6802 -7446 6818 -7412
rect 6852 -7446 6868 -7412
rect 6802 -7554 6818 -7520
rect 6852 -7554 6868 -7520
rect 6682 -7640 6689 -7604
rect 6723 -7640 6727 -7604
rect 6682 -7674 6727 -7640
rect 6682 -7710 6689 -7674
rect 6723 -7710 6727 -7674
rect 6682 -7744 6727 -7710
rect 6682 -7780 6689 -7744
rect 6723 -7780 6727 -7744
rect 6544 -7864 6560 -7830
rect 6594 -7864 6610 -7830
rect 6682 -7898 6727 -7780
rect 6941 -7604 6986 -7362
rect 7199 -7186 7244 -6944
rect 7199 -7222 7205 -7186
rect 7239 -7222 7244 -7186
rect 7199 -7256 7244 -7222
rect 7199 -7292 7205 -7256
rect 7239 -7292 7244 -7256
rect 7199 -7326 7244 -7292
rect 7199 -7362 7205 -7326
rect 7239 -7362 7244 -7326
rect 7060 -7446 7076 -7412
rect 7110 -7446 7126 -7412
rect 7060 -7554 7076 -7520
rect 7110 -7554 7126 -7520
rect 6941 -7640 6947 -7604
rect 6981 -7640 6986 -7604
rect 6941 -7674 6986 -7640
rect 6941 -7710 6947 -7674
rect 6981 -7710 6986 -7674
rect 6941 -7744 6986 -7710
rect 6941 -7780 6947 -7744
rect 6981 -7780 6986 -7744
rect 6802 -7864 6818 -7830
rect 6852 -7864 6868 -7830
rect 6941 -7898 6986 -7780
rect 7199 -7604 7244 -7362
rect 7199 -7640 7205 -7604
rect 7239 -7640 7244 -7604
rect 7199 -7674 7244 -7640
rect 7199 -7710 7205 -7674
rect 7239 -7710 7244 -7674
rect 7199 -7744 7244 -7710
rect 7199 -7780 7205 -7744
rect 7239 -7780 7244 -7744
rect 7060 -7864 7076 -7830
rect 7110 -7864 7126 -7830
rect 7199 -7898 7244 -7780
rect 7805 -5096 7850 -5052
rect 7805 -5132 7811 -5096
rect 7845 -5132 7850 -5096
rect 7805 -5166 7850 -5132
rect 7805 -5202 7811 -5166
rect 7845 -5202 7850 -5166
rect 7805 -5236 7850 -5202
rect 7805 -5272 7811 -5236
rect 7845 -5272 7850 -5236
rect 7805 -5514 7850 -5272
rect 8063 -5096 8108 -5052
rect 8063 -5132 8069 -5096
rect 8103 -5132 8108 -5096
rect 8063 -5166 8108 -5132
rect 8063 -5202 8069 -5166
rect 8103 -5202 8108 -5166
rect 8063 -5236 8108 -5202
rect 8063 -5272 8069 -5236
rect 8103 -5272 8108 -5236
rect 7924 -5356 7940 -5322
rect 7974 -5356 7990 -5322
rect 7924 -5464 7940 -5430
rect 7974 -5464 7990 -5430
rect 7805 -5550 7811 -5514
rect 7845 -5550 7850 -5514
rect 7805 -5584 7850 -5550
rect 7805 -5620 7811 -5584
rect 7845 -5620 7850 -5584
rect 7805 -5654 7850 -5620
rect 7805 -5690 7811 -5654
rect 7845 -5690 7850 -5654
rect 7805 -5932 7850 -5690
rect 8063 -5514 8108 -5272
rect 8320 -5096 8365 -5052
rect 8320 -5132 8327 -5096
rect 8361 -5132 8365 -5096
rect 8320 -5166 8365 -5132
rect 8320 -5202 8327 -5166
rect 8361 -5202 8365 -5166
rect 8320 -5237 8365 -5202
rect 8320 -5273 8327 -5237
rect 8361 -5273 8365 -5237
rect 8182 -5356 8198 -5322
rect 8232 -5356 8248 -5322
rect 8182 -5464 8198 -5430
rect 8232 -5464 8248 -5430
rect 8063 -5550 8069 -5514
rect 8103 -5550 8108 -5514
rect 8063 -5584 8108 -5550
rect 8063 -5620 8069 -5584
rect 8103 -5620 8108 -5584
rect 8063 -5654 8108 -5620
rect 8063 -5690 8069 -5654
rect 8103 -5690 8108 -5654
rect 7924 -5774 7940 -5740
rect 7974 -5774 7990 -5740
rect 7924 -5882 7940 -5848
rect 7974 -5882 7990 -5848
rect 7805 -5968 7811 -5932
rect 7845 -5968 7850 -5932
rect 7805 -6002 7850 -5968
rect 7805 -6038 7811 -6002
rect 7845 -6038 7850 -6002
rect 7805 -6072 7850 -6038
rect 7805 -6108 7811 -6072
rect 7845 -6108 7850 -6072
rect 7805 -6350 7850 -6108
rect 8063 -5932 8108 -5690
rect 8320 -5514 8365 -5273
rect 8580 -5096 8625 -5052
rect 8580 -5132 8585 -5096
rect 8619 -5132 8625 -5096
rect 8580 -5166 8625 -5132
rect 8580 -5202 8585 -5166
rect 8619 -5202 8625 -5166
rect 8580 -5236 8625 -5202
rect 8580 -5272 8585 -5236
rect 8619 -5272 8625 -5236
rect 8440 -5356 8456 -5322
rect 8490 -5356 8506 -5322
rect 8440 -5464 8456 -5430
rect 8490 -5464 8506 -5430
rect 8320 -5550 8327 -5514
rect 8361 -5550 8365 -5514
rect 8320 -5584 8365 -5550
rect 8320 -5620 8327 -5584
rect 8361 -5620 8365 -5584
rect 8320 -5655 8365 -5620
rect 8320 -5691 8327 -5655
rect 8361 -5691 8365 -5655
rect 8182 -5774 8198 -5740
rect 8232 -5774 8248 -5740
rect 8182 -5882 8198 -5848
rect 8232 -5882 8248 -5848
rect 8063 -5968 8069 -5932
rect 8103 -5968 8108 -5932
rect 8063 -6002 8108 -5968
rect 8063 -6038 8069 -6002
rect 8103 -6038 8108 -6002
rect 8063 -6072 8108 -6038
rect 8063 -6108 8069 -6072
rect 8103 -6108 8108 -6072
rect 7924 -6192 7940 -6158
rect 7974 -6192 7990 -6158
rect 7924 -6300 7940 -6266
rect 7974 -6300 7990 -6266
rect 7805 -6386 7811 -6350
rect 7845 -6386 7850 -6350
rect 7805 -6420 7850 -6386
rect 7805 -6456 7811 -6420
rect 7845 -6456 7850 -6420
rect 7805 -6490 7850 -6456
rect 7805 -6526 7811 -6490
rect 7845 -6526 7850 -6490
rect 7805 -6768 7850 -6526
rect 8063 -6350 8108 -6108
rect 8320 -5932 8365 -5691
rect 8580 -5514 8625 -5272
rect 8838 -5096 8883 -5052
rect 8838 -5132 8843 -5096
rect 8877 -5132 8883 -5096
rect 8838 -5166 8883 -5132
rect 8838 -5202 8843 -5166
rect 8877 -5202 8883 -5166
rect 8838 -5236 8883 -5202
rect 8838 -5272 8843 -5236
rect 8877 -5272 8883 -5236
rect 8698 -5356 8714 -5322
rect 8748 -5356 8764 -5322
rect 8698 -5464 8714 -5430
rect 8748 -5464 8764 -5430
rect 8580 -5550 8585 -5514
rect 8619 -5550 8625 -5514
rect 8580 -5584 8625 -5550
rect 8580 -5620 8585 -5584
rect 8619 -5620 8625 -5584
rect 8580 -5654 8625 -5620
rect 8580 -5690 8585 -5654
rect 8619 -5690 8625 -5654
rect 8440 -5774 8456 -5740
rect 8490 -5774 8506 -5740
rect 8440 -5882 8456 -5848
rect 8490 -5882 8506 -5848
rect 8320 -5968 8327 -5932
rect 8361 -5968 8365 -5932
rect 8320 -6002 8365 -5968
rect 8320 -6038 8327 -6002
rect 8361 -6038 8365 -6002
rect 8320 -6073 8365 -6038
rect 8320 -6109 8327 -6073
rect 8361 -6109 8365 -6073
rect 8182 -6192 8198 -6158
rect 8232 -6192 8248 -6158
rect 8182 -6300 8198 -6266
rect 8232 -6300 8248 -6266
rect 8063 -6386 8069 -6350
rect 8103 -6386 8108 -6350
rect 8063 -6420 8108 -6386
rect 8063 -6456 8069 -6420
rect 8103 -6456 8108 -6420
rect 8063 -6490 8108 -6456
rect 8063 -6526 8069 -6490
rect 8103 -6526 8108 -6490
rect 7924 -6610 7940 -6576
rect 7974 -6610 7990 -6576
rect 7924 -6718 7940 -6684
rect 7974 -6718 7990 -6684
rect 7805 -6804 7811 -6768
rect 7845 -6804 7850 -6768
rect 7805 -6838 7850 -6804
rect 7805 -6874 7811 -6838
rect 7845 -6874 7850 -6838
rect 7805 -6908 7850 -6874
rect 7805 -6944 7811 -6908
rect 7845 -6944 7850 -6908
rect 7805 -7186 7850 -6944
rect 8063 -6768 8108 -6526
rect 8320 -6350 8365 -6109
rect 8580 -5932 8625 -5690
rect 8838 -5514 8883 -5272
rect 9095 -5096 9140 -5052
rect 9095 -5132 9101 -5096
rect 9135 -5132 9140 -5096
rect 9095 -5166 9140 -5132
rect 9095 -5202 9101 -5166
rect 9135 -5202 9140 -5166
rect 9095 -5236 9140 -5202
rect 9095 -5272 9101 -5236
rect 9135 -5272 9140 -5236
rect 8956 -5356 8972 -5322
rect 9006 -5356 9022 -5322
rect 8956 -5464 8972 -5430
rect 9006 -5464 9022 -5430
rect 8838 -5550 8843 -5514
rect 8877 -5550 8883 -5514
rect 8838 -5584 8883 -5550
rect 8838 -5620 8843 -5584
rect 8877 -5620 8883 -5584
rect 8838 -5654 8883 -5620
rect 8838 -5690 8843 -5654
rect 8877 -5690 8883 -5654
rect 8698 -5774 8714 -5740
rect 8748 -5774 8764 -5740
rect 8698 -5882 8714 -5848
rect 8748 -5882 8764 -5848
rect 8580 -5968 8585 -5932
rect 8619 -5968 8625 -5932
rect 8580 -6002 8625 -5968
rect 8580 -6038 8585 -6002
rect 8619 -6038 8625 -6002
rect 8580 -6072 8625 -6038
rect 8580 -6108 8585 -6072
rect 8619 -6108 8625 -6072
rect 8440 -6192 8456 -6158
rect 8490 -6192 8506 -6158
rect 8440 -6300 8456 -6266
rect 8490 -6300 8506 -6266
rect 8320 -6386 8327 -6350
rect 8361 -6386 8365 -6350
rect 8320 -6420 8365 -6386
rect 8320 -6456 8327 -6420
rect 8361 -6456 8365 -6420
rect 8320 -6491 8365 -6456
rect 8320 -6527 8327 -6491
rect 8361 -6527 8365 -6491
rect 8182 -6610 8198 -6576
rect 8232 -6610 8248 -6576
rect 8182 -6718 8198 -6684
rect 8232 -6718 8248 -6684
rect 8063 -6804 8069 -6768
rect 8103 -6804 8108 -6768
rect 8063 -6838 8108 -6804
rect 8063 -6874 8069 -6838
rect 8103 -6874 8108 -6838
rect 8063 -6908 8108 -6874
rect 8063 -6944 8069 -6908
rect 8103 -6944 8108 -6908
rect 7924 -7028 7940 -6994
rect 7974 -7028 7990 -6994
rect 7924 -7136 7940 -7102
rect 7974 -7136 7990 -7102
rect 7805 -7222 7811 -7186
rect 7845 -7222 7850 -7186
rect 7805 -7256 7850 -7222
rect 7805 -7292 7811 -7256
rect 7845 -7292 7850 -7256
rect 7805 -7326 7850 -7292
rect 7805 -7362 7811 -7326
rect 7845 -7362 7850 -7326
rect 7805 -7604 7850 -7362
rect 8063 -7186 8108 -6944
rect 8320 -6768 8365 -6527
rect 8580 -6350 8625 -6108
rect 8838 -5932 8883 -5690
rect 9095 -5514 9140 -5272
rect 9352 -5096 9397 -5052
rect 9352 -5132 9359 -5096
rect 9393 -5132 9397 -5096
rect 9352 -5166 9397 -5132
rect 9352 -5202 9359 -5166
rect 9393 -5202 9397 -5166
rect 9352 -5236 9397 -5202
rect 9352 -5272 9359 -5236
rect 9393 -5272 9397 -5236
rect 9214 -5356 9230 -5322
rect 9264 -5356 9280 -5322
rect 9214 -5464 9230 -5430
rect 9264 -5464 9280 -5430
rect 9095 -5550 9101 -5514
rect 9135 -5550 9140 -5514
rect 9095 -5584 9140 -5550
rect 9095 -5620 9101 -5584
rect 9135 -5620 9140 -5584
rect 9095 -5654 9140 -5620
rect 9095 -5690 9101 -5654
rect 9135 -5690 9140 -5654
rect 8956 -5774 8972 -5740
rect 9006 -5774 9022 -5740
rect 8956 -5882 8972 -5848
rect 9006 -5882 9022 -5848
rect 8838 -5968 8843 -5932
rect 8877 -5968 8883 -5932
rect 8838 -6002 8883 -5968
rect 8838 -6038 8843 -6002
rect 8877 -6038 8883 -6002
rect 8838 -6072 8883 -6038
rect 8838 -6108 8843 -6072
rect 8877 -6108 8883 -6072
rect 8698 -6192 8714 -6158
rect 8748 -6192 8764 -6158
rect 8698 -6300 8714 -6266
rect 8748 -6300 8764 -6266
rect 8580 -6386 8585 -6350
rect 8619 -6386 8625 -6350
rect 8580 -6420 8625 -6386
rect 8580 -6456 8585 -6420
rect 8619 -6456 8625 -6420
rect 8580 -6490 8625 -6456
rect 8580 -6526 8585 -6490
rect 8619 -6526 8625 -6490
rect 8440 -6610 8456 -6576
rect 8490 -6610 8506 -6576
rect 8440 -6718 8456 -6684
rect 8490 -6718 8506 -6684
rect 8320 -6804 8327 -6768
rect 8361 -6804 8365 -6768
rect 8320 -6838 8365 -6804
rect 8320 -6874 8327 -6838
rect 8361 -6874 8365 -6838
rect 8320 -6909 8365 -6874
rect 8320 -6945 8327 -6909
rect 8361 -6945 8365 -6909
rect 8182 -7028 8198 -6994
rect 8232 -7028 8248 -6994
rect 8182 -7136 8198 -7102
rect 8232 -7136 8248 -7102
rect 8063 -7222 8069 -7186
rect 8103 -7222 8108 -7186
rect 8063 -7256 8108 -7222
rect 8063 -7292 8069 -7256
rect 8103 -7292 8108 -7256
rect 8063 -7326 8108 -7292
rect 8063 -7362 8069 -7326
rect 8103 -7362 8108 -7326
rect 7924 -7446 7940 -7412
rect 7974 -7446 7990 -7412
rect 7924 -7554 7940 -7520
rect 7974 -7554 7990 -7520
rect 7805 -7640 7811 -7604
rect 7845 -7640 7850 -7604
rect 7805 -7674 7850 -7640
rect 7805 -7710 7811 -7674
rect 7845 -7710 7850 -7674
rect 7805 -7744 7850 -7710
rect 7805 -7780 7811 -7744
rect 7845 -7780 7850 -7744
rect 7805 -8022 7850 -7780
rect 8063 -7604 8108 -7362
rect 8320 -7186 8365 -6945
rect 8580 -6768 8625 -6526
rect 8838 -6350 8883 -6108
rect 9095 -5932 9140 -5690
rect 9352 -5514 9397 -5272
rect 9611 -5096 9656 -5052
rect 9611 -5132 9617 -5096
rect 9651 -5132 9656 -5096
rect 9611 -5166 9656 -5132
rect 9611 -5202 9617 -5166
rect 9651 -5202 9656 -5166
rect 9611 -5236 9656 -5202
rect 9611 -5272 9617 -5236
rect 9651 -5272 9656 -5236
rect 9472 -5356 9488 -5322
rect 9522 -5356 9538 -5322
rect 9472 -5464 9488 -5430
rect 9522 -5464 9538 -5430
rect 9352 -5550 9359 -5514
rect 9393 -5550 9397 -5514
rect 9352 -5584 9397 -5550
rect 9352 -5620 9359 -5584
rect 9393 -5620 9397 -5584
rect 9352 -5654 9397 -5620
rect 9352 -5690 9359 -5654
rect 9393 -5690 9397 -5654
rect 9214 -5774 9230 -5740
rect 9264 -5774 9280 -5740
rect 9214 -5882 9230 -5848
rect 9264 -5882 9280 -5848
rect 9095 -5968 9101 -5932
rect 9135 -5968 9140 -5932
rect 9095 -6002 9140 -5968
rect 9095 -6038 9101 -6002
rect 9135 -6038 9140 -6002
rect 9095 -6072 9140 -6038
rect 9095 -6108 9101 -6072
rect 9135 -6108 9140 -6072
rect 8956 -6192 8972 -6158
rect 9006 -6192 9022 -6158
rect 8956 -6300 8972 -6266
rect 9006 -6300 9022 -6266
rect 8838 -6386 8843 -6350
rect 8877 -6386 8883 -6350
rect 8838 -6420 8883 -6386
rect 8838 -6456 8843 -6420
rect 8877 -6456 8883 -6420
rect 8838 -6490 8883 -6456
rect 8838 -6526 8843 -6490
rect 8877 -6526 8883 -6490
rect 8698 -6610 8714 -6576
rect 8748 -6610 8764 -6576
rect 8698 -6718 8714 -6684
rect 8748 -6718 8764 -6684
rect 8580 -6804 8585 -6768
rect 8619 -6804 8625 -6768
rect 8580 -6838 8625 -6804
rect 8580 -6874 8585 -6838
rect 8619 -6874 8625 -6838
rect 8580 -6908 8625 -6874
rect 8580 -6944 8585 -6908
rect 8619 -6944 8625 -6908
rect 8440 -7028 8456 -6994
rect 8490 -7028 8506 -6994
rect 8440 -7136 8456 -7102
rect 8490 -7136 8506 -7102
rect 8320 -7222 8327 -7186
rect 8361 -7222 8365 -7186
rect 8320 -7256 8365 -7222
rect 8320 -7292 8327 -7256
rect 8361 -7292 8365 -7256
rect 8320 -7327 8365 -7292
rect 8320 -7363 8327 -7327
rect 8361 -7363 8365 -7327
rect 8182 -7446 8198 -7412
rect 8232 -7446 8248 -7412
rect 8182 -7554 8198 -7520
rect 8232 -7554 8248 -7520
rect 8063 -7640 8069 -7604
rect 8103 -7640 8108 -7604
rect 8063 -7674 8108 -7640
rect 8063 -7710 8069 -7674
rect 8103 -7710 8108 -7674
rect 8063 -7744 8108 -7710
rect 8063 -7780 8069 -7744
rect 8103 -7780 8108 -7744
rect 7924 -7864 7940 -7830
rect 7974 -7864 7990 -7830
rect 8063 -7898 8108 -7780
rect 8320 -7604 8365 -7363
rect 8580 -7186 8625 -6944
rect 8838 -6768 8883 -6526
rect 9095 -6350 9140 -6108
rect 9352 -5932 9397 -5690
rect 9611 -5514 9656 -5272
rect 9869 -5096 9914 -4910
rect 12528 -4911 12577 -4909
rect 10587 -5045 10603 -5011
rect 10637 -5045 10653 -5011
rect 10845 -5045 10861 -5011
rect 10895 -5045 10911 -5011
rect 11103 -5045 11119 -5011
rect 11153 -5045 11169 -5011
rect 11361 -5045 11377 -5011
rect 11411 -5045 11427 -5011
rect 11619 -5045 11635 -5011
rect 11669 -5045 11685 -5011
rect 11877 -5045 11893 -5011
rect 11927 -5045 11943 -5011
rect 12135 -5045 12151 -5011
rect 12185 -5045 12201 -5011
rect 12393 -5045 12409 -5011
rect 12443 -5045 12459 -5011
rect 9869 -5132 9875 -5096
rect 9909 -5132 9914 -5096
rect 9869 -5166 9914 -5132
rect 9869 -5202 9875 -5166
rect 9909 -5202 9914 -5166
rect 9869 -5236 9914 -5202
rect 9869 -5272 9875 -5236
rect 9909 -5272 9914 -5236
rect 9730 -5356 9746 -5322
rect 9780 -5356 9796 -5322
rect 9730 -5464 9746 -5430
rect 9780 -5464 9796 -5430
rect 9611 -5550 9617 -5514
rect 9651 -5550 9656 -5514
rect 9611 -5584 9656 -5550
rect 9611 -5620 9617 -5584
rect 9651 -5620 9656 -5584
rect 9611 -5654 9656 -5620
rect 9611 -5690 9617 -5654
rect 9651 -5690 9656 -5654
rect 9472 -5774 9488 -5740
rect 9522 -5774 9538 -5740
rect 9472 -5882 9488 -5848
rect 9522 -5882 9538 -5848
rect 9352 -5968 9359 -5932
rect 9393 -5968 9397 -5932
rect 9352 -6002 9397 -5968
rect 9352 -6038 9359 -6002
rect 9393 -6038 9397 -6002
rect 9352 -6072 9397 -6038
rect 9352 -6108 9359 -6072
rect 9393 -6108 9397 -6072
rect 9214 -6192 9230 -6158
rect 9264 -6192 9280 -6158
rect 9214 -6300 9230 -6266
rect 9264 -6300 9280 -6266
rect 9095 -6386 9101 -6350
rect 9135 -6386 9140 -6350
rect 9095 -6420 9140 -6386
rect 9095 -6456 9101 -6420
rect 9135 -6456 9140 -6420
rect 9095 -6490 9140 -6456
rect 9095 -6526 9101 -6490
rect 9135 -6526 9140 -6490
rect 8956 -6610 8972 -6576
rect 9006 -6610 9022 -6576
rect 8956 -6718 8972 -6684
rect 9006 -6718 9022 -6684
rect 8838 -6804 8843 -6768
rect 8877 -6804 8883 -6768
rect 8838 -6838 8883 -6804
rect 8838 -6874 8843 -6838
rect 8877 -6874 8883 -6838
rect 8838 -6908 8883 -6874
rect 8838 -6944 8843 -6908
rect 8877 -6944 8883 -6908
rect 8698 -7028 8714 -6994
rect 8748 -7028 8764 -6994
rect 8698 -7136 8714 -7102
rect 8748 -7136 8764 -7102
rect 8580 -7222 8585 -7186
rect 8619 -7222 8625 -7186
rect 8580 -7256 8625 -7222
rect 8580 -7292 8585 -7256
rect 8619 -7292 8625 -7256
rect 8580 -7326 8625 -7292
rect 8580 -7362 8585 -7326
rect 8619 -7362 8625 -7326
rect 8440 -7446 8456 -7412
rect 8490 -7446 8506 -7412
rect 8440 -7554 8456 -7520
rect 8490 -7554 8506 -7520
rect 8320 -7640 8327 -7604
rect 8361 -7640 8365 -7604
rect 8320 -7674 8365 -7640
rect 8320 -7710 8327 -7674
rect 8361 -7710 8365 -7674
rect 8320 -7745 8365 -7710
rect 8320 -7781 8327 -7745
rect 8361 -7781 8365 -7745
rect 8182 -7864 8198 -7830
rect 8232 -7864 8248 -7830
rect 8320 -7898 8365 -7781
rect 8580 -7604 8625 -7362
rect 8838 -7186 8883 -6944
rect 9095 -6768 9140 -6526
rect 9352 -6350 9397 -6108
rect 9611 -5932 9656 -5690
rect 9869 -5514 9914 -5272
rect 9869 -5550 9875 -5514
rect 9909 -5550 9914 -5514
rect 9869 -5584 9914 -5550
rect 9869 -5620 9875 -5584
rect 9909 -5620 9914 -5584
rect 9869 -5654 9914 -5620
rect 9869 -5690 9875 -5654
rect 9909 -5690 9914 -5654
rect 9730 -5774 9746 -5740
rect 9780 -5774 9796 -5740
rect 9730 -5882 9746 -5848
rect 9780 -5882 9796 -5848
rect 9611 -5968 9617 -5932
rect 9651 -5968 9656 -5932
rect 9611 -6002 9656 -5968
rect 9611 -6038 9617 -6002
rect 9651 -6038 9656 -6002
rect 9611 -6072 9656 -6038
rect 9611 -6108 9617 -6072
rect 9651 -6108 9656 -6072
rect 9472 -6192 9488 -6158
rect 9522 -6192 9538 -6158
rect 9472 -6300 9488 -6266
rect 9522 -6300 9538 -6266
rect 9352 -6386 9359 -6350
rect 9393 -6386 9397 -6350
rect 9352 -6420 9397 -6386
rect 9352 -6456 9359 -6420
rect 9393 -6456 9397 -6420
rect 9352 -6490 9397 -6456
rect 9352 -6526 9359 -6490
rect 9393 -6526 9397 -6490
rect 9214 -6610 9230 -6576
rect 9264 -6610 9280 -6576
rect 9214 -6718 9230 -6684
rect 9264 -6718 9280 -6684
rect 9095 -6804 9101 -6768
rect 9135 -6804 9140 -6768
rect 9095 -6838 9140 -6804
rect 9095 -6874 9101 -6838
rect 9135 -6874 9140 -6838
rect 9095 -6908 9140 -6874
rect 9095 -6944 9101 -6908
rect 9135 -6944 9140 -6908
rect 8956 -7028 8972 -6994
rect 9006 -7028 9022 -6994
rect 8956 -7136 8972 -7102
rect 9006 -7136 9022 -7102
rect 8838 -7222 8843 -7186
rect 8877 -7222 8883 -7186
rect 8838 -7256 8883 -7222
rect 8838 -7292 8843 -7256
rect 8877 -7292 8883 -7256
rect 8838 -7326 8883 -7292
rect 8838 -7362 8843 -7326
rect 8877 -7362 8883 -7326
rect 8698 -7446 8714 -7412
rect 8748 -7446 8764 -7412
rect 8698 -7554 8714 -7520
rect 8748 -7554 8764 -7520
rect 8580 -7640 8585 -7604
rect 8619 -7640 8625 -7604
rect 8580 -7674 8625 -7640
rect 8580 -7710 8585 -7674
rect 8619 -7710 8625 -7674
rect 8580 -7744 8625 -7710
rect 8580 -7780 8585 -7744
rect 8619 -7780 8625 -7744
rect 8440 -7864 8456 -7830
rect 8490 -7864 8506 -7830
rect 8580 -7898 8625 -7780
rect 8838 -7604 8883 -7362
rect 9095 -7186 9140 -6944
rect 9352 -6768 9397 -6526
rect 9611 -6350 9656 -6108
rect 9869 -5932 9914 -5690
rect 9869 -5968 9875 -5932
rect 9909 -5968 9914 -5932
rect 9869 -6002 9914 -5968
rect 9869 -6038 9875 -6002
rect 9909 -6038 9914 -6002
rect 9869 -6072 9914 -6038
rect 9869 -6108 9875 -6072
rect 9909 -6108 9914 -6072
rect 9730 -6192 9746 -6158
rect 9780 -6192 9796 -6158
rect 9730 -6300 9746 -6266
rect 9780 -6300 9796 -6266
rect 9611 -6386 9617 -6350
rect 9651 -6386 9656 -6350
rect 9611 -6420 9656 -6386
rect 9611 -6456 9617 -6420
rect 9651 -6456 9656 -6420
rect 9611 -6490 9656 -6456
rect 9611 -6526 9617 -6490
rect 9651 -6526 9656 -6490
rect 9472 -6610 9488 -6576
rect 9522 -6610 9538 -6576
rect 9472 -6718 9488 -6684
rect 9522 -6718 9538 -6684
rect 9352 -6804 9359 -6768
rect 9393 -6804 9397 -6768
rect 9352 -6838 9397 -6804
rect 9352 -6874 9359 -6838
rect 9393 -6874 9397 -6838
rect 9352 -6908 9397 -6874
rect 9352 -6944 9359 -6908
rect 9393 -6944 9397 -6908
rect 9214 -7028 9230 -6994
rect 9264 -7028 9280 -6994
rect 9214 -7136 9230 -7102
rect 9264 -7136 9280 -7102
rect 9095 -7222 9101 -7186
rect 9135 -7222 9140 -7186
rect 9095 -7256 9140 -7222
rect 9095 -7292 9101 -7256
rect 9135 -7292 9140 -7256
rect 9095 -7326 9140 -7292
rect 9095 -7362 9101 -7326
rect 9135 -7362 9140 -7326
rect 8956 -7446 8972 -7412
rect 9006 -7446 9022 -7412
rect 8956 -7554 8972 -7520
rect 9006 -7554 9022 -7520
rect 8838 -7640 8843 -7604
rect 8877 -7640 8883 -7604
rect 8838 -7674 8883 -7640
rect 8838 -7710 8843 -7674
rect 8877 -7710 8883 -7674
rect 8838 -7744 8883 -7710
rect 8838 -7780 8843 -7744
rect 8877 -7780 8883 -7744
rect 8698 -7864 8714 -7830
rect 8748 -7864 8764 -7830
rect 8838 -7898 8883 -7780
rect 9095 -7604 9140 -7362
rect 9352 -7186 9397 -6944
rect 9611 -6768 9656 -6526
rect 9869 -6350 9914 -6108
rect 9869 -6386 9875 -6350
rect 9909 -6386 9914 -6350
rect 9869 -6420 9914 -6386
rect 9869 -6456 9875 -6420
rect 9909 -6456 9914 -6420
rect 9869 -6490 9914 -6456
rect 9869 -6526 9875 -6490
rect 9909 -6526 9914 -6490
rect 9730 -6610 9746 -6576
rect 9780 -6610 9796 -6576
rect 9730 -6718 9746 -6684
rect 9780 -6718 9796 -6684
rect 9611 -6804 9617 -6768
rect 9651 -6804 9656 -6768
rect 9611 -6838 9656 -6804
rect 9611 -6874 9617 -6838
rect 9651 -6874 9656 -6838
rect 9611 -6908 9656 -6874
rect 9611 -6944 9617 -6908
rect 9651 -6944 9656 -6908
rect 9472 -7028 9488 -6994
rect 9522 -7028 9538 -6994
rect 9472 -7136 9488 -7102
rect 9522 -7136 9538 -7102
rect 9352 -7222 9359 -7186
rect 9393 -7222 9397 -7186
rect 9352 -7256 9397 -7222
rect 9352 -7292 9359 -7256
rect 9393 -7292 9397 -7256
rect 9352 -7326 9397 -7292
rect 9352 -7362 9359 -7326
rect 9393 -7362 9397 -7326
rect 9214 -7446 9230 -7412
rect 9264 -7446 9280 -7412
rect 9214 -7554 9230 -7520
rect 9264 -7554 9280 -7520
rect 9095 -7640 9101 -7604
rect 9135 -7640 9140 -7604
rect 9095 -7674 9140 -7640
rect 9095 -7710 9101 -7674
rect 9135 -7710 9140 -7674
rect 9095 -7744 9140 -7710
rect 9095 -7780 9101 -7744
rect 9135 -7780 9140 -7744
rect 8956 -7864 8972 -7830
rect 9006 -7864 9022 -7830
rect 9095 -7898 9140 -7780
rect 9352 -7604 9397 -7362
rect 9611 -7186 9656 -6944
rect 9869 -6768 9914 -6526
rect 9869 -6804 9875 -6768
rect 9909 -6804 9914 -6768
rect 9869 -6838 9914 -6804
rect 9869 -6874 9875 -6838
rect 9909 -6874 9914 -6838
rect 9869 -6908 9914 -6874
rect 9869 -6944 9875 -6908
rect 9909 -6944 9914 -6908
rect 9730 -7028 9746 -6994
rect 9780 -7028 9796 -6994
rect 9730 -7136 9746 -7102
rect 9780 -7136 9796 -7102
rect 9611 -7222 9617 -7186
rect 9651 -7222 9656 -7186
rect 9611 -7256 9656 -7222
rect 9611 -7292 9617 -7256
rect 9651 -7292 9656 -7256
rect 9611 -7326 9656 -7292
rect 9611 -7362 9617 -7326
rect 9651 -7362 9656 -7326
rect 9472 -7446 9488 -7412
rect 9522 -7446 9538 -7412
rect 9472 -7554 9488 -7520
rect 9522 -7554 9538 -7520
rect 9352 -7640 9359 -7604
rect 9393 -7640 9397 -7604
rect 9352 -7674 9397 -7640
rect 9352 -7710 9359 -7674
rect 9393 -7710 9397 -7674
rect 9352 -7744 9397 -7710
rect 9352 -7780 9359 -7744
rect 9393 -7780 9397 -7744
rect 9214 -7864 9230 -7830
rect 9264 -7864 9280 -7830
rect 9352 -7898 9397 -7780
rect 9611 -7604 9656 -7362
rect 9869 -7186 9914 -6944
rect 9869 -7222 9875 -7186
rect 9909 -7222 9914 -7186
rect 9869 -7256 9914 -7222
rect 9869 -7292 9875 -7256
rect 9909 -7292 9914 -7256
rect 9869 -7326 9914 -7292
rect 9869 -7362 9875 -7326
rect 9909 -7362 9914 -7326
rect 9730 -7446 9746 -7412
rect 9780 -7446 9796 -7412
rect 9730 -7554 9746 -7520
rect 9780 -7554 9796 -7520
rect 9611 -7640 9617 -7604
rect 9651 -7640 9656 -7604
rect 9611 -7674 9656 -7640
rect 9611 -7710 9617 -7674
rect 9651 -7710 9656 -7674
rect 9611 -7744 9656 -7710
rect 9611 -7780 9617 -7744
rect 9651 -7780 9656 -7744
rect 9472 -7864 9488 -7830
rect 9522 -7864 9538 -7830
rect 9611 -7898 9656 -7780
rect 9869 -7604 9914 -7362
rect 9869 -7640 9875 -7604
rect 9909 -7640 9914 -7604
rect 9869 -7674 9914 -7640
rect 9869 -7710 9875 -7674
rect 9909 -7710 9914 -7674
rect 9869 -7744 9914 -7710
rect 9869 -7780 9875 -7744
rect 9909 -7780 9914 -7744
rect 9730 -7864 9746 -7830
rect 9780 -7864 9796 -7830
rect 9869 -7898 9914 -7780
rect 10468 -5095 10513 -5051
rect 10468 -5131 10474 -5095
rect 10508 -5131 10513 -5095
rect 10468 -5165 10513 -5131
rect 10468 -5201 10474 -5165
rect 10508 -5201 10513 -5165
rect 10468 -5235 10513 -5201
rect 10468 -5271 10474 -5235
rect 10508 -5271 10513 -5235
rect 10468 -5513 10513 -5271
rect 10726 -5095 10771 -5051
rect 10726 -5131 10732 -5095
rect 10766 -5131 10771 -5095
rect 10726 -5165 10771 -5131
rect 10726 -5201 10732 -5165
rect 10766 -5201 10771 -5165
rect 10726 -5235 10771 -5201
rect 10726 -5271 10732 -5235
rect 10766 -5271 10771 -5235
rect 10587 -5355 10603 -5321
rect 10637 -5355 10653 -5321
rect 10587 -5463 10603 -5429
rect 10637 -5463 10653 -5429
rect 10468 -5549 10474 -5513
rect 10508 -5549 10513 -5513
rect 10468 -5583 10513 -5549
rect 10468 -5619 10474 -5583
rect 10508 -5619 10513 -5583
rect 10468 -5653 10513 -5619
rect 10468 -5689 10474 -5653
rect 10508 -5689 10513 -5653
rect 10468 -5931 10513 -5689
rect 10726 -5513 10771 -5271
rect 10983 -5095 11028 -5051
rect 10983 -5131 10990 -5095
rect 11024 -5131 11028 -5095
rect 10983 -5165 11028 -5131
rect 10983 -5201 10990 -5165
rect 11024 -5201 11028 -5165
rect 10983 -5236 11028 -5201
rect 10983 -5272 10990 -5236
rect 11024 -5272 11028 -5236
rect 10845 -5355 10861 -5321
rect 10895 -5355 10911 -5321
rect 10845 -5463 10861 -5429
rect 10895 -5463 10911 -5429
rect 10726 -5549 10732 -5513
rect 10766 -5549 10771 -5513
rect 10726 -5583 10771 -5549
rect 10726 -5619 10732 -5583
rect 10766 -5619 10771 -5583
rect 10726 -5653 10771 -5619
rect 10726 -5689 10732 -5653
rect 10766 -5689 10771 -5653
rect 10587 -5773 10603 -5739
rect 10637 -5773 10653 -5739
rect 10587 -5881 10603 -5847
rect 10637 -5881 10653 -5847
rect 10468 -5967 10474 -5931
rect 10508 -5967 10513 -5931
rect 10468 -6001 10513 -5967
rect 10468 -6037 10474 -6001
rect 10508 -6037 10513 -6001
rect 10468 -6071 10513 -6037
rect 10468 -6107 10474 -6071
rect 10508 -6107 10513 -6071
rect 10468 -6349 10513 -6107
rect 10726 -5931 10771 -5689
rect 10983 -5513 11028 -5272
rect 11243 -5095 11288 -5051
rect 11243 -5131 11248 -5095
rect 11282 -5131 11288 -5095
rect 11243 -5165 11288 -5131
rect 11243 -5201 11248 -5165
rect 11282 -5201 11288 -5165
rect 11243 -5235 11288 -5201
rect 11243 -5271 11248 -5235
rect 11282 -5271 11288 -5235
rect 11103 -5355 11119 -5321
rect 11153 -5355 11169 -5321
rect 11103 -5463 11119 -5429
rect 11153 -5463 11169 -5429
rect 10983 -5549 10990 -5513
rect 11024 -5549 11028 -5513
rect 10983 -5583 11028 -5549
rect 10983 -5619 10990 -5583
rect 11024 -5619 11028 -5583
rect 10983 -5654 11028 -5619
rect 10983 -5690 10990 -5654
rect 11024 -5690 11028 -5654
rect 10845 -5773 10861 -5739
rect 10895 -5773 10911 -5739
rect 10845 -5881 10861 -5847
rect 10895 -5881 10911 -5847
rect 10726 -5967 10732 -5931
rect 10766 -5967 10771 -5931
rect 10726 -6001 10771 -5967
rect 10726 -6037 10732 -6001
rect 10766 -6037 10771 -6001
rect 10726 -6071 10771 -6037
rect 10726 -6107 10732 -6071
rect 10766 -6107 10771 -6071
rect 10587 -6191 10603 -6157
rect 10637 -6191 10653 -6157
rect 10587 -6299 10603 -6265
rect 10637 -6299 10653 -6265
rect 10468 -6385 10474 -6349
rect 10508 -6385 10513 -6349
rect 10468 -6419 10513 -6385
rect 10468 -6455 10474 -6419
rect 10508 -6455 10513 -6419
rect 10468 -6489 10513 -6455
rect 10468 -6525 10474 -6489
rect 10508 -6525 10513 -6489
rect 10468 -6767 10513 -6525
rect 10726 -6349 10771 -6107
rect 10983 -5931 11028 -5690
rect 11243 -5513 11288 -5271
rect 11501 -5095 11546 -5051
rect 11501 -5131 11506 -5095
rect 11540 -5131 11546 -5095
rect 11501 -5165 11546 -5131
rect 11501 -5201 11506 -5165
rect 11540 -5201 11546 -5165
rect 11501 -5235 11546 -5201
rect 11501 -5271 11506 -5235
rect 11540 -5271 11546 -5235
rect 11361 -5355 11377 -5321
rect 11411 -5355 11427 -5321
rect 11361 -5463 11377 -5429
rect 11411 -5463 11427 -5429
rect 11243 -5549 11248 -5513
rect 11282 -5549 11288 -5513
rect 11243 -5583 11288 -5549
rect 11243 -5619 11248 -5583
rect 11282 -5619 11288 -5583
rect 11243 -5653 11288 -5619
rect 11243 -5689 11248 -5653
rect 11282 -5689 11288 -5653
rect 11103 -5773 11119 -5739
rect 11153 -5773 11169 -5739
rect 11103 -5881 11119 -5847
rect 11153 -5881 11169 -5847
rect 10983 -5967 10990 -5931
rect 11024 -5967 11028 -5931
rect 10983 -6001 11028 -5967
rect 10983 -6037 10990 -6001
rect 11024 -6037 11028 -6001
rect 10983 -6072 11028 -6037
rect 10983 -6108 10990 -6072
rect 11024 -6108 11028 -6072
rect 10845 -6191 10861 -6157
rect 10895 -6191 10911 -6157
rect 10845 -6299 10861 -6265
rect 10895 -6299 10911 -6265
rect 10726 -6385 10732 -6349
rect 10766 -6385 10771 -6349
rect 10726 -6419 10771 -6385
rect 10726 -6455 10732 -6419
rect 10766 -6455 10771 -6419
rect 10726 -6489 10771 -6455
rect 10726 -6525 10732 -6489
rect 10766 -6525 10771 -6489
rect 10587 -6609 10603 -6575
rect 10637 -6609 10653 -6575
rect 10587 -6717 10603 -6683
rect 10637 -6717 10653 -6683
rect 10468 -6803 10474 -6767
rect 10508 -6803 10513 -6767
rect 10468 -6837 10513 -6803
rect 10468 -6873 10474 -6837
rect 10508 -6873 10513 -6837
rect 10468 -6907 10513 -6873
rect 10468 -6943 10474 -6907
rect 10508 -6943 10513 -6907
rect 10468 -7185 10513 -6943
rect 10726 -6767 10771 -6525
rect 10983 -6349 11028 -6108
rect 11243 -5931 11288 -5689
rect 11501 -5513 11546 -5271
rect 11758 -5095 11803 -5051
rect 11758 -5131 11764 -5095
rect 11798 -5131 11803 -5095
rect 11758 -5165 11803 -5131
rect 11758 -5201 11764 -5165
rect 11798 -5201 11803 -5165
rect 11758 -5235 11803 -5201
rect 11758 -5271 11764 -5235
rect 11798 -5271 11803 -5235
rect 11619 -5355 11635 -5321
rect 11669 -5355 11685 -5321
rect 11619 -5463 11635 -5429
rect 11669 -5463 11685 -5429
rect 11501 -5549 11506 -5513
rect 11540 -5549 11546 -5513
rect 11501 -5583 11546 -5549
rect 11501 -5619 11506 -5583
rect 11540 -5619 11546 -5583
rect 11501 -5653 11546 -5619
rect 11501 -5689 11506 -5653
rect 11540 -5689 11546 -5653
rect 11361 -5773 11377 -5739
rect 11411 -5773 11427 -5739
rect 11361 -5881 11377 -5847
rect 11411 -5881 11427 -5847
rect 11243 -5967 11248 -5931
rect 11282 -5967 11288 -5931
rect 11243 -6001 11288 -5967
rect 11243 -6037 11248 -6001
rect 11282 -6037 11288 -6001
rect 11243 -6071 11288 -6037
rect 11243 -6107 11248 -6071
rect 11282 -6107 11288 -6071
rect 11103 -6191 11119 -6157
rect 11153 -6191 11169 -6157
rect 11103 -6299 11119 -6265
rect 11153 -6299 11169 -6265
rect 10983 -6385 10990 -6349
rect 11024 -6385 11028 -6349
rect 10983 -6419 11028 -6385
rect 10983 -6455 10990 -6419
rect 11024 -6455 11028 -6419
rect 10983 -6490 11028 -6455
rect 10983 -6526 10990 -6490
rect 11024 -6526 11028 -6490
rect 10845 -6609 10861 -6575
rect 10895 -6609 10911 -6575
rect 10845 -6717 10861 -6683
rect 10895 -6717 10911 -6683
rect 10726 -6803 10732 -6767
rect 10766 -6803 10771 -6767
rect 10726 -6837 10771 -6803
rect 10726 -6873 10732 -6837
rect 10766 -6873 10771 -6837
rect 10726 -6907 10771 -6873
rect 10726 -6943 10732 -6907
rect 10766 -6943 10771 -6907
rect 10587 -7027 10603 -6993
rect 10637 -7027 10653 -6993
rect 10587 -7135 10603 -7101
rect 10637 -7135 10653 -7101
rect 10468 -7221 10474 -7185
rect 10508 -7221 10513 -7185
rect 10468 -7255 10513 -7221
rect 10468 -7291 10474 -7255
rect 10508 -7291 10513 -7255
rect 10468 -7325 10513 -7291
rect 10468 -7361 10474 -7325
rect 10508 -7361 10513 -7325
rect 10468 -7603 10513 -7361
rect 10726 -7185 10771 -6943
rect 10983 -6767 11028 -6526
rect 11243 -6349 11288 -6107
rect 11501 -5931 11546 -5689
rect 11758 -5513 11803 -5271
rect 12015 -5095 12060 -5051
rect 12015 -5131 12022 -5095
rect 12056 -5131 12060 -5095
rect 12015 -5165 12060 -5131
rect 12015 -5201 12022 -5165
rect 12056 -5201 12060 -5165
rect 12015 -5235 12060 -5201
rect 12015 -5271 12022 -5235
rect 12056 -5271 12060 -5235
rect 11877 -5355 11893 -5321
rect 11927 -5355 11943 -5321
rect 11877 -5463 11893 -5429
rect 11927 -5463 11943 -5429
rect 11758 -5549 11764 -5513
rect 11798 -5549 11803 -5513
rect 11758 -5583 11803 -5549
rect 11758 -5619 11764 -5583
rect 11798 -5619 11803 -5583
rect 11758 -5653 11803 -5619
rect 11758 -5689 11764 -5653
rect 11798 -5689 11803 -5653
rect 11619 -5773 11635 -5739
rect 11669 -5773 11685 -5739
rect 11619 -5881 11635 -5847
rect 11669 -5881 11685 -5847
rect 11501 -5967 11506 -5931
rect 11540 -5967 11546 -5931
rect 11501 -6001 11546 -5967
rect 11501 -6037 11506 -6001
rect 11540 -6037 11546 -6001
rect 11501 -6071 11546 -6037
rect 11501 -6107 11506 -6071
rect 11540 -6107 11546 -6071
rect 11361 -6191 11377 -6157
rect 11411 -6191 11427 -6157
rect 11361 -6299 11377 -6265
rect 11411 -6299 11427 -6265
rect 11243 -6385 11248 -6349
rect 11282 -6385 11288 -6349
rect 11243 -6419 11288 -6385
rect 11243 -6455 11248 -6419
rect 11282 -6455 11288 -6419
rect 11243 -6489 11288 -6455
rect 11243 -6525 11248 -6489
rect 11282 -6525 11288 -6489
rect 11103 -6609 11119 -6575
rect 11153 -6609 11169 -6575
rect 11103 -6717 11119 -6683
rect 11153 -6717 11169 -6683
rect 10983 -6803 10990 -6767
rect 11024 -6803 11028 -6767
rect 10983 -6837 11028 -6803
rect 10983 -6873 10990 -6837
rect 11024 -6873 11028 -6837
rect 10983 -6908 11028 -6873
rect 10983 -6944 10990 -6908
rect 11024 -6944 11028 -6908
rect 10845 -7027 10861 -6993
rect 10895 -7027 10911 -6993
rect 10845 -7135 10861 -7101
rect 10895 -7135 10911 -7101
rect 10726 -7221 10732 -7185
rect 10766 -7221 10771 -7185
rect 10726 -7255 10771 -7221
rect 10726 -7291 10732 -7255
rect 10766 -7291 10771 -7255
rect 10726 -7325 10771 -7291
rect 10726 -7361 10732 -7325
rect 10766 -7361 10771 -7325
rect 10587 -7445 10603 -7411
rect 10637 -7445 10653 -7411
rect 10587 -7553 10603 -7519
rect 10637 -7553 10653 -7519
rect 10468 -7639 10474 -7603
rect 10508 -7639 10513 -7603
rect 10468 -7673 10513 -7639
rect 10468 -7709 10474 -7673
rect 10508 -7709 10513 -7673
rect 10468 -7743 10513 -7709
rect 10468 -7779 10474 -7743
rect 10508 -7779 10513 -7743
rect 10468 -8021 10513 -7779
rect 10726 -7603 10771 -7361
rect 10983 -7185 11028 -6944
rect 11243 -6767 11288 -6525
rect 11501 -6349 11546 -6107
rect 11758 -5931 11803 -5689
rect 12015 -5513 12060 -5271
rect 12274 -5095 12319 -5051
rect 12274 -5131 12280 -5095
rect 12314 -5131 12319 -5095
rect 12274 -5165 12319 -5131
rect 12274 -5201 12280 -5165
rect 12314 -5201 12319 -5165
rect 12274 -5235 12319 -5201
rect 12274 -5271 12280 -5235
rect 12314 -5271 12319 -5235
rect 12135 -5355 12151 -5321
rect 12185 -5355 12201 -5321
rect 12135 -5463 12151 -5429
rect 12185 -5463 12201 -5429
rect 12015 -5549 12022 -5513
rect 12056 -5549 12060 -5513
rect 12015 -5583 12060 -5549
rect 12015 -5619 12022 -5583
rect 12056 -5619 12060 -5583
rect 12015 -5653 12060 -5619
rect 12015 -5689 12022 -5653
rect 12056 -5689 12060 -5653
rect 11877 -5773 11893 -5739
rect 11927 -5773 11943 -5739
rect 11877 -5881 11893 -5847
rect 11927 -5881 11943 -5847
rect 11758 -5967 11764 -5931
rect 11798 -5967 11803 -5931
rect 11758 -6001 11803 -5967
rect 11758 -6037 11764 -6001
rect 11798 -6037 11803 -6001
rect 11758 -6071 11803 -6037
rect 11758 -6107 11764 -6071
rect 11798 -6107 11803 -6071
rect 11619 -6191 11635 -6157
rect 11669 -6191 11685 -6157
rect 11619 -6299 11635 -6265
rect 11669 -6299 11685 -6265
rect 11501 -6385 11506 -6349
rect 11540 -6385 11546 -6349
rect 11501 -6419 11546 -6385
rect 11501 -6455 11506 -6419
rect 11540 -6455 11546 -6419
rect 11501 -6489 11546 -6455
rect 11501 -6525 11506 -6489
rect 11540 -6525 11546 -6489
rect 11361 -6609 11377 -6575
rect 11411 -6609 11427 -6575
rect 11361 -6717 11377 -6683
rect 11411 -6717 11427 -6683
rect 11243 -6803 11248 -6767
rect 11282 -6803 11288 -6767
rect 11243 -6837 11288 -6803
rect 11243 -6873 11248 -6837
rect 11282 -6873 11288 -6837
rect 11243 -6907 11288 -6873
rect 11243 -6943 11248 -6907
rect 11282 -6943 11288 -6907
rect 11103 -7027 11119 -6993
rect 11153 -7027 11169 -6993
rect 11103 -7135 11119 -7101
rect 11153 -7135 11169 -7101
rect 10983 -7221 10990 -7185
rect 11024 -7221 11028 -7185
rect 10983 -7255 11028 -7221
rect 10983 -7291 10990 -7255
rect 11024 -7291 11028 -7255
rect 10983 -7326 11028 -7291
rect 10983 -7362 10990 -7326
rect 11024 -7362 11028 -7326
rect 10845 -7445 10861 -7411
rect 10895 -7445 10911 -7411
rect 10845 -7553 10861 -7519
rect 10895 -7553 10911 -7519
rect 10726 -7639 10732 -7603
rect 10766 -7639 10771 -7603
rect 10726 -7673 10771 -7639
rect 10726 -7709 10732 -7673
rect 10766 -7709 10771 -7673
rect 10726 -7743 10771 -7709
rect 10726 -7779 10732 -7743
rect 10766 -7779 10771 -7743
rect 10587 -7863 10603 -7829
rect 10637 -7863 10653 -7829
rect 10726 -7897 10771 -7779
rect 10983 -7603 11028 -7362
rect 11243 -7185 11288 -6943
rect 11501 -6767 11546 -6525
rect 11758 -6349 11803 -6107
rect 12015 -5931 12060 -5689
rect 12274 -5513 12319 -5271
rect 12532 -5095 12577 -4911
rect 12532 -5131 12538 -5095
rect 12572 -5131 12577 -5095
rect 12532 -5165 12577 -5131
rect 12532 -5201 12538 -5165
rect 12572 -5201 12577 -5165
rect 12532 -5235 12577 -5201
rect 12532 -5271 12538 -5235
rect 12572 -5271 12577 -5235
rect 12393 -5355 12409 -5321
rect 12443 -5355 12459 -5321
rect 12393 -5463 12409 -5429
rect 12443 -5463 12459 -5429
rect 12274 -5549 12280 -5513
rect 12314 -5549 12319 -5513
rect 12274 -5583 12319 -5549
rect 12274 -5619 12280 -5583
rect 12314 -5619 12319 -5583
rect 12274 -5653 12319 -5619
rect 12274 -5689 12280 -5653
rect 12314 -5689 12319 -5653
rect 12135 -5773 12151 -5739
rect 12185 -5773 12201 -5739
rect 12135 -5881 12151 -5847
rect 12185 -5881 12201 -5847
rect 12015 -5967 12022 -5931
rect 12056 -5967 12060 -5931
rect 12015 -6001 12060 -5967
rect 12015 -6037 12022 -6001
rect 12056 -6037 12060 -6001
rect 12015 -6071 12060 -6037
rect 12015 -6107 12022 -6071
rect 12056 -6107 12060 -6071
rect 11877 -6191 11893 -6157
rect 11927 -6191 11943 -6157
rect 11877 -6299 11893 -6265
rect 11927 -6299 11943 -6265
rect 11758 -6385 11764 -6349
rect 11798 -6385 11803 -6349
rect 11758 -6419 11803 -6385
rect 11758 -6455 11764 -6419
rect 11798 -6455 11803 -6419
rect 11758 -6489 11803 -6455
rect 11758 -6525 11764 -6489
rect 11798 -6525 11803 -6489
rect 11619 -6609 11635 -6575
rect 11669 -6609 11685 -6575
rect 11619 -6717 11635 -6683
rect 11669 -6717 11685 -6683
rect 11501 -6803 11506 -6767
rect 11540 -6803 11546 -6767
rect 11501 -6837 11546 -6803
rect 11501 -6873 11506 -6837
rect 11540 -6873 11546 -6837
rect 11501 -6907 11546 -6873
rect 11501 -6943 11506 -6907
rect 11540 -6943 11546 -6907
rect 11361 -7027 11377 -6993
rect 11411 -7027 11427 -6993
rect 11361 -7135 11377 -7101
rect 11411 -7135 11427 -7101
rect 11243 -7221 11248 -7185
rect 11282 -7221 11288 -7185
rect 11243 -7255 11288 -7221
rect 11243 -7291 11248 -7255
rect 11282 -7291 11288 -7255
rect 11243 -7325 11288 -7291
rect 11243 -7361 11248 -7325
rect 11282 -7361 11288 -7325
rect 11103 -7445 11119 -7411
rect 11153 -7445 11169 -7411
rect 11103 -7553 11119 -7519
rect 11153 -7553 11169 -7519
rect 10983 -7639 10990 -7603
rect 11024 -7639 11028 -7603
rect 10983 -7673 11028 -7639
rect 10983 -7709 10990 -7673
rect 11024 -7709 11028 -7673
rect 10983 -7744 11028 -7709
rect 10983 -7780 10990 -7744
rect 11024 -7780 11028 -7744
rect 10845 -7863 10861 -7829
rect 10895 -7863 10911 -7829
rect 10983 -7897 11028 -7780
rect 11243 -7603 11288 -7361
rect 11501 -7185 11546 -6943
rect 11758 -6767 11803 -6525
rect 12015 -6349 12060 -6107
rect 12274 -5931 12319 -5689
rect 12532 -5513 12577 -5271
rect 12532 -5549 12538 -5513
rect 12572 -5549 12577 -5513
rect 12532 -5583 12577 -5549
rect 12532 -5619 12538 -5583
rect 12572 -5619 12577 -5583
rect 12532 -5653 12577 -5619
rect 12532 -5689 12538 -5653
rect 12572 -5689 12577 -5653
rect 12393 -5773 12409 -5739
rect 12443 -5773 12459 -5739
rect 12393 -5881 12409 -5847
rect 12443 -5881 12459 -5847
rect 12274 -5967 12280 -5931
rect 12314 -5967 12319 -5931
rect 12274 -6001 12319 -5967
rect 12274 -6037 12280 -6001
rect 12314 -6037 12319 -6001
rect 12274 -6071 12319 -6037
rect 12274 -6107 12280 -6071
rect 12314 -6107 12319 -6071
rect 12135 -6191 12151 -6157
rect 12185 -6191 12201 -6157
rect 12135 -6299 12151 -6265
rect 12185 -6299 12201 -6265
rect 12015 -6385 12022 -6349
rect 12056 -6385 12060 -6349
rect 12015 -6419 12060 -6385
rect 12015 -6455 12022 -6419
rect 12056 -6455 12060 -6419
rect 12015 -6489 12060 -6455
rect 12015 -6525 12022 -6489
rect 12056 -6525 12060 -6489
rect 11877 -6609 11893 -6575
rect 11927 -6609 11943 -6575
rect 11877 -6717 11893 -6683
rect 11927 -6717 11943 -6683
rect 11758 -6803 11764 -6767
rect 11798 -6803 11803 -6767
rect 11758 -6837 11803 -6803
rect 11758 -6873 11764 -6837
rect 11798 -6873 11803 -6837
rect 11758 -6907 11803 -6873
rect 11758 -6943 11764 -6907
rect 11798 -6943 11803 -6907
rect 11619 -7027 11635 -6993
rect 11669 -7027 11685 -6993
rect 11619 -7135 11635 -7101
rect 11669 -7135 11685 -7101
rect 11501 -7221 11506 -7185
rect 11540 -7221 11546 -7185
rect 11501 -7255 11546 -7221
rect 11501 -7291 11506 -7255
rect 11540 -7291 11546 -7255
rect 11501 -7325 11546 -7291
rect 11501 -7361 11506 -7325
rect 11540 -7361 11546 -7325
rect 11361 -7445 11377 -7411
rect 11411 -7445 11427 -7411
rect 11361 -7553 11377 -7519
rect 11411 -7553 11427 -7519
rect 11243 -7639 11248 -7603
rect 11282 -7639 11288 -7603
rect 11243 -7673 11288 -7639
rect 11243 -7709 11248 -7673
rect 11282 -7709 11288 -7673
rect 11243 -7743 11288 -7709
rect 11243 -7779 11248 -7743
rect 11282 -7779 11288 -7743
rect 11103 -7863 11119 -7829
rect 11153 -7863 11169 -7829
rect 11243 -7897 11288 -7779
rect 11501 -7603 11546 -7361
rect 11758 -7185 11803 -6943
rect 12015 -6767 12060 -6525
rect 12274 -6349 12319 -6107
rect 12532 -5931 12577 -5689
rect 12532 -5967 12538 -5931
rect 12572 -5967 12577 -5931
rect 12532 -6001 12577 -5967
rect 12532 -6037 12538 -6001
rect 12572 -6037 12577 -6001
rect 12532 -6071 12577 -6037
rect 12532 -6107 12538 -6071
rect 12572 -6107 12577 -6071
rect 12393 -6191 12409 -6157
rect 12443 -6191 12459 -6157
rect 12393 -6299 12409 -6265
rect 12443 -6299 12459 -6265
rect 12274 -6385 12280 -6349
rect 12314 -6385 12319 -6349
rect 12274 -6419 12319 -6385
rect 12274 -6455 12280 -6419
rect 12314 -6455 12319 -6419
rect 12274 -6489 12319 -6455
rect 12274 -6525 12280 -6489
rect 12314 -6525 12319 -6489
rect 12135 -6609 12151 -6575
rect 12185 -6609 12201 -6575
rect 12135 -6717 12151 -6683
rect 12185 -6717 12201 -6683
rect 12015 -6803 12022 -6767
rect 12056 -6803 12060 -6767
rect 12015 -6837 12060 -6803
rect 12015 -6873 12022 -6837
rect 12056 -6873 12060 -6837
rect 12015 -6907 12060 -6873
rect 12015 -6943 12022 -6907
rect 12056 -6943 12060 -6907
rect 11877 -7027 11893 -6993
rect 11927 -7027 11943 -6993
rect 11877 -7135 11893 -7101
rect 11927 -7135 11943 -7101
rect 11758 -7221 11764 -7185
rect 11798 -7221 11803 -7185
rect 11758 -7255 11803 -7221
rect 11758 -7291 11764 -7255
rect 11798 -7291 11803 -7255
rect 11758 -7325 11803 -7291
rect 11758 -7361 11764 -7325
rect 11798 -7361 11803 -7325
rect 11619 -7445 11635 -7411
rect 11669 -7445 11685 -7411
rect 11619 -7553 11635 -7519
rect 11669 -7553 11685 -7519
rect 11501 -7639 11506 -7603
rect 11540 -7639 11546 -7603
rect 11501 -7673 11546 -7639
rect 11501 -7709 11506 -7673
rect 11540 -7709 11546 -7673
rect 11501 -7743 11546 -7709
rect 11501 -7779 11506 -7743
rect 11540 -7779 11546 -7743
rect 11361 -7863 11377 -7829
rect 11411 -7863 11427 -7829
rect 11501 -7897 11546 -7779
rect 11758 -7603 11803 -7361
rect 12015 -7185 12060 -6943
rect 12274 -6767 12319 -6525
rect 12532 -6349 12577 -6107
rect 12532 -6385 12538 -6349
rect 12572 -6385 12577 -6349
rect 12532 -6419 12577 -6385
rect 12532 -6455 12538 -6419
rect 12572 -6455 12577 -6419
rect 12532 -6489 12577 -6455
rect 12532 -6525 12538 -6489
rect 12572 -6525 12577 -6489
rect 12393 -6609 12409 -6575
rect 12443 -6609 12459 -6575
rect 12393 -6717 12409 -6683
rect 12443 -6717 12459 -6683
rect 12274 -6803 12280 -6767
rect 12314 -6803 12319 -6767
rect 12274 -6837 12319 -6803
rect 12274 -6873 12280 -6837
rect 12314 -6873 12319 -6837
rect 12274 -6907 12319 -6873
rect 12274 -6943 12280 -6907
rect 12314 -6943 12319 -6907
rect 12135 -7027 12151 -6993
rect 12185 -7027 12201 -6993
rect 12135 -7135 12151 -7101
rect 12185 -7135 12201 -7101
rect 12015 -7221 12022 -7185
rect 12056 -7221 12060 -7185
rect 12015 -7255 12060 -7221
rect 12015 -7291 12022 -7255
rect 12056 -7291 12060 -7255
rect 12015 -7325 12060 -7291
rect 12015 -7361 12022 -7325
rect 12056 -7361 12060 -7325
rect 11877 -7445 11893 -7411
rect 11927 -7445 11943 -7411
rect 11877 -7553 11893 -7519
rect 11927 -7553 11943 -7519
rect 11758 -7639 11764 -7603
rect 11798 -7639 11803 -7603
rect 11758 -7673 11803 -7639
rect 11758 -7709 11764 -7673
rect 11798 -7709 11803 -7673
rect 11758 -7743 11803 -7709
rect 11758 -7779 11764 -7743
rect 11798 -7779 11803 -7743
rect 11619 -7863 11635 -7829
rect 11669 -7863 11685 -7829
rect 11758 -7897 11803 -7779
rect 12015 -7603 12060 -7361
rect 12274 -7185 12319 -6943
rect 12532 -6767 12577 -6525
rect 12532 -6803 12538 -6767
rect 12572 -6803 12577 -6767
rect 12532 -6837 12577 -6803
rect 12532 -6873 12538 -6837
rect 12572 -6873 12577 -6837
rect 12532 -6907 12577 -6873
rect 12532 -6943 12538 -6907
rect 12572 -6943 12577 -6907
rect 12393 -7027 12409 -6993
rect 12443 -7027 12459 -6993
rect 12393 -7135 12409 -7101
rect 12443 -7135 12459 -7101
rect 12274 -7221 12280 -7185
rect 12314 -7221 12319 -7185
rect 12274 -7255 12319 -7221
rect 12274 -7291 12280 -7255
rect 12314 -7291 12319 -7255
rect 12274 -7325 12319 -7291
rect 12274 -7361 12280 -7325
rect 12314 -7361 12319 -7325
rect 12135 -7445 12151 -7411
rect 12185 -7445 12201 -7411
rect 12135 -7553 12151 -7519
rect 12185 -7553 12201 -7519
rect 12015 -7639 12022 -7603
rect 12056 -7639 12060 -7603
rect 12015 -7673 12060 -7639
rect 12015 -7709 12022 -7673
rect 12056 -7709 12060 -7673
rect 12015 -7743 12060 -7709
rect 12015 -7779 12022 -7743
rect 12056 -7779 12060 -7743
rect 11877 -7863 11893 -7829
rect 11927 -7863 11943 -7829
rect 12015 -7897 12060 -7779
rect 12274 -7603 12319 -7361
rect 12532 -7185 12577 -6943
rect 12532 -7221 12538 -7185
rect 12572 -7221 12577 -7185
rect 12532 -7255 12577 -7221
rect 12532 -7291 12538 -7255
rect 12572 -7291 12577 -7255
rect 12532 -7325 12577 -7291
rect 12532 -7361 12538 -7325
rect 12572 -7361 12577 -7325
rect 12393 -7445 12409 -7411
rect 12443 -7445 12459 -7411
rect 12393 -7553 12409 -7519
rect 12443 -7553 12459 -7519
rect 12274 -7639 12280 -7603
rect 12314 -7639 12319 -7603
rect 12274 -7673 12319 -7639
rect 12274 -7709 12280 -7673
rect 12314 -7709 12319 -7673
rect 12274 -7743 12319 -7709
rect 12274 -7779 12280 -7743
rect 12314 -7779 12319 -7743
rect 12135 -7863 12151 -7829
rect 12185 -7863 12201 -7829
rect 12274 -7897 12319 -7779
rect 12532 -7603 12577 -7361
rect 12532 -7639 12538 -7603
rect 12572 -7639 12577 -7603
rect 12532 -7673 12577 -7639
rect 12532 -7709 12538 -7673
rect 12572 -7709 12577 -7673
rect 12532 -7743 12577 -7709
rect 12532 -7779 12538 -7743
rect 12572 -7779 12577 -7743
rect 12393 -7863 12409 -7829
rect 12443 -7863 12459 -7829
rect 12532 -7897 12577 -7779
rect 5135 -8117 6361 -8022
rect 7805 -8117 9031 -8022
rect 10468 -8116 11694 -8021
rect 5134 -8206 5150 -8172
rect 5184 -8206 5200 -8172
rect 5674 -8206 5690 -8172
rect 5724 -8206 5740 -8172
rect 6154 -8206 6165 -8172
rect 6215 -8206 6220 -8172
rect 4995 -8258 5057 -8236
rect 4995 -8292 5021 -8258
rect 5055 -8292 5057 -8258
rect 4995 -8326 5057 -8292
rect 4995 -8362 5021 -8326
rect 5055 -8362 5057 -8326
rect 4995 -8396 5057 -8362
rect 4995 -8430 5021 -8396
rect 5055 -8430 5057 -8396
rect 4995 -8472 5057 -8430
rect 5273 -8258 5341 -8238
rect 5273 -8292 5279 -8258
rect 5313 -8292 5341 -8258
rect 5273 -8326 5341 -8292
rect 5273 -8362 5279 -8326
rect 5313 -8362 5341 -8326
rect 5273 -8396 5341 -8362
rect 5273 -8430 5279 -8396
rect 5313 -8430 5341 -8396
rect 5273 -8474 5341 -8430
rect 5535 -8258 5597 -8236
rect 5535 -8292 5561 -8258
rect 5595 -8292 5597 -8258
rect 5535 -8326 5597 -8292
rect 5535 -8362 5561 -8326
rect 5595 -8362 5597 -8326
rect 5535 -8396 5597 -8362
rect 5535 -8430 5561 -8396
rect 5595 -8430 5597 -8396
rect 5535 -8472 5597 -8430
rect 5813 -8258 5881 -8238
rect 5813 -8292 5819 -8258
rect 5853 -8292 5881 -8258
rect 5813 -8326 5881 -8292
rect 5813 -8362 5819 -8326
rect 5853 -8362 5881 -8326
rect 5813 -8396 5881 -8362
rect 5813 -8430 5819 -8396
rect 5853 -8430 5881 -8396
rect 5813 -8474 5881 -8430
rect 6015 -8258 6077 -8236
rect 6015 -8292 6041 -8258
rect 6075 -8292 6077 -8258
rect 6015 -8326 6077 -8292
rect 6015 -8362 6041 -8326
rect 6075 -8362 6077 -8326
rect 6015 -8396 6077 -8362
rect 6015 -8430 6041 -8396
rect 6075 -8430 6077 -8396
rect 5134 -8516 5150 -8482
rect 5184 -8516 5200 -8482
rect 5674 -8516 5690 -8482
rect 5724 -8516 5740 -8482
rect 6015 -8601 6077 -8430
rect 6293 -8258 6361 -8117
rect 6657 -8204 6673 -8170
rect 6707 -8204 6723 -8170
rect 7167 -8194 7183 -8160
rect 7217 -8194 7233 -8160
rect 7804 -8206 7820 -8172
rect 7854 -8206 7870 -8172
rect 8344 -8206 8360 -8172
rect 8394 -8206 8410 -8172
rect 8824 -8206 8835 -8172
rect 8885 -8206 8890 -8172
rect 6293 -8292 6299 -8258
rect 6333 -8292 6361 -8258
rect 6293 -8326 6361 -8292
rect 6293 -8362 6299 -8326
rect 6333 -8362 6361 -8326
rect 6293 -8396 6361 -8362
rect 6293 -8430 6299 -8396
rect 6333 -8430 6361 -8396
rect 6293 -8474 6361 -8430
rect 6518 -8256 6580 -8234
rect 6518 -8290 6544 -8256
rect 6578 -8290 6580 -8256
rect 6518 -8324 6580 -8290
rect 6518 -8360 6544 -8324
rect 6578 -8360 6580 -8324
rect 6518 -8394 6580 -8360
rect 6518 -8428 6544 -8394
rect 6578 -8428 6580 -8394
rect 6518 -8470 6580 -8428
rect 6796 -8256 6864 -8236
rect 6796 -8290 6802 -8256
rect 6836 -8290 6864 -8256
rect 6796 -8324 6864 -8290
rect 6796 -8360 6802 -8324
rect 6836 -8360 6864 -8324
rect 6796 -8394 6864 -8360
rect 6796 -8428 6802 -8394
rect 6836 -8428 6864 -8394
rect 6796 -8472 6864 -8428
rect 7028 -8246 7090 -8224
rect 7028 -8280 7054 -8246
rect 7088 -8280 7090 -8246
rect 7028 -8314 7090 -8280
rect 7028 -8350 7054 -8314
rect 7088 -8350 7090 -8314
rect 7028 -8384 7090 -8350
rect 7028 -8418 7054 -8384
rect 7088 -8418 7090 -8384
rect 7028 -8460 7090 -8418
rect 7306 -8246 7374 -8226
rect 7306 -8280 7312 -8246
rect 7346 -8280 7374 -8246
rect 7306 -8314 7374 -8280
rect 7306 -8350 7312 -8314
rect 7346 -8350 7374 -8314
rect 7306 -8384 7374 -8350
rect 7306 -8418 7312 -8384
rect 7346 -8418 7374 -8384
rect 7306 -8462 7374 -8418
rect 7665 -8258 7727 -8236
rect 7665 -8292 7691 -8258
rect 7725 -8292 7727 -8258
rect 7665 -8326 7727 -8292
rect 7665 -8362 7691 -8326
rect 7725 -8362 7727 -8326
rect 7665 -8396 7727 -8362
rect 7665 -8430 7691 -8396
rect 7725 -8430 7727 -8396
rect 6154 -8516 6166 -8482
rect 6206 -8516 6220 -8482
rect 6657 -8514 6673 -8480
rect 6707 -8514 6723 -8480
rect 7167 -8504 7183 -8470
rect 7217 -8504 7233 -8470
rect 7665 -8472 7727 -8430
rect 7943 -8258 8011 -8238
rect 7943 -8292 7949 -8258
rect 7983 -8292 8011 -8258
rect 7943 -8326 8011 -8292
rect 7943 -8362 7949 -8326
rect 7983 -8362 8011 -8326
rect 7943 -8396 8011 -8362
rect 7943 -8430 7949 -8396
rect 7983 -8430 8011 -8396
rect 7943 -8474 8011 -8430
rect 8205 -8258 8267 -8236
rect 8205 -8292 8231 -8258
rect 8265 -8292 8267 -8258
rect 8205 -8326 8267 -8292
rect 8205 -8362 8231 -8326
rect 8265 -8362 8267 -8326
rect 8205 -8396 8267 -8362
rect 8205 -8430 8231 -8396
rect 8265 -8430 8267 -8396
rect 8205 -8472 8267 -8430
rect 8483 -8258 8551 -8238
rect 8483 -8292 8489 -8258
rect 8523 -8292 8551 -8258
rect 8483 -8326 8551 -8292
rect 8483 -8362 8489 -8326
rect 8523 -8362 8551 -8326
rect 8483 -8396 8551 -8362
rect 8483 -8430 8489 -8396
rect 8523 -8430 8551 -8396
rect 8483 -8474 8551 -8430
rect 8685 -8258 8747 -8236
rect 8685 -8292 8711 -8258
rect 8745 -8292 8747 -8258
rect 8685 -8326 8747 -8292
rect 8685 -8362 8711 -8326
rect 8745 -8362 8747 -8326
rect 8685 -8396 8747 -8362
rect 8685 -8430 8711 -8396
rect 8745 -8430 8747 -8396
rect 7804 -8516 7820 -8482
rect 7854 -8516 7870 -8482
rect 8344 -8516 8360 -8482
rect 8394 -8516 8410 -8482
rect 8685 -8542 8747 -8430
rect 8963 -8258 9031 -8117
rect 9327 -8204 9343 -8170
rect 9377 -8204 9393 -8170
rect 9837 -8194 9853 -8160
rect 9887 -8194 9903 -8160
rect 10467 -8205 10483 -8171
rect 10517 -8205 10533 -8171
rect 11007 -8205 11023 -8171
rect 11057 -8205 11073 -8171
rect 11487 -8205 11498 -8171
rect 11548 -8205 11553 -8171
rect 8963 -8292 8969 -8258
rect 9003 -8292 9031 -8258
rect 8963 -8326 9031 -8292
rect 8963 -8362 8969 -8326
rect 9003 -8362 9031 -8326
rect 8963 -8396 9031 -8362
rect 8963 -8430 8969 -8396
rect 9003 -8430 9031 -8396
rect 8963 -8474 9031 -8430
rect 9188 -8256 9250 -8234
rect 9188 -8290 9214 -8256
rect 9248 -8290 9250 -8256
rect 9188 -8324 9250 -8290
rect 9188 -8360 9214 -8324
rect 9248 -8360 9250 -8324
rect 9188 -8394 9250 -8360
rect 9188 -8428 9214 -8394
rect 9248 -8428 9250 -8394
rect 9188 -8470 9250 -8428
rect 9466 -8256 9534 -8236
rect 9466 -8290 9472 -8256
rect 9506 -8290 9534 -8256
rect 9466 -8324 9534 -8290
rect 9466 -8360 9472 -8324
rect 9506 -8360 9534 -8324
rect 9466 -8394 9534 -8360
rect 9466 -8428 9472 -8394
rect 9506 -8428 9534 -8394
rect 9466 -8472 9534 -8428
rect 9698 -8246 9760 -8224
rect 9698 -8280 9724 -8246
rect 9758 -8280 9760 -8246
rect 9698 -8314 9760 -8280
rect 9698 -8350 9724 -8314
rect 9758 -8350 9760 -8314
rect 9698 -8384 9760 -8350
rect 9698 -8418 9724 -8384
rect 9758 -8418 9760 -8384
rect 9698 -8460 9760 -8418
rect 9976 -8246 10044 -8226
rect 9976 -8280 9982 -8246
rect 10016 -8280 10044 -8246
rect 9976 -8314 10044 -8280
rect 9976 -8350 9982 -8314
rect 10016 -8350 10044 -8314
rect 9976 -8384 10044 -8350
rect 9976 -8418 9982 -8384
rect 10016 -8418 10044 -8384
rect 9976 -8462 10044 -8418
rect 10328 -8257 10390 -8235
rect 10328 -8291 10354 -8257
rect 10388 -8291 10390 -8257
rect 10328 -8325 10390 -8291
rect 10328 -8361 10354 -8325
rect 10388 -8361 10390 -8325
rect 10328 -8395 10390 -8361
rect 10328 -8429 10354 -8395
rect 10388 -8429 10390 -8395
rect 8824 -8516 8836 -8482
rect 8880 -8516 8890 -8482
rect 9327 -8514 9343 -8480
rect 9377 -8514 9393 -8480
rect 9837 -8504 9853 -8470
rect 9887 -8504 9903 -8470
rect 10328 -8471 10390 -8429
rect 10606 -8257 10674 -8237
rect 10606 -8291 10612 -8257
rect 10646 -8291 10674 -8257
rect 10606 -8325 10674 -8291
rect 10606 -8361 10612 -8325
rect 10646 -8361 10674 -8325
rect 10606 -8395 10674 -8361
rect 10606 -8429 10612 -8395
rect 10646 -8429 10674 -8395
rect 10606 -8473 10674 -8429
rect 10868 -8257 10930 -8235
rect 10868 -8291 10894 -8257
rect 10928 -8291 10930 -8257
rect 10868 -8325 10930 -8291
rect 10868 -8361 10894 -8325
rect 10928 -8361 10930 -8325
rect 10868 -8395 10930 -8361
rect 10868 -8429 10894 -8395
rect 10928 -8429 10930 -8395
rect 10868 -8471 10930 -8429
rect 11146 -8257 11214 -8237
rect 11146 -8291 11152 -8257
rect 11186 -8291 11214 -8257
rect 11146 -8325 11214 -8291
rect 11146 -8361 11152 -8325
rect 11186 -8361 11214 -8325
rect 11146 -8395 11214 -8361
rect 11146 -8429 11152 -8395
rect 11186 -8429 11214 -8395
rect 11146 -8473 11214 -8429
rect 11348 -8257 11410 -8235
rect 11348 -8291 11374 -8257
rect 11408 -8291 11410 -8257
rect 11348 -8325 11410 -8291
rect 11348 -8361 11374 -8325
rect 11408 -8361 11410 -8325
rect 11348 -8395 11410 -8361
rect 11348 -8429 11374 -8395
rect 11408 -8429 11410 -8395
rect 10467 -8515 10483 -8481
rect 10517 -8515 10533 -8481
rect 11007 -8515 11023 -8481
rect 11057 -8515 11073 -8481
rect 8684 -8601 8747 -8542
rect 11348 -8601 11410 -8429
rect 11626 -8257 11694 -8116
rect 11990 -8203 12006 -8169
rect 12040 -8203 12056 -8169
rect 12500 -8193 12516 -8159
rect 12550 -8193 12566 -8159
rect 11626 -8291 11632 -8257
rect 11666 -8291 11694 -8257
rect 11626 -8325 11694 -8291
rect 11626 -8361 11632 -8325
rect 11666 -8361 11694 -8325
rect 11626 -8395 11694 -8361
rect 11626 -8429 11632 -8395
rect 11666 -8429 11694 -8395
rect 11626 -8473 11694 -8429
rect 11851 -8255 11913 -8233
rect 11851 -8289 11877 -8255
rect 11911 -8289 11913 -8255
rect 11851 -8323 11913 -8289
rect 11851 -8359 11877 -8323
rect 11911 -8359 11913 -8323
rect 11851 -8393 11913 -8359
rect 11851 -8427 11877 -8393
rect 11911 -8427 11913 -8393
rect 11851 -8469 11913 -8427
rect 12129 -8255 12197 -8235
rect 12129 -8289 12135 -8255
rect 12169 -8289 12197 -8255
rect 12129 -8323 12197 -8289
rect 12129 -8359 12135 -8323
rect 12169 -8359 12197 -8323
rect 12129 -8393 12197 -8359
rect 12129 -8427 12135 -8393
rect 12169 -8427 12197 -8393
rect 12129 -8471 12197 -8427
rect 12361 -8245 12423 -8223
rect 12361 -8279 12387 -8245
rect 12421 -8279 12423 -8245
rect 12361 -8313 12423 -8279
rect 12361 -8349 12387 -8313
rect 12421 -8349 12423 -8313
rect 12361 -8383 12423 -8349
rect 12361 -8417 12387 -8383
rect 12421 -8417 12423 -8383
rect 12361 -8459 12423 -8417
rect 12639 -8245 12707 -8225
rect 12639 -8279 12645 -8245
rect 12679 -8279 12707 -8245
rect 12639 -8313 12707 -8279
rect 12639 -8349 12645 -8313
rect 12679 -8349 12707 -8313
rect 12639 -8383 12707 -8349
rect 12639 -8417 12645 -8383
rect 12679 -8417 12707 -8383
rect 12639 -8461 12707 -8417
rect 11487 -8515 11498 -8481
rect 11542 -8515 11553 -8481
rect 11990 -8513 12006 -8479
rect 12040 -8513 12056 -8479
rect 12500 -8503 12516 -8469
rect 12550 -8503 12566 -8469
rect 4851 -8608 12841 -8601
rect 4848 -8702 6000 -8608
rect 6092 -8702 8670 -8608
rect 8762 -8702 11336 -8608
rect 11428 -8702 12908 -8608
rect 4848 -8796 12908 -8702
rect 14124 8623 15448 8668
rect 14064 8589 14080 8623
rect 14018 8539 14052 8555
rect 14018 7147 14052 7163
rect 14124 7113 15448 8589
rect 15941 8623 17272 8668
rect 17306 8589 17322 8623
rect 14064 7079 14080 7113
rect 14018 7029 14052 7045
rect 14018 5637 14052 5653
rect 14124 5603 15448 7079
rect 14064 5569 14080 5603
rect 14018 5519 14052 5535
rect 14018 4127 14052 4143
rect 14124 4093 15448 5569
rect 14064 4059 14080 4093
rect 14018 4009 14052 4025
rect 14018 2617 14052 2633
rect 14124 2583 15448 4059
rect 14064 2549 14080 2583
rect 14018 2499 14052 2515
rect 14018 1107 14052 1123
rect 14124 1073 15448 2549
rect 14064 1039 14080 1073
rect 14018 989 14052 1005
rect 14018 -403 14052 -387
rect 14124 -437 15448 1039
rect 14064 -471 14080 -437
rect 14018 -521 14052 -505
rect 14018 -1913 14052 -1897
rect 14124 -1947 15448 -471
rect 14064 -1981 14080 -1947
rect 14018 -2031 14052 -2015
rect 14018 -3423 14052 -3407
rect 14124 -3457 15448 -1981
rect 14064 -3491 14080 -3457
rect 14018 -3541 14052 -3525
rect 14018 -4933 14052 -4917
rect 14124 -4967 15448 -3491
rect 14064 -5001 14080 -4967
rect 14018 -5051 14052 -5035
rect 14018 -6443 14052 -6427
rect 14124 -6477 15448 -5001
rect 14064 -6511 14080 -6477
rect 14018 -6561 14052 -6545
rect 14018 -7953 14052 -7937
rect 14124 -7987 15448 -6511
rect 14064 -8021 14080 -7987
rect 14018 -8071 14052 -8055
rect 14018 -9463 14052 -9447
rect 14124 -9497 15448 -8021
rect 14064 -9531 14080 -9497
rect 14124 -9547 15448 -9531
rect 15670 8539 15719 8556
rect 15670 7163 15676 8539
rect 15710 7163 15719 8539
rect 15670 7029 15719 7163
rect 15670 5653 15676 7029
rect 15710 5653 15719 7029
rect 15670 5519 15719 5653
rect 15670 4143 15676 5519
rect 15710 4143 15719 5519
rect 15670 4009 15719 4143
rect 15670 2633 15676 4009
rect 15710 2633 15719 4009
rect 15670 2499 15719 2633
rect 15670 1123 15676 2499
rect 15710 1123 15719 2499
rect 15670 989 15719 1123
rect 15670 -387 15676 989
rect 15710 -387 15719 989
rect 15670 -521 15719 -387
rect 15670 -1897 15676 -521
rect 15710 -1897 15719 -521
rect 15670 -2031 15719 -1897
rect 15670 -3407 15676 -2031
rect 15710 -3407 15719 -2031
rect 15670 -3541 15719 -3407
rect 15670 -4917 15676 -3541
rect 15710 -4917 15719 -3541
rect 15670 -5051 15719 -4917
rect 15670 -6427 15676 -5051
rect 15710 -6427 15719 -5051
rect 15670 -6561 15719 -6427
rect 15670 -7937 15676 -6561
rect 15710 -7937 15719 -6561
rect 15670 -8071 15719 -7937
rect 15670 -9447 15676 -8071
rect 15710 -9447 15719 -8071
rect 15670 -9547 15719 -9447
rect 15941 8503 17272 8589
rect 17334 8539 17368 8555
rect 15941 7113 17268 8503
rect 17334 7147 17368 7163
rect 17306 7079 17322 7113
rect 15941 5603 17268 7079
rect 17334 7029 17368 7045
rect 17334 5637 17368 5653
rect 17306 5569 17322 5603
rect 15941 4093 17268 5569
rect 17334 5519 17368 5535
rect 17334 4127 17368 4143
rect 17306 4059 17322 4093
rect 15941 2583 17268 4059
rect 17334 4009 17368 4025
rect 17334 2617 17368 2633
rect 17306 2549 17322 2583
rect 15941 1073 17268 2549
rect 17334 2499 17368 2515
rect 17334 1107 17368 1123
rect 17306 1039 17322 1073
rect 15941 -437 17268 1039
rect 17334 989 17368 1005
rect 17334 -403 17368 -387
rect 17306 -471 17322 -437
rect 15941 -1947 17268 -471
rect 17334 -521 17368 -505
rect 17334 -1913 17368 -1897
rect 17306 -1981 17322 -1947
rect 15941 -3457 17268 -1981
rect 17334 -2031 17368 -2015
rect 17334 -3423 17368 -3407
rect 17306 -3491 17322 -3457
rect 15941 -4967 17268 -3491
rect 17334 -3541 17368 -3525
rect 17334 -4933 17368 -4917
rect 17306 -5001 17322 -4967
rect 15941 -6477 17268 -5001
rect 17334 -5051 17368 -5035
rect 17334 -6443 17368 -6427
rect 17306 -6511 17322 -6477
rect 15941 -7987 17268 -6511
rect 17334 -6561 17368 -6545
rect 17334 -7953 17368 -7937
rect 17306 -8021 17322 -7987
rect 15941 -9497 17268 -8021
rect 17334 -8071 17368 -8055
rect 17334 -9463 17368 -9447
rect 17306 -9531 17322 -9497
rect 15941 -9547 17268 -9531
<< viali >>
rect 282 8628 318 8655
rect 282 -9538 283 8628
rect 283 -9538 317 8628
rect 317 -9538 318 8628
rect 397 7162 431 8538
rect 3826 8628 3862 8654
rect 397 5652 431 7028
rect 397 4142 431 5518
rect 397 2632 431 4008
rect 397 1122 431 2498
rect 397 -388 431 988
rect 397 -1898 431 -522
rect 397 -3408 431 -2032
rect 397 -4918 431 -3542
rect 397 -6428 431 -5052
rect 397 -7938 431 -6562
rect 397 -9448 431 -8072
rect 282 -9598 318 -9538
rect 2055 7162 2089 8538
rect 2055 5652 2089 7028
rect 2055 4142 2089 5518
rect 2055 2632 2089 4008
rect 2055 1122 2089 2498
rect 2055 -388 2089 988
rect 2055 -1898 2089 -522
rect 2055 -3408 2089 -2032
rect 2055 -4918 2089 -3542
rect 2055 -6428 2089 -5052
rect 2055 -7938 2089 -6562
rect 2055 -9448 2089 -8072
rect 3713 7162 3747 8538
rect 3713 5652 3747 7028
rect 3713 4142 3747 5518
rect 3713 2632 3747 4008
rect 3713 1122 3747 2498
rect 3713 -388 3747 988
rect 3713 -1898 3747 -522
rect 3713 -3408 3747 -2032
rect 3713 -4918 3747 -3542
rect 3713 -6428 3747 -5052
rect 3713 -7938 3747 -6562
rect 3713 -9448 3747 -8072
rect 3826 -9538 3827 8628
rect 3827 -9538 3861 8628
rect 3861 -9538 3862 8628
rect 6204 8545 6238 8579
rect 6204 8217 6238 8251
rect 9092 8544 9126 8578
rect 9350 8544 9384 8578
rect 9092 8216 9126 8250
rect 9608 8544 9642 8578
rect 9866 8544 9900 8578
rect 10124 8544 10158 8578
rect 9350 8216 9384 8250
rect 9608 8216 9642 8250
rect 9866 8216 9900 8250
rect 10124 8216 10158 8250
rect 5064 7498 5237 7516
rect 5064 7236 5083 7498
rect 5083 7236 5220 7498
rect 5220 7236 5237 7498
rect 6121 7605 6201 7606
rect 6121 7571 6201 7605
rect 6121 7545 6201 7571
rect 6122 7367 6202 7385
rect 6122 7333 6202 7367
rect 6122 7324 6202 7333
rect 5064 7214 5237 7236
rect 8795 7571 8893 7602
rect 8795 7519 8893 7571
rect 8795 7367 8893 7407
rect 8795 7333 8893 7367
rect 8795 7324 8893 7333
rect 13903 8629 13938 8655
rect 11447 7572 11545 7602
rect 11447 7519 11545 7572
rect 11447 7368 11545 7407
rect 11447 7334 11545 7368
rect 11447 7324 11545 7334
rect 12464 7479 12679 7503
rect 8783 6728 8878 6807
rect 11456 6728 11551 6807
rect 12464 7217 12502 7479
rect 12502 7217 12639 7479
rect 12639 7217 12679 7479
rect 12464 7184 12679 7217
rect 12692 6742 12860 6920
rect 5270 6575 5304 6609
rect 5528 6575 5562 6609
rect 5786 6575 5820 6609
rect 6044 6575 6078 6609
rect 6302 6575 6336 6609
rect 6560 6575 6594 6609
rect 6818 6575 6852 6609
rect 7076 6575 7110 6609
rect 5270 6265 5304 6299
rect 5270 6157 5304 6191
rect 5528 6265 5562 6299
rect 5528 6157 5562 6191
rect 5270 5847 5304 5881
rect 5270 5739 5304 5773
rect 5786 6265 5820 6299
rect 5786 6157 5820 6191
rect 5528 5847 5562 5881
rect 5528 5739 5562 5773
rect 5270 5429 5304 5463
rect 5270 5321 5304 5355
rect 6044 6265 6078 6299
rect 6044 6157 6078 6191
rect 5786 5847 5820 5881
rect 5786 5739 5820 5773
rect 5528 5429 5562 5463
rect 5528 5321 5562 5355
rect 5270 5011 5304 5045
rect 5270 4903 5304 4937
rect 6302 6265 6336 6299
rect 6302 6157 6336 6191
rect 6044 5847 6078 5881
rect 6044 5739 6078 5773
rect 5786 5429 5820 5463
rect 5786 5321 5820 5355
rect 5528 5011 5562 5045
rect 5528 4903 5562 4937
rect 5270 4593 5304 4627
rect 5270 4485 5304 4519
rect 6560 6265 6594 6299
rect 6560 6157 6594 6191
rect 6302 5847 6336 5881
rect 6302 5739 6336 5773
rect 6044 5429 6078 5463
rect 6044 5321 6078 5355
rect 5786 5011 5820 5045
rect 5786 4903 5820 4937
rect 5528 4593 5562 4627
rect 5528 4485 5562 4519
rect 5270 4175 5304 4209
rect 5270 4067 5304 4101
rect 6818 6265 6852 6299
rect 6818 6157 6852 6191
rect 6560 5847 6594 5881
rect 6560 5739 6594 5773
rect 6302 5429 6336 5463
rect 6302 5321 6336 5355
rect 6044 5011 6078 5045
rect 6044 4903 6078 4937
rect 5786 4593 5820 4627
rect 5786 4485 5820 4519
rect 5528 4175 5562 4209
rect 5528 4067 5562 4101
rect 5270 3757 5304 3791
rect 7940 6575 7974 6609
rect 8198 6575 8232 6609
rect 8456 6575 8490 6609
rect 8714 6575 8748 6609
rect 8972 6575 9006 6609
rect 9230 6575 9264 6609
rect 9488 6575 9522 6609
rect 9746 6575 9780 6609
rect 7076 6265 7110 6299
rect 7076 6157 7110 6191
rect 6818 5847 6852 5881
rect 6818 5739 6852 5773
rect 6560 5429 6594 5463
rect 6560 5321 6594 5355
rect 6302 5011 6336 5045
rect 6302 4903 6336 4937
rect 6044 4593 6078 4627
rect 6044 4485 6078 4519
rect 5786 4175 5820 4209
rect 5786 4067 5820 4101
rect 5528 3757 5562 3791
rect 7076 5847 7110 5881
rect 7076 5739 7110 5773
rect 6818 5429 6852 5463
rect 6818 5321 6852 5355
rect 6560 5011 6594 5045
rect 6560 4903 6594 4937
rect 6302 4593 6336 4627
rect 6302 4485 6336 4519
rect 6044 4175 6078 4209
rect 6044 4067 6078 4101
rect 5786 3757 5820 3791
rect 7076 5429 7110 5463
rect 7076 5321 7110 5355
rect 6818 5011 6852 5045
rect 6818 4903 6852 4937
rect 6560 4593 6594 4627
rect 6560 4485 6594 4519
rect 6302 4175 6336 4209
rect 6302 4067 6336 4101
rect 6044 3757 6078 3791
rect 7076 5011 7110 5045
rect 7076 4903 7110 4937
rect 6818 4593 6852 4627
rect 6818 4485 6852 4519
rect 6560 4175 6594 4209
rect 6560 4067 6594 4101
rect 6302 3757 6336 3791
rect 7076 4593 7110 4627
rect 7076 4485 7110 4519
rect 6818 4175 6852 4209
rect 6818 4067 6852 4101
rect 6560 3757 6594 3791
rect 7076 4175 7110 4209
rect 7076 4067 7110 4101
rect 6818 3757 6852 3791
rect 7076 3757 7110 3791
rect 7940 6265 7974 6299
rect 7940 6157 7974 6191
rect 8198 6265 8232 6299
rect 8198 6157 8232 6191
rect 7940 5847 7974 5881
rect 7940 5739 7974 5773
rect 8456 6265 8490 6299
rect 8456 6157 8490 6191
rect 8198 5847 8232 5881
rect 8198 5739 8232 5773
rect 7940 5429 7974 5463
rect 7940 5321 7974 5355
rect 8714 6265 8748 6299
rect 8714 6157 8748 6191
rect 8456 5847 8490 5881
rect 8456 5739 8490 5773
rect 8198 5429 8232 5463
rect 8198 5321 8232 5355
rect 7940 5011 7974 5045
rect 7940 4903 7974 4937
rect 8972 6265 9006 6299
rect 8972 6157 9006 6191
rect 8714 5847 8748 5881
rect 8714 5739 8748 5773
rect 8456 5429 8490 5463
rect 8456 5321 8490 5355
rect 8198 5011 8232 5045
rect 8198 4903 8232 4937
rect 7940 4593 7974 4627
rect 7940 4485 7974 4519
rect 9230 6265 9264 6299
rect 9230 6157 9264 6191
rect 8972 5847 9006 5881
rect 8972 5739 9006 5773
rect 8714 5429 8748 5463
rect 8714 5321 8748 5355
rect 8456 5011 8490 5045
rect 8456 4903 8490 4937
rect 8198 4593 8232 4627
rect 8198 4485 8232 4519
rect 7940 4175 7974 4209
rect 7940 4067 7974 4101
rect 9488 6265 9522 6299
rect 9488 6157 9522 6191
rect 9230 5847 9264 5881
rect 9230 5739 9264 5773
rect 8972 5429 9006 5463
rect 8972 5321 9006 5355
rect 8714 5011 8748 5045
rect 8714 4903 8748 4937
rect 8456 4593 8490 4627
rect 8456 4485 8490 4519
rect 8198 4175 8232 4209
rect 8198 4067 8232 4101
rect 7940 3757 7974 3791
rect 10603 6576 10637 6610
rect 10861 6576 10895 6610
rect 11119 6576 11153 6610
rect 11377 6576 11411 6610
rect 11635 6576 11669 6610
rect 11893 6576 11927 6610
rect 12151 6576 12185 6610
rect 12409 6576 12443 6610
rect 9746 6265 9780 6299
rect 9746 6157 9780 6191
rect 9488 5847 9522 5881
rect 9488 5739 9522 5773
rect 9230 5429 9264 5463
rect 9230 5321 9264 5355
rect 8972 5011 9006 5045
rect 8972 4903 9006 4937
rect 8714 4593 8748 4627
rect 8714 4485 8748 4519
rect 8456 4175 8490 4209
rect 8456 4067 8490 4101
rect 8198 3757 8232 3791
rect 9746 5847 9780 5881
rect 9746 5739 9780 5773
rect 9488 5429 9522 5463
rect 9488 5321 9522 5355
rect 9230 5011 9264 5045
rect 9230 4903 9264 4937
rect 8972 4593 9006 4627
rect 8972 4485 9006 4519
rect 8714 4175 8748 4209
rect 8714 4067 8748 4101
rect 8456 3757 8490 3791
rect 9746 5429 9780 5463
rect 9746 5321 9780 5355
rect 9488 5011 9522 5045
rect 9488 4903 9522 4937
rect 9230 4593 9264 4627
rect 9230 4485 9264 4519
rect 8972 4175 9006 4209
rect 8972 4067 9006 4101
rect 8714 3757 8748 3791
rect 9746 5011 9780 5045
rect 9746 4903 9780 4937
rect 9488 4593 9522 4627
rect 9488 4485 9522 4519
rect 9230 4175 9264 4209
rect 9230 4067 9264 4101
rect 8972 3757 9006 3791
rect 9746 4593 9780 4627
rect 9746 4485 9780 4519
rect 9488 4175 9522 4209
rect 9488 4067 9522 4101
rect 9230 3757 9264 3791
rect 9746 4175 9780 4209
rect 9746 4067 9780 4101
rect 9488 3757 9522 3791
rect 9746 3757 9780 3791
rect 10603 6266 10637 6300
rect 10603 6158 10637 6192
rect 10861 6266 10895 6300
rect 10861 6158 10895 6192
rect 10603 5848 10637 5882
rect 10603 5740 10637 5774
rect 11119 6266 11153 6300
rect 11119 6158 11153 6192
rect 10861 5848 10895 5882
rect 10861 5740 10895 5774
rect 10603 5430 10637 5464
rect 10603 5322 10637 5356
rect 11377 6266 11411 6300
rect 11377 6158 11411 6192
rect 11119 5848 11153 5882
rect 11119 5740 11153 5774
rect 10861 5430 10895 5464
rect 10861 5322 10895 5356
rect 10603 5012 10637 5046
rect 10603 4904 10637 4938
rect 11635 6266 11669 6300
rect 11635 6158 11669 6192
rect 11377 5848 11411 5882
rect 11377 5740 11411 5774
rect 11119 5430 11153 5464
rect 11119 5322 11153 5356
rect 10861 5012 10895 5046
rect 10861 4904 10895 4938
rect 10603 4594 10637 4628
rect 10603 4486 10637 4520
rect 11893 6266 11927 6300
rect 11893 6158 11927 6192
rect 11635 5848 11669 5882
rect 11635 5740 11669 5774
rect 11377 5430 11411 5464
rect 11377 5322 11411 5356
rect 11119 5012 11153 5046
rect 11119 4904 11153 4938
rect 10861 4594 10895 4628
rect 10861 4486 10895 4520
rect 10603 4176 10637 4210
rect 10603 4068 10637 4102
rect 12151 6266 12185 6300
rect 12151 6158 12185 6192
rect 11893 5848 11927 5882
rect 11893 5740 11927 5774
rect 11635 5430 11669 5464
rect 11635 5322 11669 5356
rect 11377 5012 11411 5046
rect 11377 4904 11411 4938
rect 11119 4594 11153 4628
rect 11119 4486 11153 4520
rect 10861 4176 10895 4210
rect 10861 4068 10895 4102
rect 10603 3758 10637 3792
rect 12409 6266 12443 6300
rect 12409 6158 12443 6192
rect 12151 5848 12185 5882
rect 12151 5740 12185 5774
rect 11893 5430 11927 5464
rect 11893 5322 11927 5356
rect 11635 5012 11669 5046
rect 11635 4904 11669 4938
rect 11377 4594 11411 4628
rect 11377 4486 11411 4520
rect 11119 4176 11153 4210
rect 11119 4068 11153 4102
rect 10861 3758 10895 3792
rect 12409 5848 12443 5882
rect 12409 5740 12443 5774
rect 12151 5430 12185 5464
rect 12151 5322 12185 5356
rect 11893 5012 11927 5046
rect 11893 4904 11927 4938
rect 11635 4594 11669 4628
rect 11635 4486 11669 4520
rect 11377 4176 11411 4210
rect 11377 4068 11411 4102
rect 11119 3758 11153 3792
rect 12409 5430 12443 5464
rect 12409 5322 12443 5356
rect 12151 5012 12185 5046
rect 12151 4904 12185 4938
rect 11893 4594 11927 4628
rect 11893 4486 11927 4520
rect 11635 4176 11669 4210
rect 11635 4068 11669 4102
rect 11377 3758 11411 3792
rect 12409 5012 12443 5046
rect 12409 4904 12443 4938
rect 12151 4594 12185 4628
rect 12151 4486 12185 4520
rect 11893 4176 11927 4210
rect 11893 4068 11927 4102
rect 11635 3758 11669 3792
rect 12409 4594 12443 4628
rect 12409 4486 12443 4520
rect 12151 4176 12185 4210
rect 12151 4068 12185 4102
rect 11893 3758 11927 3792
rect 12409 4176 12443 4210
rect 12409 4068 12443 4102
rect 12151 3758 12185 3792
rect 12409 3758 12443 3792
rect 6165 3415 6170 3449
rect 6170 3415 6204 3449
rect 6204 3415 6215 3449
rect 6165 3409 6215 3415
rect 8835 3415 8840 3449
rect 8840 3415 8874 3449
rect 8874 3415 8885 3449
rect 8835 3409 8885 3415
rect 6168 3139 6206 3142
rect 6168 3105 6170 3139
rect 6170 3105 6204 3139
rect 6204 3105 6206 3139
rect 6168 3102 6206 3105
rect 11498 3416 11503 3450
rect 11503 3416 11537 3450
rect 11537 3416 11548 3450
rect 11498 3410 11548 3416
rect 8838 3139 8876 3142
rect 8838 3105 8840 3139
rect 8840 3105 8874 3139
rect 8874 3105 8876 3139
rect 8838 3102 8876 3105
rect 11500 3140 11538 3142
rect 11500 3106 11503 3140
rect 11503 3106 11537 3140
rect 11537 3106 11538 3140
rect 11500 3102 11538 3106
rect 5998 2906 6104 3012
rect 8662 2906 8768 3012
rect 11324 2906 11430 3012
rect 5019 1932 5202 1953
rect 5019 1670 5042 1932
rect 5042 1670 5179 1932
rect 5179 1670 5202 1932
rect 6121 1923 6201 1924
rect 6121 1889 6201 1923
rect 6121 1863 6201 1889
rect 6120 1685 6200 1703
rect 5019 1648 5202 1670
rect 6120 1651 6200 1685
rect 6120 1642 6200 1651
rect 8776 1889 8874 1920
rect 8776 1837 8874 1889
rect 11451 1890 11549 1920
rect 11451 1837 11549 1890
rect 8776 1685 8874 1725
rect 8776 1651 8874 1685
rect 8776 1642 8874 1651
rect 4884 1002 5042 1166
rect 11451 1686 11549 1725
rect 11451 1652 11549 1686
rect 11451 1642 11549 1652
rect 7590 982 7708 1116
rect 5270 858 5304 892
rect 5528 858 5562 892
rect 5786 858 5820 892
rect 6044 858 6078 892
rect 6302 858 6336 892
rect 6560 858 6594 892
rect 6818 858 6852 892
rect 7076 858 7110 892
rect 5270 548 5304 582
rect 5270 440 5304 474
rect 5528 548 5562 582
rect 5528 440 5562 474
rect 5270 130 5304 164
rect 5270 22 5304 56
rect 5786 548 5820 582
rect 5786 440 5820 474
rect 5528 130 5562 164
rect 5528 22 5562 56
rect 5270 -288 5304 -254
rect 5270 -396 5304 -362
rect 6044 548 6078 582
rect 6044 440 6078 474
rect 5786 130 5820 164
rect 5786 22 5820 56
rect 5528 -288 5562 -254
rect 5528 -396 5562 -362
rect 5270 -706 5304 -672
rect 5270 -814 5304 -780
rect 6302 548 6336 582
rect 6302 440 6336 474
rect 6044 130 6078 164
rect 6044 22 6078 56
rect 5786 -288 5820 -254
rect 5786 -396 5820 -362
rect 5528 -706 5562 -672
rect 5528 -814 5562 -780
rect 5270 -1124 5304 -1090
rect 5270 -1232 5304 -1198
rect 6560 548 6594 582
rect 6560 440 6594 474
rect 6302 130 6336 164
rect 6302 22 6336 56
rect 6044 -288 6078 -254
rect 6044 -396 6078 -362
rect 5786 -706 5820 -672
rect 5786 -814 5820 -780
rect 5528 -1124 5562 -1090
rect 5528 -1232 5562 -1198
rect 5270 -1542 5304 -1508
rect 5270 -1650 5304 -1616
rect 10196 982 10308 1106
rect 7940 858 7974 892
rect 8198 858 8232 892
rect 8456 858 8490 892
rect 8714 858 8748 892
rect 8972 858 9006 892
rect 9230 858 9264 892
rect 9488 858 9522 892
rect 9746 858 9780 892
rect 6818 548 6852 582
rect 6818 440 6852 474
rect 6560 130 6594 164
rect 6560 22 6594 56
rect 6302 -288 6336 -254
rect 6302 -396 6336 -362
rect 6044 -706 6078 -672
rect 6044 -814 6078 -780
rect 5786 -1124 5820 -1090
rect 5786 -1232 5820 -1198
rect 5528 -1542 5562 -1508
rect 5528 -1650 5562 -1616
rect 5270 -1960 5304 -1926
rect 7076 548 7110 582
rect 7076 440 7110 474
rect 6818 130 6852 164
rect 6818 22 6852 56
rect 6560 -288 6594 -254
rect 6560 -396 6594 -362
rect 6302 -706 6336 -672
rect 6302 -814 6336 -780
rect 6044 -1124 6078 -1090
rect 6044 -1232 6078 -1198
rect 5786 -1542 5820 -1508
rect 5786 -1650 5820 -1616
rect 5528 -1960 5562 -1926
rect 7076 130 7110 164
rect 7076 22 7110 56
rect 6818 -288 6852 -254
rect 6818 -396 6852 -362
rect 6560 -706 6594 -672
rect 6560 -814 6594 -780
rect 6302 -1124 6336 -1090
rect 6302 -1232 6336 -1198
rect 6044 -1542 6078 -1508
rect 6044 -1650 6078 -1616
rect 5786 -1960 5820 -1926
rect 7076 -288 7110 -254
rect 7076 -396 7110 -362
rect 6818 -706 6852 -672
rect 6818 -814 6852 -780
rect 6560 -1124 6594 -1090
rect 6560 -1232 6594 -1198
rect 6302 -1542 6336 -1508
rect 6302 -1650 6336 -1616
rect 6044 -1960 6078 -1926
rect 7076 -706 7110 -672
rect 7076 -814 7110 -780
rect 6818 -1124 6852 -1090
rect 6818 -1232 6852 -1198
rect 6560 -1542 6594 -1508
rect 6560 -1650 6594 -1616
rect 6302 -1960 6336 -1926
rect 7076 -1124 7110 -1090
rect 7076 -1232 7110 -1198
rect 6818 -1542 6852 -1508
rect 6818 -1650 6852 -1616
rect 6560 -1960 6594 -1926
rect 7076 -1542 7110 -1508
rect 7076 -1650 7110 -1616
rect 6818 -1960 6852 -1926
rect 7940 548 7974 582
rect 7940 440 7974 474
rect 8198 548 8232 582
rect 8198 440 8232 474
rect 7940 130 7974 164
rect 7940 22 7974 56
rect 8456 548 8490 582
rect 8456 440 8490 474
rect 8198 130 8232 164
rect 8198 22 8232 56
rect 7940 -288 7974 -254
rect 7940 -396 7974 -362
rect 8714 548 8748 582
rect 8714 440 8748 474
rect 8456 130 8490 164
rect 8456 22 8490 56
rect 8198 -288 8232 -254
rect 8198 -396 8232 -362
rect 7940 -706 7974 -672
rect 7940 -814 7974 -780
rect 8972 548 9006 582
rect 8972 440 9006 474
rect 8714 130 8748 164
rect 8714 22 8748 56
rect 8456 -288 8490 -254
rect 8456 -396 8490 -362
rect 8198 -706 8232 -672
rect 8198 -814 8232 -780
rect 7940 -1124 7974 -1090
rect 7940 -1232 7974 -1198
rect 9230 548 9264 582
rect 9230 440 9264 474
rect 8972 130 9006 164
rect 8972 22 9006 56
rect 8714 -288 8748 -254
rect 8714 -396 8748 -362
rect 8456 -706 8490 -672
rect 8456 -814 8490 -780
rect 8198 -1124 8232 -1090
rect 8198 -1232 8232 -1198
rect 7940 -1542 7974 -1508
rect 7940 -1650 7974 -1616
rect 7076 -1960 7110 -1926
rect 10603 859 10637 893
rect 10861 859 10895 893
rect 11119 859 11153 893
rect 11377 859 11411 893
rect 11635 859 11669 893
rect 11893 859 11927 893
rect 12151 859 12185 893
rect 12409 859 12443 893
rect 9488 548 9522 582
rect 9488 440 9522 474
rect 9230 130 9264 164
rect 9230 22 9264 56
rect 8972 -288 9006 -254
rect 8972 -396 9006 -362
rect 8714 -706 8748 -672
rect 8714 -814 8748 -780
rect 8456 -1124 8490 -1090
rect 8456 -1232 8490 -1198
rect 8198 -1542 8232 -1508
rect 8198 -1650 8232 -1616
rect 7940 -1960 7974 -1926
rect 9746 548 9780 582
rect 9746 440 9780 474
rect 9488 130 9522 164
rect 9488 22 9522 56
rect 9230 -288 9264 -254
rect 9230 -396 9264 -362
rect 8972 -706 9006 -672
rect 8972 -814 9006 -780
rect 8714 -1124 8748 -1090
rect 8714 -1232 8748 -1198
rect 8456 -1542 8490 -1508
rect 8456 -1650 8490 -1616
rect 8198 -1960 8232 -1926
rect 9746 130 9780 164
rect 9746 22 9780 56
rect 9488 -288 9522 -254
rect 9488 -396 9522 -362
rect 9230 -706 9264 -672
rect 9230 -814 9264 -780
rect 8972 -1124 9006 -1090
rect 8972 -1232 9006 -1198
rect 8714 -1542 8748 -1508
rect 8714 -1650 8748 -1616
rect 8456 -1960 8490 -1926
rect 9746 -288 9780 -254
rect 9746 -396 9780 -362
rect 9488 -706 9522 -672
rect 9488 -814 9522 -780
rect 9230 -1124 9264 -1090
rect 9230 -1232 9264 -1198
rect 8972 -1542 9006 -1508
rect 8972 -1650 9006 -1616
rect 8714 -1960 8748 -1926
rect 9746 -706 9780 -672
rect 9746 -814 9780 -780
rect 9488 -1124 9522 -1090
rect 9488 -1232 9522 -1198
rect 9230 -1542 9264 -1508
rect 9230 -1650 9264 -1616
rect 8972 -1960 9006 -1926
rect 9746 -1124 9780 -1090
rect 9746 -1232 9780 -1198
rect 9488 -1542 9522 -1508
rect 9488 -1650 9522 -1616
rect 9230 -1960 9264 -1926
rect 9746 -1542 9780 -1508
rect 9746 -1650 9780 -1616
rect 9488 -1960 9522 -1926
rect 10603 549 10637 583
rect 10603 441 10637 475
rect 10861 549 10895 583
rect 10861 441 10895 475
rect 10603 131 10637 165
rect 10603 23 10637 57
rect 11119 549 11153 583
rect 11119 441 11153 475
rect 10861 131 10895 165
rect 10861 23 10895 57
rect 10603 -287 10637 -253
rect 10603 -395 10637 -361
rect 11377 549 11411 583
rect 11377 441 11411 475
rect 11119 131 11153 165
rect 11119 23 11153 57
rect 10861 -287 10895 -253
rect 10861 -395 10895 -361
rect 10603 -705 10637 -671
rect 10603 -813 10637 -779
rect 11635 549 11669 583
rect 11635 441 11669 475
rect 11377 131 11411 165
rect 11377 23 11411 57
rect 11119 -287 11153 -253
rect 11119 -395 11153 -361
rect 10861 -705 10895 -671
rect 10861 -813 10895 -779
rect 10603 -1123 10637 -1089
rect 10603 -1231 10637 -1197
rect 11893 549 11927 583
rect 11893 441 11927 475
rect 11635 131 11669 165
rect 11635 23 11669 57
rect 11377 -287 11411 -253
rect 11377 -395 11411 -361
rect 11119 -705 11153 -671
rect 11119 -813 11153 -779
rect 10861 -1123 10895 -1089
rect 10861 -1231 10895 -1197
rect 10603 -1541 10637 -1507
rect 10603 -1649 10637 -1615
rect 9746 -1960 9780 -1926
rect 12151 549 12185 583
rect 12151 441 12185 475
rect 11893 131 11927 165
rect 11893 23 11927 57
rect 11635 -287 11669 -253
rect 11635 -395 11669 -361
rect 11377 -705 11411 -671
rect 11377 -813 11411 -779
rect 11119 -1123 11153 -1089
rect 11119 -1231 11153 -1197
rect 10861 -1541 10895 -1507
rect 10861 -1649 10895 -1615
rect 10603 -1959 10637 -1925
rect 12409 549 12443 583
rect 12409 441 12443 475
rect 12151 131 12185 165
rect 12151 23 12185 57
rect 11893 -287 11927 -253
rect 11893 -395 11927 -361
rect 11635 -705 11669 -671
rect 11635 -813 11669 -779
rect 11377 -1123 11411 -1089
rect 11377 -1231 11411 -1197
rect 11119 -1541 11153 -1507
rect 11119 -1649 11153 -1615
rect 10861 -1959 10895 -1925
rect 12409 131 12443 165
rect 12409 23 12443 57
rect 12151 -287 12185 -253
rect 12151 -395 12185 -361
rect 11893 -705 11927 -671
rect 11893 -813 11927 -779
rect 11635 -1123 11669 -1089
rect 11635 -1231 11669 -1197
rect 11377 -1541 11411 -1507
rect 11377 -1649 11411 -1615
rect 11119 -1959 11153 -1925
rect 12409 -287 12443 -253
rect 12409 -395 12443 -361
rect 12151 -705 12185 -671
rect 12151 -813 12185 -779
rect 11893 -1123 11927 -1089
rect 11893 -1231 11927 -1197
rect 11635 -1541 11669 -1507
rect 11635 -1649 11669 -1615
rect 11377 -1959 11411 -1925
rect 12409 -705 12443 -671
rect 12409 -813 12443 -779
rect 12151 -1123 12185 -1089
rect 12151 -1231 12185 -1197
rect 11893 -1541 11927 -1507
rect 11893 -1649 11927 -1615
rect 11635 -1959 11669 -1925
rect 12409 -1123 12443 -1089
rect 12409 -1231 12443 -1197
rect 12151 -1541 12185 -1507
rect 12151 -1649 12185 -1615
rect 11893 -1959 11927 -1925
rect 12409 -1541 12443 -1507
rect 12409 -1649 12443 -1615
rect 12151 -1959 12185 -1925
rect 12409 -1959 12443 -1925
rect 6165 -2302 6170 -2268
rect 6170 -2302 6204 -2268
rect 6204 -2302 6215 -2268
rect 6165 -2308 6215 -2302
rect 8835 -2302 8840 -2268
rect 8840 -2302 8874 -2268
rect 8874 -2302 8885 -2268
rect 8835 -2308 8885 -2302
rect 6168 -2578 6208 -2576
rect 6168 -2612 6170 -2578
rect 6170 -2612 6204 -2578
rect 6204 -2612 6208 -2578
rect 6168 -2614 6208 -2612
rect 11498 -2301 11503 -2267
rect 11503 -2301 11537 -2267
rect 11537 -2301 11548 -2267
rect 11498 -2307 11548 -2301
rect 8838 -2578 8878 -2576
rect 8838 -2612 8840 -2578
rect 8840 -2612 8874 -2578
rect 8874 -2612 8878 -2578
rect 8838 -2614 8878 -2612
rect 11498 -2577 11540 -2574
rect 11498 -2611 11503 -2577
rect 11503 -2611 11537 -2577
rect 11537 -2611 11540 -2577
rect 11498 -2616 11540 -2611
rect 5992 -2712 6098 -2707
rect 5992 -2806 6000 -2712
rect 6000 -2806 6092 -2712
rect 6092 -2806 6098 -2712
rect 8668 -2806 8760 -2712
rect 11334 -2806 11426 -2712
rect 5992 -2813 6098 -2806
rect 4998 -3951 5141 -3950
rect 4998 -4212 5001 -3951
rect 5001 -4212 5137 -3951
rect 5137 -4212 5141 -3951
rect 4998 -4214 5141 -4212
rect 6121 -4002 6201 -4001
rect 6121 -4036 6201 -4002
rect 6121 -4062 6201 -4036
rect 6122 -4240 6202 -4222
rect 6122 -4274 6202 -4240
rect 6122 -4283 6202 -4274
rect 8795 -4036 8893 -4005
rect 8795 -4088 8893 -4036
rect 8795 -4240 8893 -4200
rect 8795 -4274 8893 -4240
rect 8795 -4283 8893 -4274
rect 12726 -3402 12760 -3368
rect 13116 -3404 13150 -3370
rect 12275 -3406 12477 -3404
rect 12275 -3719 12276 -3406
rect 12276 -3719 12477 -3406
rect 12915 -3578 12986 -3574
rect 12915 -3640 12928 -3578
rect 12928 -3640 12984 -3578
rect 12984 -3640 12986 -3578
rect 12915 -3646 12986 -3640
rect 12726 -3866 12760 -3832
rect 13116 -3868 13150 -3834
rect 11447 -4035 11545 -4005
rect 11447 -4088 11545 -4035
rect 12876 -4046 12930 -4008
rect 13264 -4054 13312 -4010
rect 11447 -4239 11545 -4200
rect 11447 -4273 11545 -4239
rect 11447 -4283 11545 -4273
rect 12730 -4198 12764 -4164
rect 13120 -4198 13154 -4164
rect 12551 -4314 12554 -4242
rect 12554 -4314 12598 -4242
rect 12598 -4314 12607 -4242
rect 12551 -4315 12607 -4314
rect 12943 -4314 12944 -4242
rect 12944 -4314 12988 -4242
rect 12988 -4314 12989 -4242
rect 12943 -4315 12989 -4314
rect 12730 -4392 12764 -4358
rect 13120 -4392 13154 -4358
rect 8783 -4893 8878 -4814
rect 11456 -4893 11551 -4814
rect 12570 -4858 12820 -4568
rect 13192 -4860 13442 -4570
rect 5270 -5046 5304 -5012
rect 5528 -5046 5562 -5012
rect 5786 -5046 5820 -5012
rect 6044 -5046 6078 -5012
rect 6302 -5046 6336 -5012
rect 6560 -5046 6594 -5012
rect 6818 -5046 6852 -5012
rect 7076 -5046 7110 -5012
rect 5270 -5356 5304 -5322
rect 5270 -5464 5304 -5430
rect 5528 -5356 5562 -5322
rect 5528 -5464 5562 -5430
rect 5270 -5774 5304 -5740
rect 5270 -5882 5304 -5848
rect 5786 -5356 5820 -5322
rect 5786 -5464 5820 -5430
rect 5528 -5774 5562 -5740
rect 5528 -5882 5562 -5848
rect 5270 -6192 5304 -6158
rect 5270 -6300 5304 -6266
rect 6044 -5356 6078 -5322
rect 6044 -5464 6078 -5430
rect 5786 -5774 5820 -5740
rect 5786 -5882 5820 -5848
rect 5528 -6192 5562 -6158
rect 5528 -6300 5562 -6266
rect 5270 -6610 5304 -6576
rect 5270 -6718 5304 -6684
rect 6302 -5356 6336 -5322
rect 6302 -5464 6336 -5430
rect 6044 -5774 6078 -5740
rect 6044 -5882 6078 -5848
rect 5786 -6192 5820 -6158
rect 5786 -6300 5820 -6266
rect 5528 -6610 5562 -6576
rect 5528 -6718 5562 -6684
rect 5270 -7028 5304 -6994
rect 5270 -7136 5304 -7102
rect 6560 -5356 6594 -5322
rect 6560 -5464 6594 -5430
rect 6302 -5774 6336 -5740
rect 6302 -5882 6336 -5848
rect 6044 -6192 6078 -6158
rect 6044 -6300 6078 -6266
rect 5786 -6610 5820 -6576
rect 5786 -6718 5820 -6684
rect 5528 -7028 5562 -6994
rect 5528 -7136 5562 -7102
rect 5270 -7446 5304 -7412
rect 5270 -7554 5304 -7520
rect 6818 -5356 6852 -5322
rect 6818 -5464 6852 -5430
rect 6560 -5774 6594 -5740
rect 6560 -5882 6594 -5848
rect 6302 -6192 6336 -6158
rect 6302 -6300 6336 -6266
rect 6044 -6610 6078 -6576
rect 6044 -6718 6078 -6684
rect 5786 -7028 5820 -6994
rect 5786 -7136 5820 -7102
rect 5528 -7446 5562 -7412
rect 5528 -7554 5562 -7520
rect 5270 -7864 5304 -7830
rect 7940 -5046 7974 -5012
rect 8198 -5046 8232 -5012
rect 8456 -5046 8490 -5012
rect 8714 -5046 8748 -5012
rect 8972 -5046 9006 -5012
rect 9230 -5046 9264 -5012
rect 9488 -5046 9522 -5012
rect 9746 -5046 9780 -5012
rect 7076 -5356 7110 -5322
rect 7076 -5464 7110 -5430
rect 6818 -5774 6852 -5740
rect 6818 -5882 6852 -5848
rect 6560 -6192 6594 -6158
rect 6560 -6300 6594 -6266
rect 6302 -6610 6336 -6576
rect 6302 -6718 6336 -6684
rect 6044 -7028 6078 -6994
rect 6044 -7136 6078 -7102
rect 5786 -7446 5820 -7412
rect 5786 -7554 5820 -7520
rect 5528 -7864 5562 -7830
rect 7076 -5774 7110 -5740
rect 7076 -5882 7110 -5848
rect 6818 -6192 6852 -6158
rect 6818 -6300 6852 -6266
rect 6560 -6610 6594 -6576
rect 6560 -6718 6594 -6684
rect 6302 -7028 6336 -6994
rect 6302 -7136 6336 -7102
rect 6044 -7446 6078 -7412
rect 6044 -7554 6078 -7520
rect 5786 -7864 5820 -7830
rect 7076 -6192 7110 -6158
rect 7076 -6300 7110 -6266
rect 6818 -6610 6852 -6576
rect 6818 -6718 6852 -6684
rect 6560 -7028 6594 -6994
rect 6560 -7136 6594 -7102
rect 6302 -7446 6336 -7412
rect 6302 -7554 6336 -7520
rect 6044 -7864 6078 -7830
rect 7076 -6610 7110 -6576
rect 7076 -6718 7110 -6684
rect 6818 -7028 6852 -6994
rect 6818 -7136 6852 -7102
rect 6560 -7446 6594 -7412
rect 6560 -7554 6594 -7520
rect 6302 -7864 6336 -7830
rect 7076 -7028 7110 -6994
rect 7076 -7136 7110 -7102
rect 6818 -7446 6852 -7412
rect 6818 -7554 6852 -7520
rect 6560 -7864 6594 -7830
rect 7076 -7446 7110 -7412
rect 7076 -7554 7110 -7520
rect 6818 -7864 6852 -7830
rect 7076 -7864 7110 -7830
rect 7940 -5356 7974 -5322
rect 7940 -5464 7974 -5430
rect 8198 -5356 8232 -5322
rect 8198 -5464 8232 -5430
rect 7940 -5774 7974 -5740
rect 7940 -5882 7974 -5848
rect 8456 -5356 8490 -5322
rect 8456 -5464 8490 -5430
rect 8198 -5774 8232 -5740
rect 8198 -5882 8232 -5848
rect 7940 -6192 7974 -6158
rect 7940 -6300 7974 -6266
rect 8714 -5356 8748 -5322
rect 8714 -5464 8748 -5430
rect 8456 -5774 8490 -5740
rect 8456 -5882 8490 -5848
rect 8198 -6192 8232 -6158
rect 8198 -6300 8232 -6266
rect 7940 -6610 7974 -6576
rect 7940 -6718 7974 -6684
rect 8972 -5356 9006 -5322
rect 8972 -5464 9006 -5430
rect 8714 -5774 8748 -5740
rect 8714 -5882 8748 -5848
rect 8456 -6192 8490 -6158
rect 8456 -6300 8490 -6266
rect 8198 -6610 8232 -6576
rect 8198 -6718 8232 -6684
rect 7940 -7028 7974 -6994
rect 7940 -7136 7974 -7102
rect 9230 -5356 9264 -5322
rect 9230 -5464 9264 -5430
rect 8972 -5774 9006 -5740
rect 8972 -5882 9006 -5848
rect 8714 -6192 8748 -6158
rect 8714 -6300 8748 -6266
rect 8456 -6610 8490 -6576
rect 8456 -6718 8490 -6684
rect 8198 -7028 8232 -6994
rect 8198 -7136 8232 -7102
rect 7940 -7446 7974 -7412
rect 7940 -7554 7974 -7520
rect 9488 -5356 9522 -5322
rect 9488 -5464 9522 -5430
rect 9230 -5774 9264 -5740
rect 9230 -5882 9264 -5848
rect 8972 -6192 9006 -6158
rect 8972 -6300 9006 -6266
rect 8714 -6610 8748 -6576
rect 8714 -6718 8748 -6684
rect 8456 -7028 8490 -6994
rect 8456 -7136 8490 -7102
rect 8198 -7446 8232 -7412
rect 8198 -7554 8232 -7520
rect 7940 -7864 7974 -7830
rect 10603 -5045 10637 -5011
rect 10861 -5045 10895 -5011
rect 11119 -5045 11153 -5011
rect 11377 -5045 11411 -5011
rect 11635 -5045 11669 -5011
rect 11893 -5045 11927 -5011
rect 12151 -5045 12185 -5011
rect 12409 -5045 12443 -5011
rect 9746 -5356 9780 -5322
rect 9746 -5464 9780 -5430
rect 9488 -5774 9522 -5740
rect 9488 -5882 9522 -5848
rect 9230 -6192 9264 -6158
rect 9230 -6300 9264 -6266
rect 8972 -6610 9006 -6576
rect 8972 -6718 9006 -6684
rect 8714 -7028 8748 -6994
rect 8714 -7136 8748 -7102
rect 8456 -7446 8490 -7412
rect 8456 -7554 8490 -7520
rect 8198 -7864 8232 -7830
rect 9746 -5774 9780 -5740
rect 9746 -5882 9780 -5848
rect 9488 -6192 9522 -6158
rect 9488 -6300 9522 -6266
rect 9230 -6610 9264 -6576
rect 9230 -6718 9264 -6684
rect 8972 -7028 9006 -6994
rect 8972 -7136 9006 -7102
rect 8714 -7446 8748 -7412
rect 8714 -7554 8748 -7520
rect 8456 -7864 8490 -7830
rect 9746 -6192 9780 -6158
rect 9746 -6300 9780 -6266
rect 9488 -6610 9522 -6576
rect 9488 -6718 9522 -6684
rect 9230 -7028 9264 -6994
rect 9230 -7136 9264 -7102
rect 8972 -7446 9006 -7412
rect 8972 -7554 9006 -7520
rect 8714 -7864 8748 -7830
rect 9746 -6610 9780 -6576
rect 9746 -6718 9780 -6684
rect 9488 -7028 9522 -6994
rect 9488 -7136 9522 -7102
rect 9230 -7446 9264 -7412
rect 9230 -7554 9264 -7520
rect 8972 -7864 9006 -7830
rect 9746 -7028 9780 -6994
rect 9746 -7136 9780 -7102
rect 9488 -7446 9522 -7412
rect 9488 -7554 9522 -7520
rect 9230 -7864 9264 -7830
rect 9746 -7446 9780 -7412
rect 9746 -7554 9780 -7520
rect 9488 -7864 9522 -7830
rect 9746 -7864 9780 -7830
rect 10603 -5355 10637 -5321
rect 10603 -5463 10637 -5429
rect 10861 -5355 10895 -5321
rect 10861 -5463 10895 -5429
rect 10603 -5773 10637 -5739
rect 10603 -5881 10637 -5847
rect 11119 -5355 11153 -5321
rect 11119 -5463 11153 -5429
rect 10861 -5773 10895 -5739
rect 10861 -5881 10895 -5847
rect 10603 -6191 10637 -6157
rect 10603 -6299 10637 -6265
rect 11377 -5355 11411 -5321
rect 11377 -5463 11411 -5429
rect 11119 -5773 11153 -5739
rect 11119 -5881 11153 -5847
rect 10861 -6191 10895 -6157
rect 10861 -6299 10895 -6265
rect 10603 -6609 10637 -6575
rect 10603 -6717 10637 -6683
rect 11635 -5355 11669 -5321
rect 11635 -5463 11669 -5429
rect 11377 -5773 11411 -5739
rect 11377 -5881 11411 -5847
rect 11119 -6191 11153 -6157
rect 11119 -6299 11153 -6265
rect 10861 -6609 10895 -6575
rect 10861 -6717 10895 -6683
rect 10603 -7027 10637 -6993
rect 10603 -7135 10637 -7101
rect 11893 -5355 11927 -5321
rect 11893 -5463 11927 -5429
rect 11635 -5773 11669 -5739
rect 11635 -5881 11669 -5847
rect 11377 -6191 11411 -6157
rect 11377 -6299 11411 -6265
rect 11119 -6609 11153 -6575
rect 11119 -6717 11153 -6683
rect 10861 -7027 10895 -6993
rect 10861 -7135 10895 -7101
rect 10603 -7445 10637 -7411
rect 10603 -7553 10637 -7519
rect 12151 -5355 12185 -5321
rect 12151 -5463 12185 -5429
rect 11893 -5773 11927 -5739
rect 11893 -5881 11927 -5847
rect 11635 -6191 11669 -6157
rect 11635 -6299 11669 -6265
rect 11377 -6609 11411 -6575
rect 11377 -6717 11411 -6683
rect 11119 -7027 11153 -6993
rect 11119 -7135 11153 -7101
rect 10861 -7445 10895 -7411
rect 10861 -7553 10895 -7519
rect 10603 -7863 10637 -7829
rect 12409 -5355 12443 -5321
rect 12409 -5463 12443 -5429
rect 12151 -5773 12185 -5739
rect 12151 -5881 12185 -5847
rect 11893 -6191 11927 -6157
rect 11893 -6299 11927 -6265
rect 11635 -6609 11669 -6575
rect 11635 -6717 11669 -6683
rect 11377 -7027 11411 -6993
rect 11377 -7135 11411 -7101
rect 11119 -7445 11153 -7411
rect 11119 -7553 11153 -7519
rect 10861 -7863 10895 -7829
rect 12409 -5773 12443 -5739
rect 12409 -5881 12443 -5847
rect 12151 -6191 12185 -6157
rect 12151 -6299 12185 -6265
rect 11893 -6609 11927 -6575
rect 11893 -6717 11927 -6683
rect 11635 -7027 11669 -6993
rect 11635 -7135 11669 -7101
rect 11377 -7445 11411 -7411
rect 11377 -7553 11411 -7519
rect 11119 -7863 11153 -7829
rect 12409 -6191 12443 -6157
rect 12409 -6299 12443 -6265
rect 12151 -6609 12185 -6575
rect 12151 -6717 12185 -6683
rect 11893 -7027 11927 -6993
rect 11893 -7135 11927 -7101
rect 11635 -7445 11669 -7411
rect 11635 -7553 11669 -7519
rect 11377 -7863 11411 -7829
rect 12409 -6609 12443 -6575
rect 12409 -6717 12443 -6683
rect 12151 -7027 12185 -6993
rect 12151 -7135 12185 -7101
rect 11893 -7445 11927 -7411
rect 11893 -7553 11927 -7519
rect 11635 -7863 11669 -7829
rect 12409 -7027 12443 -6993
rect 12409 -7135 12443 -7101
rect 12151 -7445 12185 -7411
rect 12151 -7553 12185 -7519
rect 11893 -7863 11927 -7829
rect 12409 -7445 12443 -7411
rect 12409 -7553 12443 -7519
rect 12151 -7863 12185 -7829
rect 12409 -7863 12443 -7829
rect 6165 -8206 6170 -8172
rect 6170 -8206 6204 -8172
rect 6204 -8206 6215 -8172
rect 6165 -8212 6215 -8206
rect 8835 -8206 8840 -8172
rect 8840 -8206 8874 -8172
rect 8874 -8206 8885 -8172
rect 8835 -8212 8885 -8206
rect 6166 -8482 6206 -8481
rect 6166 -8516 6170 -8482
rect 6170 -8516 6204 -8482
rect 6204 -8516 6206 -8482
rect 6166 -8517 6206 -8516
rect 11498 -8205 11503 -8171
rect 11503 -8205 11537 -8171
rect 11537 -8205 11548 -8171
rect 11498 -8211 11548 -8205
rect 8836 -8482 8880 -8478
rect 8836 -8516 8840 -8482
rect 8840 -8516 8874 -8482
rect 8874 -8516 8880 -8482
rect 8836 -8521 8880 -8516
rect 11498 -8481 11542 -8477
rect 11498 -8515 11503 -8481
rect 11503 -8515 11537 -8481
rect 11537 -8515 11542 -8481
rect 11498 -8519 11542 -8515
rect 6000 -8702 6092 -8608
rect 8670 -8702 8762 -8608
rect 11336 -8702 11428 -8608
rect 3826 -9598 3862 -9538
rect 13903 -9537 13904 8629
rect 13904 -9537 13938 8629
rect 14018 7163 14052 8539
rect 17447 8629 17482 8655
rect 14018 5653 14052 7029
rect 14018 4143 14052 5519
rect 14018 2633 14052 4009
rect 14018 1123 14052 2499
rect 14018 -387 14052 989
rect 14018 -1897 14052 -521
rect 14018 -3407 14052 -2031
rect 14018 -4917 14052 -3541
rect 14018 -6427 14052 -5051
rect 14018 -7937 14052 -6561
rect 14018 -9447 14052 -8071
rect 13903 -9591 13938 -9537
rect 15676 7163 15710 8539
rect 15676 5653 15710 7029
rect 15676 4143 15710 5519
rect 15676 2633 15710 4009
rect 15676 1123 15710 2499
rect 15676 -387 15710 989
rect 15676 -1897 15710 -521
rect 15676 -3407 15710 -2031
rect 15676 -4917 15710 -3541
rect 15676 -6427 15710 -5051
rect 15676 -7937 15710 -6561
rect 15676 -9447 15710 -8071
rect 17334 7163 17368 8539
rect 17334 5653 17368 7029
rect 17334 4143 17368 5519
rect 17334 2633 17368 4009
rect 17334 1123 17368 2499
rect 17334 -387 17368 989
rect 17334 -1897 17368 -521
rect 17334 -3407 17368 -2031
rect 17334 -4917 17368 -3541
rect 17334 -6427 17368 -5051
rect 17334 -7937 17368 -6561
rect 17334 -9447 17368 -8071
rect 17447 -9537 17448 8629
rect 17448 -9537 17482 8629
rect 17447 -9591 17482 -9537
rect 274 -9600 3862 -9598
rect 274 -9634 379 -9600
rect 379 -9634 3765 -9600
rect 3765 -9634 3862 -9600
rect 274 -9635 3862 -9634
rect 13902 -9599 17487 -9591
rect 13902 -9633 14000 -9599
rect 14000 -9633 17386 -9599
rect 17386 -9633 17487 -9599
rect 274 -9641 3861 -9635
rect 13902 -9636 17487 -9633
<< metal1 >>
rect 244 8655 3900 8667
rect 244 -9598 282 8655
rect 318 8654 3900 8655
rect 318 8538 3826 8654
rect 318 7162 397 8538
rect 431 7162 2055 8538
rect 2089 7162 3713 8538
rect 3747 7162 3826 8538
rect 318 7028 3826 7162
rect 318 5652 397 7028
rect 431 5652 2055 7028
rect 2089 5652 3713 7028
rect 3747 5652 3826 7028
rect 318 5518 3826 5652
rect 318 4142 397 5518
rect 431 4142 2055 5518
rect 2089 4142 3713 5518
rect 3747 4142 3826 5518
rect 318 4008 3826 4142
rect 318 2632 397 4008
rect 431 3196 2055 4008
rect 2089 3196 3713 4008
rect 431 2706 1441 3196
rect 2738 2706 3713 3196
rect 431 2632 2055 2706
rect 2089 2632 3713 2706
rect 3747 2632 3826 4008
rect 318 2498 3826 2632
rect 318 1122 397 2498
rect 431 1122 2055 2498
rect 2089 1122 3713 2498
rect 3747 1122 3826 2498
rect 318 988 3826 1122
rect 318 -388 397 988
rect 431 -388 2055 988
rect 2089 -388 3713 988
rect 3747 -388 3826 988
rect 318 -522 3826 -388
rect 318 -1898 397 -522
rect 431 -1898 2055 -522
rect 2089 -1898 3713 -522
rect 3747 -1898 3826 -522
rect 318 -2032 3826 -1898
rect 318 -3408 397 -2032
rect 431 -3408 2055 -2032
rect 2089 -3408 3713 -2032
rect 3747 -3408 3826 -2032
rect 318 -3542 3826 -3408
rect 318 -4918 397 -3542
rect 431 -4918 2055 -3542
rect 2089 -4918 3713 -3542
rect 3747 -4918 3826 -3542
rect 318 -5052 3826 -4918
rect 318 -6428 397 -5052
rect 431 -6428 2055 -5052
rect 2089 -6428 3713 -5052
rect 3747 -6428 3826 -5052
rect 318 -6562 3826 -6428
rect 318 -7938 397 -6562
rect 431 -7938 2055 -6562
rect 2089 -7938 3713 -6562
rect 3747 -7938 3826 -6562
rect 318 -8072 3826 -7938
rect 318 -9448 397 -8072
rect 431 -9448 2055 -8072
rect 2089 -9448 3713 -8072
rect 3747 -9448 3826 -8072
rect 318 -9598 3826 -9448
rect 244 -9641 274 -9598
rect 3862 -9635 3900 8654
rect 13862 8655 17519 8663
rect 8817 8610 10506 8619
rect 5886 8579 6433 8605
rect 5886 8545 6204 8579
rect 6238 8545 6433 8579
rect 5886 8484 6433 8545
rect 5886 8323 5925 8484
rect 5988 8483 6314 8484
rect 5988 8324 6051 8483
rect 6131 8324 6202 8483
rect 6282 8325 6314 8483
rect 6394 8325 6433 8484
rect 6282 8324 6433 8325
rect 5988 8323 6433 8324
rect 5886 8251 6433 8323
rect 5886 8217 6204 8251
rect 6238 8217 6433 8251
rect 5886 8191 6433 8217
rect 8816 8578 10506 8610
rect 8816 8544 9092 8578
rect 9126 8544 9350 8578
rect 9384 8544 9608 8578
rect 9642 8544 9866 8578
rect 9900 8544 10124 8578
rect 10158 8544 10506 8578
rect 8816 8517 10506 8544
rect 8816 8291 8924 8517
rect 10483 8291 10506 8517
rect 8816 8289 10369 8291
rect 10482 8289 10506 8291
rect 8816 8250 10506 8289
rect 8816 8216 9092 8250
rect 9126 8216 9350 8250
rect 9384 8216 9608 8250
rect 9642 8216 9866 8250
rect 9900 8216 10124 8250
rect 10158 8216 10506 8250
rect 8816 8181 10506 8216
rect 8817 8178 10506 8181
rect 6099 7606 6225 7614
rect 6099 7545 6121 7606
rect 6201 7545 6225 7606
rect 5012 7519 5290 7538
rect 5012 7206 5030 7519
rect 5269 7206 5290 7519
rect 6099 7385 6225 7545
rect 6099 7324 6122 7385
rect 6202 7324 6225 7385
rect 6099 7231 6225 7324
rect 5012 7187 5290 7206
rect 6098 6852 6225 7231
rect 8775 7602 8901 7615
rect 8775 7519 8795 7602
rect 8893 7519 8901 7602
rect 8775 7407 8901 7519
rect 8775 7324 8795 7407
rect 8893 7324 8901 7407
rect 8775 7220 8901 7324
rect 11431 7602 11557 7614
rect 11431 7519 11447 7602
rect 11545 7519 11557 7602
rect 11431 7407 11557 7519
rect 11431 7324 11447 7407
rect 11545 7324 11557 7407
rect 11431 7231 11557 7324
rect 8775 6855 8900 7220
rect 4014 6824 4406 6830
rect 6098 6824 6226 6852
rect 4014 6688 6226 6824
rect 8771 6807 8900 6855
rect 8771 6728 8783 6807
rect 8878 6728 8900 6807
rect 8771 6711 8900 6728
rect 4014 5560 4406 6688
rect 4014 5342 4070 5560
rect 4316 5342 4406 5560
rect 4014 5324 4406 5342
rect 4885 6648 5045 6649
rect 6098 6648 6224 6688
rect 7335 6648 7495 6649
rect 4885 6609 7495 6648
rect 4885 6575 5270 6609
rect 5304 6575 5528 6609
rect 5562 6575 5786 6609
rect 5820 6575 6044 6609
rect 6078 6575 6302 6609
rect 6336 6575 6560 6609
rect 6594 6575 6818 6609
rect 6852 6575 7076 6609
rect 7110 6575 7495 6609
rect 4885 6549 7495 6575
rect 4885 6320 5045 6549
rect 7335 6320 7495 6549
rect 4885 6299 7495 6320
rect 4885 6265 5270 6299
rect 5304 6265 5528 6299
rect 5562 6265 5786 6299
rect 5820 6265 6044 6299
rect 6078 6265 6302 6299
rect 6336 6265 6560 6299
rect 6594 6265 6818 6299
rect 6852 6265 7076 6299
rect 7110 6265 7495 6299
rect 4885 6191 7495 6265
rect 4885 6157 5270 6191
rect 5304 6157 5528 6191
rect 5562 6157 5786 6191
rect 5820 6157 6044 6191
rect 6078 6157 6302 6191
rect 6336 6157 6560 6191
rect 6594 6157 6818 6191
rect 6852 6157 7076 6191
rect 7110 6157 7495 6191
rect 4885 6129 7495 6157
rect 4885 5910 5045 6129
rect 7335 5910 7495 6129
rect 4885 5881 7495 5910
rect 4885 5847 5270 5881
rect 5304 5847 5528 5881
rect 5562 5847 5786 5881
rect 5820 5847 6044 5881
rect 6078 5847 6302 5881
rect 6336 5847 6560 5881
rect 6594 5847 6818 5881
rect 6852 5847 7076 5881
rect 7110 5847 7495 5881
rect 4885 5773 7495 5847
rect 4885 5739 5270 5773
rect 5304 5739 5528 5773
rect 5562 5739 5786 5773
rect 5820 5739 6044 5773
rect 6078 5739 6302 5773
rect 6336 5739 6560 5773
rect 6594 5739 6818 5773
rect 6852 5739 7076 5773
rect 7110 5739 7495 5773
rect 4885 5719 7495 5739
rect 4885 5480 5045 5719
rect 7335 5480 7495 5719
rect 4885 5463 7495 5480
rect 4885 5429 5270 5463
rect 5304 5429 5528 5463
rect 5562 5429 5786 5463
rect 5820 5429 6044 5463
rect 6078 5429 6302 5463
rect 6336 5429 6560 5463
rect 6594 5429 6818 5463
rect 6852 5429 7076 5463
rect 7110 5429 7495 5463
rect 4885 5355 7495 5429
rect 4885 5321 5270 5355
rect 5304 5321 5528 5355
rect 5562 5321 5786 5355
rect 5820 5321 6044 5355
rect 6078 5321 6302 5355
rect 6336 5321 6560 5355
rect 6594 5321 6818 5355
rect 6852 5321 7076 5355
rect 7110 5321 7495 5355
rect 4885 5289 7495 5321
rect 4885 5070 5045 5289
rect 7335 5070 7495 5289
rect 4885 5045 7495 5070
rect 4885 5011 5270 5045
rect 5304 5011 5528 5045
rect 5562 5011 5786 5045
rect 5820 5011 6044 5045
rect 6078 5011 6302 5045
rect 6336 5011 6560 5045
rect 6594 5011 6818 5045
rect 6852 5011 7076 5045
rect 7110 5011 7495 5045
rect 4885 4937 7495 5011
rect 4885 4903 5270 4937
rect 5304 4903 5528 4937
rect 5562 4903 5786 4937
rect 5820 4903 6044 4937
rect 6078 4903 6302 4937
rect 6336 4903 6560 4937
rect 6594 4903 6818 4937
rect 6852 4903 7076 4937
rect 7110 4903 7495 4937
rect 4885 4879 7495 4903
rect 4885 4650 5045 4879
rect 7335 4650 7495 4879
rect 4885 4627 7495 4650
rect 4885 4593 5270 4627
rect 5304 4593 5528 4627
rect 5562 4593 5786 4627
rect 5820 4593 6044 4627
rect 6078 4593 6302 4627
rect 6336 4593 6560 4627
rect 6594 4593 6818 4627
rect 6852 4593 7076 4627
rect 7110 4593 7495 4627
rect 4885 4519 7495 4593
rect 4885 4485 5270 4519
rect 5304 4485 5528 4519
rect 5562 4485 5786 4519
rect 5820 4485 6044 4519
rect 6078 4485 6302 4519
rect 6336 4485 6560 4519
rect 6594 4485 6818 4519
rect 6852 4485 7076 4519
rect 7110 4485 7495 4519
rect 4885 4459 7495 4485
rect 4885 4240 5045 4459
rect 7335 4240 7495 4459
rect 4885 4209 7495 4240
rect 4885 4175 5270 4209
rect 5304 4175 5528 4209
rect 5562 4175 5786 4209
rect 5820 4175 6044 4209
rect 6078 4175 6302 4209
rect 6336 4175 6560 4209
rect 6594 4175 6818 4209
rect 6852 4175 7076 4209
rect 7110 4175 7495 4209
rect 4885 4101 7495 4175
rect 4885 4067 5270 4101
rect 5304 4067 5528 4101
rect 5562 4067 5786 4101
rect 5820 4067 6044 4101
rect 6078 4067 6302 4101
rect 6336 4067 6560 4101
rect 6594 4067 6818 4101
rect 6852 4067 7076 4101
rect 7110 4067 7495 4101
rect 4885 4049 7495 4067
rect 4885 3819 5045 4049
rect 7335 3819 7495 4049
rect 4885 3791 7495 3819
rect 4885 3757 5270 3791
rect 5304 3757 5528 3791
rect 5562 3757 5786 3791
rect 5820 3757 6044 3791
rect 6078 3757 6302 3791
rect 6336 3757 6560 3791
rect 6594 3757 6818 3791
rect 6852 3757 7076 3791
rect 7110 3757 7495 3791
rect 4885 3689 7495 3757
rect 7555 6648 7715 6649
rect 8774 6648 8900 6711
rect 11430 6818 11557 7231
rect 12426 7504 12727 7528
rect 12426 7183 12461 7504
rect 12683 7183 12727 7504
rect 12426 7157 12727 7183
rect 12672 6920 13550 6964
rect 11430 6807 11570 6818
rect 11430 6728 11456 6807
rect 11551 6728 11570 6807
rect 11430 6711 11570 6728
rect 12672 6742 12692 6920
rect 12860 6744 13352 6920
rect 13514 6744 13550 6920
rect 12860 6742 13550 6744
rect 10218 6649 10378 6650
rect 11430 6649 11556 6711
rect 12672 6710 13550 6742
rect 12668 6649 12828 6650
rect 10005 6648 10165 6649
rect 7555 6609 10165 6648
rect 7555 6575 7940 6609
rect 7974 6575 8198 6609
rect 8232 6575 8456 6609
rect 8490 6575 8714 6609
rect 8748 6575 8972 6609
rect 9006 6575 9230 6609
rect 9264 6575 9488 6609
rect 9522 6575 9746 6609
rect 9780 6575 10165 6609
rect 7555 6549 10165 6575
rect 7555 6320 7715 6549
rect 10005 6320 10165 6549
rect 7555 6299 10165 6320
rect 7555 6265 7940 6299
rect 7974 6265 8198 6299
rect 8232 6265 8456 6299
rect 8490 6265 8714 6299
rect 8748 6265 8972 6299
rect 9006 6265 9230 6299
rect 9264 6265 9488 6299
rect 9522 6265 9746 6299
rect 9780 6265 10165 6299
rect 7555 6191 10165 6265
rect 7555 6157 7940 6191
rect 7974 6157 8198 6191
rect 8232 6157 8456 6191
rect 8490 6157 8714 6191
rect 8748 6157 8972 6191
rect 9006 6157 9230 6191
rect 9264 6157 9488 6191
rect 9522 6157 9746 6191
rect 9780 6157 10165 6191
rect 7555 6129 10165 6157
rect 7555 5910 7715 6129
rect 10005 5910 10165 6129
rect 7555 5881 10165 5910
rect 7555 5847 7940 5881
rect 7974 5847 8198 5881
rect 8232 5847 8456 5881
rect 8490 5847 8714 5881
rect 8748 5847 8972 5881
rect 9006 5847 9230 5881
rect 9264 5847 9488 5881
rect 9522 5847 9746 5881
rect 9780 5847 10165 5881
rect 7555 5773 10165 5847
rect 7555 5739 7940 5773
rect 7974 5739 8198 5773
rect 8232 5739 8456 5773
rect 8490 5739 8714 5773
rect 8748 5739 8972 5773
rect 9006 5739 9230 5773
rect 9264 5739 9488 5773
rect 9522 5739 9746 5773
rect 9780 5739 10165 5773
rect 7555 5719 10165 5739
rect 7555 5480 7715 5719
rect 10005 5480 10165 5719
rect 7555 5463 10165 5480
rect 7555 5429 7940 5463
rect 7974 5429 8198 5463
rect 8232 5429 8456 5463
rect 8490 5429 8714 5463
rect 8748 5429 8972 5463
rect 9006 5429 9230 5463
rect 9264 5429 9488 5463
rect 9522 5429 9746 5463
rect 9780 5429 10165 5463
rect 7555 5355 10165 5429
rect 7555 5321 7940 5355
rect 7974 5321 8198 5355
rect 8232 5321 8456 5355
rect 8490 5321 8714 5355
rect 8748 5321 8972 5355
rect 9006 5321 9230 5355
rect 9264 5321 9488 5355
rect 9522 5321 9746 5355
rect 9780 5321 10165 5355
rect 7555 5289 10165 5321
rect 7555 5070 7715 5289
rect 10005 5070 10165 5289
rect 7555 5045 10165 5070
rect 7555 5011 7940 5045
rect 7974 5011 8198 5045
rect 8232 5011 8456 5045
rect 8490 5011 8714 5045
rect 8748 5011 8972 5045
rect 9006 5011 9230 5045
rect 9264 5011 9488 5045
rect 9522 5011 9746 5045
rect 9780 5011 10165 5045
rect 7555 4937 10165 5011
rect 7555 4903 7940 4937
rect 7974 4903 8198 4937
rect 8232 4903 8456 4937
rect 8490 4903 8714 4937
rect 8748 4903 8972 4937
rect 9006 4903 9230 4937
rect 9264 4903 9488 4937
rect 9522 4903 9746 4937
rect 9780 4903 10165 4937
rect 7555 4879 10165 4903
rect 7555 4650 7715 4879
rect 10005 4650 10165 4879
rect 7555 4627 10165 4650
rect 7555 4593 7940 4627
rect 7974 4593 8198 4627
rect 8232 4593 8456 4627
rect 8490 4593 8714 4627
rect 8748 4593 8972 4627
rect 9006 4593 9230 4627
rect 9264 4593 9488 4627
rect 9522 4593 9746 4627
rect 9780 4593 10165 4627
rect 7555 4519 10165 4593
rect 7555 4485 7940 4519
rect 7974 4485 8198 4519
rect 8232 4485 8456 4519
rect 8490 4485 8714 4519
rect 8748 4485 8972 4519
rect 9006 4485 9230 4519
rect 9264 4485 9488 4519
rect 9522 4485 9746 4519
rect 9780 4485 10165 4519
rect 7555 4459 10165 4485
rect 7555 4240 7715 4459
rect 10005 4240 10165 4459
rect 7555 4209 10165 4240
rect 7555 4175 7940 4209
rect 7974 4175 8198 4209
rect 8232 4175 8456 4209
rect 8490 4175 8714 4209
rect 8748 4175 8972 4209
rect 9006 4175 9230 4209
rect 9264 4175 9488 4209
rect 9522 4175 9746 4209
rect 9780 4175 10165 4209
rect 7555 4101 10165 4175
rect 7555 4067 7940 4101
rect 7974 4067 8198 4101
rect 8232 4067 8456 4101
rect 8490 4067 8714 4101
rect 8748 4067 8972 4101
rect 9006 4067 9230 4101
rect 9264 4067 9488 4101
rect 9522 4067 9746 4101
rect 9780 4067 10165 4101
rect 7555 4049 10165 4067
rect 7555 3819 7715 4049
rect 10005 3819 10165 4049
rect 7555 3791 10165 3819
rect 7555 3757 7940 3791
rect 7974 3757 8198 3791
rect 8232 3757 8456 3791
rect 8490 3757 8714 3791
rect 8748 3757 8972 3791
rect 9006 3757 9230 3791
rect 9264 3757 9488 3791
rect 9522 3757 9746 3791
rect 9780 3757 10165 3791
rect 7555 3689 10165 3757
rect 10218 6610 12828 6649
rect 10218 6576 10603 6610
rect 10637 6576 10861 6610
rect 10895 6576 11119 6610
rect 11153 6576 11377 6610
rect 11411 6576 11635 6610
rect 11669 6576 11893 6610
rect 11927 6576 12151 6610
rect 12185 6576 12409 6610
rect 12443 6576 12828 6610
rect 10218 6550 12828 6576
rect 10218 6321 10378 6550
rect 12668 6321 12828 6550
rect 10218 6300 12828 6321
rect 10218 6266 10603 6300
rect 10637 6266 10861 6300
rect 10895 6266 11119 6300
rect 11153 6266 11377 6300
rect 11411 6266 11635 6300
rect 11669 6266 11893 6300
rect 11927 6266 12151 6300
rect 12185 6266 12409 6300
rect 12443 6266 12828 6300
rect 10218 6192 12828 6266
rect 10218 6158 10603 6192
rect 10637 6158 10861 6192
rect 10895 6158 11119 6192
rect 11153 6158 11377 6192
rect 11411 6158 11635 6192
rect 11669 6158 11893 6192
rect 11927 6158 12151 6192
rect 12185 6158 12409 6192
rect 12443 6158 12828 6192
rect 10218 6130 12828 6158
rect 10218 5911 10378 6130
rect 12668 5911 12828 6130
rect 10218 5882 12828 5911
rect 10218 5848 10603 5882
rect 10637 5848 10861 5882
rect 10895 5848 11119 5882
rect 11153 5848 11377 5882
rect 11411 5848 11635 5882
rect 11669 5848 11893 5882
rect 11927 5848 12151 5882
rect 12185 5848 12409 5882
rect 12443 5848 12828 5882
rect 10218 5774 12828 5848
rect 10218 5740 10603 5774
rect 10637 5740 10861 5774
rect 10895 5740 11119 5774
rect 11153 5740 11377 5774
rect 11411 5740 11635 5774
rect 11669 5740 11893 5774
rect 11927 5740 12151 5774
rect 12185 5740 12409 5774
rect 12443 5740 12828 5774
rect 10218 5720 12828 5740
rect 10218 5481 10378 5720
rect 12668 5481 12828 5720
rect 10218 5464 12828 5481
rect 10218 5430 10603 5464
rect 10637 5430 10861 5464
rect 10895 5430 11119 5464
rect 11153 5430 11377 5464
rect 11411 5430 11635 5464
rect 11669 5430 11893 5464
rect 11927 5430 12151 5464
rect 12185 5430 12409 5464
rect 12443 5430 12828 5464
rect 10218 5356 12828 5430
rect 10218 5322 10603 5356
rect 10637 5322 10861 5356
rect 10895 5322 11119 5356
rect 11153 5322 11377 5356
rect 11411 5322 11635 5356
rect 11669 5322 11893 5356
rect 11927 5322 12151 5356
rect 12185 5322 12409 5356
rect 12443 5322 12828 5356
rect 10218 5290 12828 5322
rect 10218 5071 10378 5290
rect 12668 5071 12828 5290
rect 10218 5046 12828 5071
rect 10218 5012 10603 5046
rect 10637 5012 10861 5046
rect 10895 5012 11119 5046
rect 11153 5012 11377 5046
rect 11411 5012 11635 5046
rect 11669 5012 11893 5046
rect 11927 5012 12151 5046
rect 12185 5012 12409 5046
rect 12443 5012 12828 5046
rect 10218 4938 12828 5012
rect 10218 4904 10603 4938
rect 10637 4904 10861 4938
rect 10895 4904 11119 4938
rect 11153 4904 11377 4938
rect 11411 4904 11635 4938
rect 11669 4904 11893 4938
rect 11927 4904 12151 4938
rect 12185 4904 12409 4938
rect 12443 4904 12828 4938
rect 10218 4880 12828 4904
rect 10218 4651 10378 4880
rect 12668 4651 12828 4880
rect 10218 4628 12828 4651
rect 10218 4594 10603 4628
rect 10637 4594 10861 4628
rect 10895 4594 11119 4628
rect 11153 4594 11377 4628
rect 11411 4594 11635 4628
rect 11669 4594 11893 4628
rect 11927 4594 12151 4628
rect 12185 4594 12409 4628
rect 12443 4594 12828 4628
rect 10218 4520 12828 4594
rect 10218 4486 10603 4520
rect 10637 4486 10861 4520
rect 10895 4486 11119 4520
rect 11153 4486 11377 4520
rect 11411 4486 11635 4520
rect 11669 4486 11893 4520
rect 11927 4486 12151 4520
rect 12185 4486 12409 4520
rect 12443 4486 12828 4520
rect 10218 4460 12828 4486
rect 10218 4241 10378 4460
rect 12668 4241 12828 4460
rect 10218 4210 12828 4241
rect 10218 4176 10603 4210
rect 10637 4176 10861 4210
rect 10895 4176 11119 4210
rect 11153 4176 11377 4210
rect 11411 4176 11635 4210
rect 11669 4176 11893 4210
rect 11927 4176 12151 4210
rect 12185 4176 12409 4210
rect 12443 4176 12828 4210
rect 10218 4102 12828 4176
rect 10218 4068 10603 4102
rect 10637 4068 10861 4102
rect 10895 4068 11119 4102
rect 11153 4068 11377 4102
rect 11411 4068 11635 4102
rect 11669 4068 11893 4102
rect 11927 4068 12151 4102
rect 12185 4068 12409 4102
rect 12443 4068 12828 4102
rect 10218 4050 12828 4068
rect 10218 3820 10378 4050
rect 12668 3820 12828 4050
rect 10218 3792 12828 3820
rect 10218 3758 10603 3792
rect 10637 3758 10861 3792
rect 10895 3758 11119 3792
rect 11153 3758 11377 3792
rect 11411 3758 11635 3792
rect 11669 3758 11893 3792
rect 11927 3758 12151 3792
rect 12185 3758 12409 3792
rect 12443 3758 12828 3792
rect 10218 3690 12828 3758
rect 13322 5994 13550 6010
rect 13322 5818 13352 5994
rect 13514 5818 13550 5994
rect 6135 3449 6245 3689
rect 6135 3409 6165 3449
rect 6215 3409 6245 3449
rect 6135 3142 6245 3409
rect 6135 3102 6168 3142
rect 6206 3102 6245 3142
rect 6135 3081 6245 3102
rect 8805 3449 8915 3689
rect 8805 3409 8835 3449
rect 8885 3409 8915 3449
rect 8805 3142 8915 3409
rect 8805 3102 8838 3142
rect 8876 3102 8915 3142
rect 8805 3078 8915 3102
rect 11468 3450 11578 3690
rect 11468 3410 11498 3450
rect 11548 3410 11578 3450
rect 11468 3142 11578 3410
rect 11468 3102 11500 3142
rect 11538 3102 11578 3142
rect 11468 3087 11578 3102
rect 5978 3012 6122 3020
rect 5978 2906 5998 3012
rect 6104 2906 6122 3012
rect 5978 2896 6122 2906
rect 8644 3012 8788 3020
rect 8644 2906 8662 3012
rect 8768 2906 8788 3012
rect 8644 2896 8788 2906
rect 11305 3012 11451 3020
rect 11305 2906 11324 3012
rect 11430 2906 11451 3012
rect 11305 2895 11451 2906
rect 13322 2156 13550 5818
rect 13318 2112 13550 2156
rect 4979 1953 5257 1967
rect 4979 1648 5019 1953
rect 5202 1648 5257 1953
rect 13318 1936 13352 2112
rect 13514 1936 13550 2112
rect 4979 1616 5257 1648
rect 6097 1924 6223 1932
rect 6097 1863 6121 1924
rect 6201 1863 6223 1924
rect 6097 1703 6223 1863
rect 6097 1642 6120 1703
rect 6200 1642 6223 1703
rect 6097 1635 6223 1642
rect 8768 1920 8894 1933
rect 8768 1837 8776 1920
rect 8874 1837 8894 1920
rect 8768 1725 8894 1837
rect 8768 1642 8776 1725
rect 8874 1642 8894 1725
rect 8768 1635 8894 1642
rect 11439 1920 11565 1932
rect 11439 1837 11451 1920
rect 11549 1837 11565 1920
rect 13318 1902 13550 1936
rect 11439 1725 11565 1837
rect 11439 1642 11451 1725
rect 11549 1642 11565 1725
rect 11439 1635 11565 1642
rect 4060 1166 5084 1200
rect 4060 1114 4884 1166
rect 4060 938 4098 1114
rect 4260 1002 4884 1114
rect 5042 1002 5084 1166
rect 4260 980 5084 1002
rect 6098 1144 6224 1635
rect 8774 1144 8900 1635
rect 6098 1116 7746 1144
rect 6098 982 7590 1116
rect 7708 982 7746 1116
rect 8774 1106 10330 1144
rect 8774 1101 10196 1106
rect 8771 994 10196 1101
rect 4260 938 4296 980
rect 4060 904 4296 938
rect 6098 972 7746 982
rect 8774 982 10196 994
rect 10308 982 10330 1106
rect 4885 931 5045 932
rect 6098 931 6224 972
rect 8774 968 10330 982
rect 11430 1134 11556 1635
rect 13322 1186 13550 1202
rect 13322 1134 13352 1186
rect 11430 1010 13352 1134
rect 13514 1010 13550 1186
rect 11430 994 13550 1010
rect 11430 992 13320 994
rect 7335 931 7495 932
rect 4885 892 7495 931
rect 4885 858 5270 892
rect 5304 858 5528 892
rect 5562 858 5786 892
rect 5820 858 6044 892
rect 6078 858 6302 892
rect 6336 858 6560 892
rect 6594 858 6818 892
rect 6852 858 7076 892
rect 7110 858 7495 892
rect 4885 832 7495 858
rect 4885 603 5045 832
rect 7335 603 7495 832
rect 4885 582 7495 603
rect 4885 548 5270 582
rect 5304 548 5528 582
rect 5562 548 5786 582
rect 5820 548 6044 582
rect 6078 548 6302 582
rect 6336 548 6560 582
rect 6594 548 6818 582
rect 6852 548 7076 582
rect 7110 548 7495 582
rect 4885 474 7495 548
rect 4885 440 5270 474
rect 5304 440 5528 474
rect 5562 440 5786 474
rect 5820 440 6044 474
rect 6078 440 6302 474
rect 6336 440 6560 474
rect 6594 440 6818 474
rect 6852 440 7076 474
rect 7110 440 7495 474
rect 4885 412 7495 440
rect 4068 188 4296 204
rect 4068 12 4098 188
rect 4260 12 4296 188
rect 4068 -3868 4296 12
rect 4885 193 5045 412
rect 7335 193 7495 412
rect 4885 164 7495 193
rect 4885 130 5270 164
rect 5304 130 5528 164
rect 5562 130 5786 164
rect 5820 130 6044 164
rect 6078 130 6302 164
rect 6336 130 6560 164
rect 6594 130 6818 164
rect 6852 130 7076 164
rect 7110 130 7495 164
rect 4885 56 7495 130
rect 4885 22 5270 56
rect 5304 22 5528 56
rect 5562 22 5786 56
rect 5820 22 6044 56
rect 6078 22 6302 56
rect 6336 22 6560 56
rect 6594 22 6818 56
rect 6852 22 7076 56
rect 7110 22 7495 56
rect 4885 2 7495 22
rect 4885 -237 5045 2
rect 7335 -237 7495 2
rect 4885 -254 7495 -237
rect 4885 -288 5270 -254
rect 5304 -288 5528 -254
rect 5562 -288 5786 -254
rect 5820 -288 6044 -254
rect 6078 -288 6302 -254
rect 6336 -288 6560 -254
rect 6594 -288 6818 -254
rect 6852 -288 7076 -254
rect 7110 -288 7495 -254
rect 4885 -362 7495 -288
rect 4885 -396 5270 -362
rect 5304 -396 5528 -362
rect 5562 -396 5786 -362
rect 5820 -396 6044 -362
rect 6078 -396 6302 -362
rect 6336 -396 6560 -362
rect 6594 -396 6818 -362
rect 6852 -396 7076 -362
rect 7110 -396 7495 -362
rect 4885 -428 7495 -396
rect 4885 -647 5045 -428
rect 7335 -647 7495 -428
rect 4885 -672 7495 -647
rect 4885 -706 5270 -672
rect 5304 -706 5528 -672
rect 5562 -706 5786 -672
rect 5820 -706 6044 -672
rect 6078 -706 6302 -672
rect 6336 -706 6560 -672
rect 6594 -706 6818 -672
rect 6852 -706 7076 -672
rect 7110 -706 7495 -672
rect 4885 -780 7495 -706
rect 4885 -814 5270 -780
rect 5304 -814 5528 -780
rect 5562 -814 5786 -780
rect 5820 -814 6044 -780
rect 6078 -814 6302 -780
rect 6336 -814 6560 -780
rect 6594 -814 6818 -780
rect 6852 -814 7076 -780
rect 7110 -814 7495 -780
rect 4885 -838 7495 -814
rect 4885 -1067 5045 -838
rect 7335 -1067 7495 -838
rect 4885 -1090 7495 -1067
rect 4885 -1124 5270 -1090
rect 5304 -1124 5528 -1090
rect 5562 -1124 5786 -1090
rect 5820 -1124 6044 -1090
rect 6078 -1124 6302 -1090
rect 6336 -1124 6560 -1090
rect 6594 -1124 6818 -1090
rect 6852 -1124 7076 -1090
rect 7110 -1124 7495 -1090
rect 4885 -1198 7495 -1124
rect 4885 -1232 5270 -1198
rect 5304 -1232 5528 -1198
rect 5562 -1232 5786 -1198
rect 5820 -1232 6044 -1198
rect 6078 -1232 6302 -1198
rect 6336 -1232 6560 -1198
rect 6594 -1232 6818 -1198
rect 6852 -1232 7076 -1198
rect 7110 -1232 7495 -1198
rect 4885 -1258 7495 -1232
rect 4885 -1477 5045 -1258
rect 7335 -1477 7495 -1258
rect 4885 -1508 7495 -1477
rect 4885 -1542 5270 -1508
rect 5304 -1542 5528 -1508
rect 5562 -1542 5786 -1508
rect 5820 -1542 6044 -1508
rect 6078 -1542 6302 -1508
rect 6336 -1542 6560 -1508
rect 6594 -1542 6818 -1508
rect 6852 -1542 7076 -1508
rect 7110 -1542 7495 -1508
rect 4885 -1616 7495 -1542
rect 4885 -1650 5270 -1616
rect 5304 -1650 5528 -1616
rect 5562 -1650 5786 -1616
rect 5820 -1650 6044 -1616
rect 6078 -1650 6302 -1616
rect 6336 -1650 6560 -1616
rect 6594 -1650 6818 -1616
rect 6852 -1650 7076 -1616
rect 7110 -1650 7495 -1616
rect 4885 -1668 7495 -1650
rect 4885 -1898 5045 -1668
rect 7335 -1898 7495 -1668
rect 4885 -1926 7495 -1898
rect 4885 -1960 5270 -1926
rect 5304 -1960 5528 -1926
rect 5562 -1960 5786 -1926
rect 5820 -1960 6044 -1926
rect 6078 -1960 6302 -1926
rect 6336 -1960 6560 -1926
rect 6594 -1960 6818 -1926
rect 6852 -1960 7076 -1926
rect 7110 -1960 7495 -1926
rect 4885 -2028 7495 -1960
rect 7555 931 7715 932
rect 8774 931 8900 968
rect 10218 932 10378 933
rect 11430 932 11556 992
rect 12668 932 12828 933
rect 10005 931 10165 932
rect 7555 892 10165 931
rect 7555 858 7940 892
rect 7974 858 8198 892
rect 8232 858 8456 892
rect 8490 858 8714 892
rect 8748 858 8972 892
rect 9006 858 9230 892
rect 9264 858 9488 892
rect 9522 858 9746 892
rect 9780 858 10165 892
rect 7555 832 10165 858
rect 7555 603 7715 832
rect 10005 603 10165 832
rect 7555 582 10165 603
rect 7555 548 7940 582
rect 7974 548 8198 582
rect 8232 548 8456 582
rect 8490 548 8714 582
rect 8748 548 8972 582
rect 9006 548 9230 582
rect 9264 548 9488 582
rect 9522 548 9746 582
rect 9780 548 10165 582
rect 7555 474 10165 548
rect 7555 440 7940 474
rect 7974 440 8198 474
rect 8232 440 8456 474
rect 8490 440 8714 474
rect 8748 440 8972 474
rect 9006 440 9230 474
rect 9264 440 9488 474
rect 9522 440 9746 474
rect 9780 440 10165 474
rect 7555 412 10165 440
rect 7555 193 7715 412
rect 10005 193 10165 412
rect 7555 164 10165 193
rect 7555 130 7940 164
rect 7974 130 8198 164
rect 8232 130 8456 164
rect 8490 130 8714 164
rect 8748 130 8972 164
rect 9006 130 9230 164
rect 9264 130 9488 164
rect 9522 130 9746 164
rect 9780 130 10165 164
rect 7555 56 10165 130
rect 7555 22 7940 56
rect 7974 22 8198 56
rect 8232 22 8456 56
rect 8490 22 8714 56
rect 8748 22 8972 56
rect 9006 22 9230 56
rect 9264 22 9488 56
rect 9522 22 9746 56
rect 9780 22 10165 56
rect 7555 2 10165 22
rect 7555 -237 7715 2
rect 10005 -237 10165 2
rect 7555 -254 10165 -237
rect 7555 -288 7940 -254
rect 7974 -288 8198 -254
rect 8232 -288 8456 -254
rect 8490 -288 8714 -254
rect 8748 -288 8972 -254
rect 9006 -288 9230 -254
rect 9264 -288 9488 -254
rect 9522 -288 9746 -254
rect 9780 -288 10165 -254
rect 7555 -362 10165 -288
rect 7555 -396 7940 -362
rect 7974 -396 8198 -362
rect 8232 -396 8456 -362
rect 8490 -396 8714 -362
rect 8748 -396 8972 -362
rect 9006 -396 9230 -362
rect 9264 -396 9488 -362
rect 9522 -396 9746 -362
rect 9780 -396 10165 -362
rect 7555 -428 10165 -396
rect 7555 -647 7715 -428
rect 10005 -647 10165 -428
rect 7555 -672 10165 -647
rect 7555 -706 7940 -672
rect 7974 -706 8198 -672
rect 8232 -706 8456 -672
rect 8490 -706 8714 -672
rect 8748 -706 8972 -672
rect 9006 -706 9230 -672
rect 9264 -706 9488 -672
rect 9522 -706 9746 -672
rect 9780 -706 10165 -672
rect 7555 -780 10165 -706
rect 7555 -814 7940 -780
rect 7974 -814 8198 -780
rect 8232 -814 8456 -780
rect 8490 -814 8714 -780
rect 8748 -814 8972 -780
rect 9006 -814 9230 -780
rect 9264 -814 9488 -780
rect 9522 -814 9746 -780
rect 9780 -814 10165 -780
rect 7555 -838 10165 -814
rect 7555 -1067 7715 -838
rect 10005 -1067 10165 -838
rect 7555 -1090 10165 -1067
rect 7555 -1124 7940 -1090
rect 7974 -1124 8198 -1090
rect 8232 -1124 8456 -1090
rect 8490 -1124 8714 -1090
rect 8748 -1124 8972 -1090
rect 9006 -1124 9230 -1090
rect 9264 -1124 9488 -1090
rect 9522 -1124 9746 -1090
rect 9780 -1124 10165 -1090
rect 7555 -1198 10165 -1124
rect 7555 -1232 7940 -1198
rect 7974 -1232 8198 -1198
rect 8232 -1232 8456 -1198
rect 8490 -1232 8714 -1198
rect 8748 -1232 8972 -1198
rect 9006 -1232 9230 -1198
rect 9264 -1232 9488 -1198
rect 9522 -1232 9746 -1198
rect 9780 -1232 10165 -1198
rect 7555 -1258 10165 -1232
rect 7555 -1477 7715 -1258
rect 10005 -1477 10165 -1258
rect 7555 -1508 10165 -1477
rect 7555 -1542 7940 -1508
rect 7974 -1542 8198 -1508
rect 8232 -1542 8456 -1508
rect 8490 -1542 8714 -1508
rect 8748 -1542 8972 -1508
rect 9006 -1542 9230 -1508
rect 9264 -1542 9488 -1508
rect 9522 -1542 9746 -1508
rect 9780 -1542 10165 -1508
rect 7555 -1616 10165 -1542
rect 7555 -1650 7940 -1616
rect 7974 -1650 8198 -1616
rect 8232 -1650 8456 -1616
rect 8490 -1650 8714 -1616
rect 8748 -1650 8972 -1616
rect 9006 -1650 9230 -1616
rect 9264 -1650 9488 -1616
rect 9522 -1650 9746 -1616
rect 9780 -1650 10165 -1616
rect 7555 -1668 10165 -1650
rect 7555 -1898 7715 -1668
rect 10005 -1898 10165 -1668
rect 7555 -1926 10165 -1898
rect 7555 -1960 7940 -1926
rect 7974 -1960 8198 -1926
rect 8232 -1960 8456 -1926
rect 8490 -1960 8714 -1926
rect 8748 -1960 8972 -1926
rect 9006 -1960 9230 -1926
rect 9264 -1960 9488 -1926
rect 9522 -1960 9746 -1926
rect 9780 -1960 10165 -1926
rect 7555 -2028 10165 -1960
rect 10218 893 12828 932
rect 10218 859 10603 893
rect 10637 859 10861 893
rect 10895 859 11119 893
rect 11153 859 11377 893
rect 11411 859 11635 893
rect 11669 859 11893 893
rect 11927 859 12151 893
rect 12185 859 12409 893
rect 12443 859 12828 893
rect 10218 833 12828 859
rect 10218 604 10378 833
rect 12668 604 12828 833
rect 10218 583 12828 604
rect 10218 549 10603 583
rect 10637 549 10861 583
rect 10895 549 11119 583
rect 11153 549 11377 583
rect 11411 549 11635 583
rect 11669 549 11893 583
rect 11927 549 12151 583
rect 12185 549 12409 583
rect 12443 549 12828 583
rect 10218 475 12828 549
rect 10218 441 10603 475
rect 10637 441 10861 475
rect 10895 441 11119 475
rect 11153 441 11377 475
rect 11411 441 11635 475
rect 11669 441 11893 475
rect 11927 441 12151 475
rect 12185 441 12409 475
rect 12443 441 12828 475
rect 10218 413 12828 441
rect 10218 194 10378 413
rect 12668 194 12828 413
rect 10218 165 12828 194
rect 10218 131 10603 165
rect 10637 131 10861 165
rect 10895 131 11119 165
rect 11153 131 11377 165
rect 11411 131 11635 165
rect 11669 131 11893 165
rect 11927 131 12151 165
rect 12185 131 12409 165
rect 12443 131 12828 165
rect 10218 57 12828 131
rect 10218 23 10603 57
rect 10637 23 10861 57
rect 10895 23 11119 57
rect 11153 23 11377 57
rect 11411 23 11635 57
rect 11669 23 11893 57
rect 11927 23 12151 57
rect 12185 23 12409 57
rect 12443 23 12828 57
rect 10218 3 12828 23
rect 10218 -236 10378 3
rect 12668 -236 12828 3
rect 10218 -253 12828 -236
rect 10218 -287 10603 -253
rect 10637 -287 10861 -253
rect 10895 -287 11119 -253
rect 11153 -287 11377 -253
rect 11411 -287 11635 -253
rect 11669 -287 11893 -253
rect 11927 -287 12151 -253
rect 12185 -287 12409 -253
rect 12443 -287 12828 -253
rect 10218 -361 12828 -287
rect 10218 -395 10603 -361
rect 10637 -395 10861 -361
rect 10895 -395 11119 -361
rect 11153 -395 11377 -361
rect 11411 -395 11635 -361
rect 11669 -395 11893 -361
rect 11927 -395 12151 -361
rect 12185 -395 12409 -361
rect 12443 -395 12828 -361
rect 10218 -427 12828 -395
rect 10218 -646 10378 -427
rect 12668 -646 12828 -427
rect 10218 -671 12828 -646
rect 10218 -705 10603 -671
rect 10637 -705 10861 -671
rect 10895 -705 11119 -671
rect 11153 -705 11377 -671
rect 11411 -705 11635 -671
rect 11669 -705 11893 -671
rect 11927 -705 12151 -671
rect 12185 -705 12409 -671
rect 12443 -705 12828 -671
rect 10218 -779 12828 -705
rect 10218 -813 10603 -779
rect 10637 -813 10861 -779
rect 10895 -813 11119 -779
rect 11153 -813 11377 -779
rect 11411 -813 11635 -779
rect 11669 -813 11893 -779
rect 11927 -813 12151 -779
rect 12185 -813 12409 -779
rect 12443 -813 12828 -779
rect 10218 -837 12828 -813
rect 10218 -1066 10378 -837
rect 12668 -1066 12828 -837
rect 10218 -1089 12828 -1066
rect 10218 -1123 10603 -1089
rect 10637 -1123 10861 -1089
rect 10895 -1123 11119 -1089
rect 11153 -1123 11377 -1089
rect 11411 -1123 11635 -1089
rect 11669 -1123 11893 -1089
rect 11927 -1123 12151 -1089
rect 12185 -1123 12409 -1089
rect 12443 -1123 12828 -1089
rect 10218 -1197 12828 -1123
rect 10218 -1231 10603 -1197
rect 10637 -1231 10861 -1197
rect 10895 -1231 11119 -1197
rect 11153 -1231 11377 -1197
rect 11411 -1231 11635 -1197
rect 11669 -1231 11893 -1197
rect 11927 -1231 12151 -1197
rect 12185 -1231 12409 -1197
rect 12443 -1231 12828 -1197
rect 10218 -1257 12828 -1231
rect 10218 -1476 10378 -1257
rect 12668 -1476 12828 -1257
rect 10218 -1507 12828 -1476
rect 10218 -1541 10603 -1507
rect 10637 -1541 10861 -1507
rect 10895 -1541 11119 -1507
rect 11153 -1541 11377 -1507
rect 11411 -1541 11635 -1507
rect 11669 -1541 11893 -1507
rect 11927 -1541 12151 -1507
rect 12185 -1541 12409 -1507
rect 12443 -1541 12828 -1507
rect 10218 -1615 12828 -1541
rect 10218 -1649 10603 -1615
rect 10637 -1649 10861 -1615
rect 10895 -1649 11119 -1615
rect 11153 -1649 11377 -1615
rect 11411 -1649 11635 -1615
rect 11669 -1649 11893 -1615
rect 11927 -1649 12151 -1615
rect 12185 -1649 12409 -1615
rect 12443 -1649 12828 -1615
rect 10218 -1667 12828 -1649
rect 10218 -1897 10378 -1667
rect 12668 -1897 12828 -1667
rect 10218 -1925 12828 -1897
rect 10218 -1959 10603 -1925
rect 10637 -1959 10861 -1925
rect 10895 -1959 11119 -1925
rect 11153 -1959 11377 -1925
rect 11411 -1959 11635 -1925
rect 11669 -1959 11893 -1925
rect 11927 -1959 12151 -1925
rect 12185 -1959 12409 -1925
rect 12443 -1959 12828 -1925
rect 10218 -2027 12828 -1959
rect 6135 -2268 6245 -2028
rect 6135 -2292 6165 -2268
rect 6134 -2308 6165 -2292
rect 6215 -2292 6245 -2268
rect 8805 -2268 8915 -2028
rect 8805 -2274 8835 -2268
rect 6215 -2308 6246 -2292
rect 6134 -2576 6246 -2308
rect 6134 -2614 6168 -2576
rect 6208 -2614 6246 -2576
rect 6134 -2648 6246 -2614
rect 8804 -2308 8835 -2274
rect 8885 -2274 8915 -2268
rect 11468 -2267 11578 -2027
rect 8885 -2308 8916 -2274
rect 8804 -2576 8916 -2308
rect 8804 -2614 8838 -2576
rect 8878 -2614 8916 -2576
rect 8804 -2636 8916 -2614
rect 11468 -2307 11498 -2267
rect 11548 -2307 11578 -2267
rect 11468 -2574 11578 -2307
rect 11468 -2616 11498 -2574
rect 11540 -2616 11578 -2574
rect 11468 -2630 11578 -2616
rect 5970 -2707 6124 -2697
rect 5970 -2813 5992 -2707
rect 6098 -2813 6124 -2707
rect 5970 -2824 6124 -2813
rect 8654 -2712 8779 -2696
rect 8654 -2806 8668 -2712
rect 8760 -2806 8779 -2712
rect 8654 -2818 8779 -2806
rect 11318 -2712 11443 -2692
rect 11318 -2806 11334 -2712
rect 11426 -2806 11443 -2712
rect 11318 -2818 11443 -2806
rect 12678 -3368 12800 -3340
rect 12234 -3404 12518 -3376
rect 12234 -3405 12275 -3404
rect 12477 -3405 12518 -3404
rect 12234 -3722 12270 -3405
rect 12486 -3722 12518 -3405
rect 12234 -3738 12518 -3722
rect 12678 -3402 12726 -3368
rect 12760 -3402 12800 -3368
rect 4068 -4044 4098 -3868
rect 4260 -4044 4296 -3868
rect 12678 -3832 12800 -3402
rect 13068 -3370 13212 -3342
rect 13068 -3404 13116 -3370
rect 13150 -3404 13212 -3370
rect 12898 -3574 13002 -3555
rect 12898 -3646 12915 -3574
rect 12986 -3646 13002 -3574
rect 12898 -3666 13002 -3646
rect 12678 -3866 12726 -3832
rect 12760 -3866 12800 -3832
rect 4068 -4078 4296 -4044
rect 4978 -3946 5165 -3929
rect 4978 -4218 4991 -3946
rect 5147 -4218 5165 -3946
rect 4978 -4246 5165 -4218
rect 6099 -4001 6225 -3993
rect 6099 -4062 6121 -4001
rect 6201 -4062 6225 -4001
rect 6099 -4222 6225 -4062
rect 6099 -4283 6122 -4222
rect 6202 -4283 6225 -4222
rect 6099 -4700 6225 -4283
rect 4068 -4716 6225 -4700
rect 4068 -4892 4098 -4716
rect 4260 -4743 6225 -4716
rect 8775 -4005 8901 -3992
rect 8775 -4088 8795 -4005
rect 8893 -4088 8901 -4005
rect 8775 -4200 8901 -4088
rect 8775 -4283 8795 -4200
rect 8893 -4283 8901 -4200
rect 8775 -4741 8901 -4283
rect 11431 -4005 11557 -3993
rect 11431 -4088 11447 -4005
rect 11545 -4088 11557 -4005
rect 11431 -4200 11557 -4088
rect 11431 -4283 11447 -4200
rect 11545 -4283 11557 -4200
rect 12678 -4164 12800 -3866
rect 13068 -3834 13212 -3404
rect 13068 -3868 13116 -3834
rect 13150 -3868 13212 -3834
rect 13068 -3996 13212 -3868
rect 12864 -4008 13212 -3996
rect 13393 -3998 13787 -3997
rect 12864 -4046 12876 -4008
rect 12930 -4046 13212 -4008
rect 12864 -4056 13212 -4046
rect 12864 -4058 12950 -4056
rect 12678 -4198 12730 -4164
rect 12764 -4198 12800 -4164
rect 11431 -4364 11557 -4283
rect 12528 -4242 12631 -4216
rect 12528 -4315 12551 -4242
rect 12607 -4315 12631 -4242
rect 12528 -4342 12631 -4315
rect 4260 -4892 6224 -4743
rect 8774 -4761 8901 -4741
rect 8774 -4803 8900 -4761
rect 4068 -4910 6224 -4892
rect 8771 -4814 8900 -4803
rect 8771 -4893 8783 -4814
rect 8878 -4893 8900 -4814
rect 8771 -4910 8900 -4893
rect 4884 -4973 5050 -4970
rect 6098 -4973 6224 -4910
rect 7335 -4973 7495 -4972
rect 4884 -5012 7495 -4973
rect 4884 -5046 5270 -5012
rect 5304 -5046 5528 -5012
rect 5562 -5046 5786 -5012
rect 5820 -5046 6044 -5012
rect 6078 -5046 6302 -5012
rect 6336 -5046 6560 -5012
rect 6594 -5046 6818 -5012
rect 6852 -5046 7076 -5012
rect 7110 -5046 7495 -5012
rect 4884 -5071 7495 -5046
rect 4885 -5072 7495 -5071
rect 4885 -5301 5045 -5072
rect 7335 -5301 7495 -5072
rect 4885 -5322 7495 -5301
rect 4885 -5356 5270 -5322
rect 5304 -5356 5528 -5322
rect 5562 -5356 5786 -5322
rect 5820 -5356 6044 -5322
rect 6078 -5356 6302 -5322
rect 6336 -5356 6560 -5322
rect 6594 -5356 6818 -5322
rect 6852 -5356 7076 -5322
rect 7110 -5356 7495 -5322
rect 4885 -5430 7495 -5356
rect 4885 -5464 5270 -5430
rect 5304 -5464 5528 -5430
rect 5562 -5464 5786 -5430
rect 5820 -5464 6044 -5430
rect 6078 -5464 6302 -5430
rect 6336 -5464 6560 -5430
rect 6594 -5464 6818 -5430
rect 6852 -5464 7076 -5430
rect 7110 -5464 7495 -5430
rect 4885 -5492 7495 -5464
rect 4885 -5711 5045 -5492
rect 7335 -5711 7495 -5492
rect 4885 -5740 7495 -5711
rect 4885 -5774 5270 -5740
rect 5304 -5774 5528 -5740
rect 5562 -5774 5786 -5740
rect 5820 -5774 6044 -5740
rect 6078 -5774 6302 -5740
rect 6336 -5774 6560 -5740
rect 6594 -5774 6818 -5740
rect 6852 -5774 7076 -5740
rect 7110 -5774 7495 -5740
rect 4885 -5848 7495 -5774
rect 4885 -5882 5270 -5848
rect 5304 -5882 5528 -5848
rect 5562 -5882 5786 -5848
rect 5820 -5882 6044 -5848
rect 6078 -5882 6302 -5848
rect 6336 -5882 6560 -5848
rect 6594 -5882 6818 -5848
rect 6852 -5882 7076 -5848
rect 7110 -5882 7495 -5848
rect 4885 -5902 7495 -5882
rect 4885 -6141 5045 -5902
rect 7335 -6141 7495 -5902
rect 4885 -6158 7495 -6141
rect 4885 -6192 5270 -6158
rect 5304 -6192 5528 -6158
rect 5562 -6192 5786 -6158
rect 5820 -6192 6044 -6158
rect 6078 -6192 6302 -6158
rect 6336 -6192 6560 -6158
rect 6594 -6192 6818 -6158
rect 6852 -6192 7076 -6158
rect 7110 -6192 7495 -6158
rect 4885 -6266 7495 -6192
rect 4885 -6300 5270 -6266
rect 5304 -6300 5528 -6266
rect 5562 -6300 5786 -6266
rect 5820 -6300 6044 -6266
rect 6078 -6300 6302 -6266
rect 6336 -6300 6560 -6266
rect 6594 -6300 6818 -6266
rect 6852 -6300 7076 -6266
rect 7110 -6300 7495 -6266
rect 4885 -6332 7495 -6300
rect 4885 -6551 5045 -6332
rect 7335 -6551 7495 -6332
rect 4885 -6576 7495 -6551
rect 4885 -6610 5270 -6576
rect 5304 -6610 5528 -6576
rect 5562 -6610 5786 -6576
rect 5820 -6610 6044 -6576
rect 6078 -6610 6302 -6576
rect 6336 -6610 6560 -6576
rect 6594 -6610 6818 -6576
rect 6852 -6610 7076 -6576
rect 7110 -6610 7495 -6576
rect 4885 -6684 7495 -6610
rect 4885 -6718 5270 -6684
rect 5304 -6718 5528 -6684
rect 5562 -6718 5786 -6684
rect 5820 -6718 6044 -6684
rect 6078 -6718 6302 -6684
rect 6336 -6718 6560 -6684
rect 6594 -6718 6818 -6684
rect 6852 -6718 7076 -6684
rect 7110 -6718 7495 -6684
rect 4885 -6742 7495 -6718
rect 4885 -6971 5045 -6742
rect 7335 -6971 7495 -6742
rect 4885 -6994 7495 -6971
rect 4885 -7028 5270 -6994
rect 5304 -7028 5528 -6994
rect 5562 -7028 5786 -6994
rect 5820 -7028 6044 -6994
rect 6078 -7028 6302 -6994
rect 6336 -7028 6560 -6994
rect 6594 -7028 6818 -6994
rect 6852 -7028 7076 -6994
rect 7110 -7028 7495 -6994
rect 4885 -7102 7495 -7028
rect 4885 -7136 5270 -7102
rect 5304 -7136 5528 -7102
rect 5562 -7136 5786 -7102
rect 5820 -7136 6044 -7102
rect 6078 -7136 6302 -7102
rect 6336 -7136 6560 -7102
rect 6594 -7136 6818 -7102
rect 6852 -7136 7076 -7102
rect 7110 -7136 7495 -7102
rect 4885 -7162 7495 -7136
rect 4885 -7381 5045 -7162
rect 7335 -7381 7495 -7162
rect 4885 -7412 7495 -7381
rect 4885 -7446 5270 -7412
rect 5304 -7446 5528 -7412
rect 5562 -7446 5786 -7412
rect 5820 -7446 6044 -7412
rect 6078 -7446 6302 -7412
rect 6336 -7446 6560 -7412
rect 6594 -7446 6818 -7412
rect 6852 -7446 7076 -7412
rect 7110 -7446 7495 -7412
rect 4885 -7520 7495 -7446
rect 4885 -7554 5270 -7520
rect 5304 -7554 5528 -7520
rect 5562 -7554 5786 -7520
rect 5820 -7554 6044 -7520
rect 6078 -7554 6302 -7520
rect 6336 -7554 6560 -7520
rect 6594 -7554 6818 -7520
rect 6852 -7554 7076 -7520
rect 7110 -7554 7495 -7520
rect 4885 -7572 7495 -7554
rect 4885 -7802 5045 -7572
rect 7335 -7802 7495 -7572
rect 4885 -7830 7495 -7802
rect 4885 -7864 5270 -7830
rect 5304 -7864 5528 -7830
rect 5562 -7864 5786 -7830
rect 5820 -7864 6044 -7830
rect 6078 -7864 6302 -7830
rect 6336 -7864 6560 -7830
rect 6594 -7864 6818 -7830
rect 6852 -7864 7076 -7830
rect 7110 -7864 7495 -7830
rect 4885 -7932 7495 -7864
rect 7555 -4973 7715 -4972
rect 8774 -4973 8900 -4910
rect 11430 -4767 11557 -4364
rect 12678 -4358 12800 -4198
rect 13068 -4164 13212 -4056
rect 13250 -4010 13787 -3998
rect 13250 -4054 13264 -4010
rect 13312 -4054 13787 -4010
rect 13250 -4062 13787 -4054
rect 13068 -4198 13120 -4164
rect 13154 -4198 13212 -4164
rect 12915 -4242 13018 -4214
rect 12915 -4315 12940 -4242
rect 12996 -4315 13018 -4242
rect 12915 -4340 13018 -4315
rect 12678 -4392 12730 -4358
rect 12764 -4392 12800 -4358
rect 12678 -4520 12800 -4392
rect 13068 -4358 13212 -4198
rect 13068 -4392 13120 -4358
rect 13154 -4392 13212 -4358
rect 13068 -4420 13212 -4392
rect 12526 -4568 13526 -4520
rect 11430 -4803 11556 -4767
rect 11430 -4814 11570 -4803
rect 11430 -4893 11456 -4814
rect 11551 -4893 11570 -4814
rect 11430 -4910 11570 -4893
rect 12526 -4858 12570 -4568
rect 12820 -4570 13526 -4568
rect 12820 -4858 13192 -4570
rect 12526 -4866 13192 -4858
rect 13444 -4866 13526 -4570
rect 10218 -4972 10378 -4971
rect 11430 -4972 11556 -4910
rect 12526 -4912 13526 -4866
rect 12668 -4972 12828 -4971
rect 10005 -4973 10165 -4972
rect 7555 -5012 10165 -4973
rect 7555 -5046 7940 -5012
rect 7974 -5046 8198 -5012
rect 8232 -5046 8456 -5012
rect 8490 -5046 8714 -5012
rect 8748 -5046 8972 -5012
rect 9006 -5046 9230 -5012
rect 9264 -5046 9488 -5012
rect 9522 -5046 9746 -5012
rect 9780 -5046 10165 -5012
rect 7555 -5072 10165 -5046
rect 7555 -5301 7715 -5072
rect 10005 -5301 10165 -5072
rect 7555 -5322 10165 -5301
rect 7555 -5356 7940 -5322
rect 7974 -5356 8198 -5322
rect 8232 -5356 8456 -5322
rect 8490 -5356 8714 -5322
rect 8748 -5356 8972 -5322
rect 9006 -5356 9230 -5322
rect 9264 -5356 9488 -5322
rect 9522 -5356 9746 -5322
rect 9780 -5356 10165 -5322
rect 7555 -5430 10165 -5356
rect 7555 -5464 7940 -5430
rect 7974 -5464 8198 -5430
rect 8232 -5464 8456 -5430
rect 8490 -5464 8714 -5430
rect 8748 -5464 8972 -5430
rect 9006 -5464 9230 -5430
rect 9264 -5464 9488 -5430
rect 9522 -5464 9746 -5430
rect 9780 -5464 10165 -5430
rect 7555 -5492 10165 -5464
rect 7555 -5711 7715 -5492
rect 10005 -5711 10165 -5492
rect 7555 -5740 10165 -5711
rect 7555 -5774 7940 -5740
rect 7974 -5774 8198 -5740
rect 8232 -5774 8456 -5740
rect 8490 -5774 8714 -5740
rect 8748 -5774 8972 -5740
rect 9006 -5774 9230 -5740
rect 9264 -5774 9488 -5740
rect 9522 -5774 9746 -5740
rect 9780 -5774 10165 -5740
rect 7555 -5848 10165 -5774
rect 7555 -5882 7940 -5848
rect 7974 -5882 8198 -5848
rect 8232 -5882 8456 -5848
rect 8490 -5882 8714 -5848
rect 8748 -5882 8972 -5848
rect 9006 -5882 9230 -5848
rect 9264 -5882 9488 -5848
rect 9522 -5882 9746 -5848
rect 9780 -5882 10165 -5848
rect 7555 -5902 10165 -5882
rect 7555 -6141 7715 -5902
rect 10005 -6141 10165 -5902
rect 7555 -6158 10165 -6141
rect 7555 -6192 7940 -6158
rect 7974 -6192 8198 -6158
rect 8232 -6192 8456 -6158
rect 8490 -6192 8714 -6158
rect 8748 -6192 8972 -6158
rect 9006 -6192 9230 -6158
rect 9264 -6192 9488 -6158
rect 9522 -6192 9746 -6158
rect 9780 -6192 10165 -6158
rect 7555 -6266 10165 -6192
rect 7555 -6300 7940 -6266
rect 7974 -6300 8198 -6266
rect 8232 -6300 8456 -6266
rect 8490 -6300 8714 -6266
rect 8748 -6300 8972 -6266
rect 9006 -6300 9230 -6266
rect 9264 -6300 9488 -6266
rect 9522 -6300 9746 -6266
rect 9780 -6300 10165 -6266
rect 7555 -6332 10165 -6300
rect 7555 -6551 7715 -6332
rect 10005 -6551 10165 -6332
rect 7555 -6576 10165 -6551
rect 7555 -6610 7940 -6576
rect 7974 -6610 8198 -6576
rect 8232 -6610 8456 -6576
rect 8490 -6610 8714 -6576
rect 8748 -6610 8972 -6576
rect 9006 -6610 9230 -6576
rect 9264 -6610 9488 -6576
rect 9522 -6610 9746 -6576
rect 9780 -6610 10165 -6576
rect 7555 -6684 10165 -6610
rect 7555 -6718 7940 -6684
rect 7974 -6718 8198 -6684
rect 8232 -6718 8456 -6684
rect 8490 -6718 8714 -6684
rect 8748 -6718 8972 -6684
rect 9006 -6718 9230 -6684
rect 9264 -6718 9488 -6684
rect 9522 -6718 9746 -6684
rect 9780 -6718 10165 -6684
rect 7555 -6742 10165 -6718
rect 7555 -6971 7715 -6742
rect 10005 -6971 10165 -6742
rect 7555 -6994 10165 -6971
rect 7555 -7028 7940 -6994
rect 7974 -7028 8198 -6994
rect 8232 -7028 8456 -6994
rect 8490 -7028 8714 -6994
rect 8748 -7028 8972 -6994
rect 9006 -7028 9230 -6994
rect 9264 -7028 9488 -6994
rect 9522 -7028 9746 -6994
rect 9780 -7028 10165 -6994
rect 7555 -7102 10165 -7028
rect 7555 -7136 7940 -7102
rect 7974 -7136 8198 -7102
rect 8232 -7136 8456 -7102
rect 8490 -7136 8714 -7102
rect 8748 -7136 8972 -7102
rect 9006 -7136 9230 -7102
rect 9264 -7136 9488 -7102
rect 9522 -7136 9746 -7102
rect 9780 -7136 10165 -7102
rect 7555 -7162 10165 -7136
rect 7555 -7381 7715 -7162
rect 10005 -7381 10165 -7162
rect 7555 -7412 10165 -7381
rect 7555 -7446 7940 -7412
rect 7974 -7446 8198 -7412
rect 8232 -7446 8456 -7412
rect 8490 -7446 8714 -7412
rect 8748 -7446 8972 -7412
rect 9006 -7446 9230 -7412
rect 9264 -7446 9488 -7412
rect 9522 -7446 9746 -7412
rect 9780 -7446 10165 -7412
rect 7555 -7520 10165 -7446
rect 7555 -7554 7940 -7520
rect 7974 -7554 8198 -7520
rect 8232 -7554 8456 -7520
rect 8490 -7554 8714 -7520
rect 8748 -7554 8972 -7520
rect 9006 -7554 9230 -7520
rect 9264 -7554 9488 -7520
rect 9522 -7554 9746 -7520
rect 9780 -7554 10165 -7520
rect 7555 -7572 10165 -7554
rect 7555 -7802 7715 -7572
rect 10005 -7802 10165 -7572
rect 7555 -7830 10165 -7802
rect 7555 -7864 7940 -7830
rect 7974 -7864 8198 -7830
rect 8232 -7864 8456 -7830
rect 8490 -7864 8714 -7830
rect 8748 -7864 8972 -7830
rect 9006 -7864 9230 -7830
rect 9264 -7864 9488 -7830
rect 9522 -7864 9746 -7830
rect 9780 -7864 10165 -7830
rect 7555 -7932 10165 -7864
rect 10218 -5011 12828 -4972
rect 10218 -5045 10603 -5011
rect 10637 -5045 10861 -5011
rect 10895 -5045 11119 -5011
rect 11153 -5045 11377 -5011
rect 11411 -5045 11635 -5011
rect 11669 -5045 11893 -5011
rect 11927 -5045 12151 -5011
rect 12185 -5045 12409 -5011
rect 12443 -5045 12828 -5011
rect 10218 -5071 12828 -5045
rect 10218 -5300 10378 -5071
rect 12668 -5300 12828 -5071
rect 10218 -5321 12828 -5300
rect 10218 -5355 10603 -5321
rect 10637 -5355 10861 -5321
rect 10895 -5355 11119 -5321
rect 11153 -5355 11377 -5321
rect 11411 -5355 11635 -5321
rect 11669 -5355 11893 -5321
rect 11927 -5355 12151 -5321
rect 12185 -5355 12409 -5321
rect 12443 -5355 12828 -5321
rect 10218 -5429 12828 -5355
rect 10218 -5463 10603 -5429
rect 10637 -5463 10861 -5429
rect 10895 -5463 11119 -5429
rect 11153 -5463 11377 -5429
rect 11411 -5463 11635 -5429
rect 11669 -5463 11893 -5429
rect 11927 -5463 12151 -5429
rect 12185 -5463 12409 -5429
rect 12443 -5463 12828 -5429
rect 10218 -5491 12828 -5463
rect 10218 -5710 10378 -5491
rect 12668 -5710 12828 -5491
rect 10218 -5739 12828 -5710
rect 10218 -5773 10603 -5739
rect 10637 -5773 10861 -5739
rect 10895 -5773 11119 -5739
rect 11153 -5773 11377 -5739
rect 11411 -5773 11635 -5739
rect 11669 -5773 11893 -5739
rect 11927 -5773 12151 -5739
rect 12185 -5773 12409 -5739
rect 12443 -5773 12828 -5739
rect 10218 -5847 12828 -5773
rect 10218 -5881 10603 -5847
rect 10637 -5881 10861 -5847
rect 10895 -5881 11119 -5847
rect 11153 -5881 11377 -5847
rect 11411 -5881 11635 -5847
rect 11669 -5881 11893 -5847
rect 11927 -5881 12151 -5847
rect 12185 -5881 12409 -5847
rect 12443 -5881 12828 -5847
rect 10218 -5901 12828 -5881
rect 10218 -6140 10378 -5901
rect 12668 -6140 12828 -5901
rect 10218 -6157 12828 -6140
rect 10218 -6191 10603 -6157
rect 10637 -6191 10861 -6157
rect 10895 -6191 11119 -6157
rect 11153 -6191 11377 -6157
rect 11411 -6191 11635 -6157
rect 11669 -6191 11893 -6157
rect 11927 -6191 12151 -6157
rect 12185 -6191 12409 -6157
rect 12443 -6191 12828 -6157
rect 10218 -6265 12828 -6191
rect 10218 -6299 10603 -6265
rect 10637 -6299 10861 -6265
rect 10895 -6299 11119 -6265
rect 11153 -6299 11377 -6265
rect 11411 -6299 11635 -6265
rect 11669 -6299 11893 -6265
rect 11927 -6299 12151 -6265
rect 12185 -6299 12409 -6265
rect 12443 -6299 12828 -6265
rect 10218 -6331 12828 -6299
rect 10218 -6550 10378 -6331
rect 12668 -6550 12828 -6331
rect 10218 -6575 12828 -6550
rect 10218 -6609 10603 -6575
rect 10637 -6609 10861 -6575
rect 10895 -6609 11119 -6575
rect 11153 -6609 11377 -6575
rect 11411 -6609 11635 -6575
rect 11669 -6609 11893 -6575
rect 11927 -6609 12151 -6575
rect 12185 -6609 12409 -6575
rect 12443 -6609 12828 -6575
rect 10218 -6683 12828 -6609
rect 10218 -6717 10603 -6683
rect 10637 -6717 10861 -6683
rect 10895 -6717 11119 -6683
rect 11153 -6717 11377 -6683
rect 11411 -6717 11635 -6683
rect 11669 -6717 11893 -6683
rect 11927 -6717 12151 -6683
rect 12185 -6717 12409 -6683
rect 12443 -6717 12828 -6683
rect 10218 -6741 12828 -6717
rect 10218 -6970 10378 -6741
rect 12668 -6970 12828 -6741
rect 10218 -6993 12828 -6970
rect 10218 -7027 10603 -6993
rect 10637 -7027 10861 -6993
rect 10895 -7027 11119 -6993
rect 11153 -7027 11377 -6993
rect 11411 -7027 11635 -6993
rect 11669 -7027 11893 -6993
rect 11927 -7027 12151 -6993
rect 12185 -7027 12409 -6993
rect 12443 -7027 12828 -6993
rect 10218 -7101 12828 -7027
rect 10218 -7135 10603 -7101
rect 10637 -7135 10861 -7101
rect 10895 -7135 11119 -7101
rect 11153 -7135 11377 -7101
rect 11411 -7135 11635 -7101
rect 11669 -7135 11893 -7101
rect 11927 -7135 12151 -7101
rect 12185 -7135 12409 -7101
rect 12443 -7135 12828 -7101
rect 10218 -7161 12828 -7135
rect 10218 -7380 10378 -7161
rect 12668 -7380 12828 -7161
rect 10218 -7411 12828 -7380
rect 10218 -7445 10603 -7411
rect 10637 -7445 10861 -7411
rect 10895 -7445 11119 -7411
rect 11153 -7445 11377 -7411
rect 11411 -7445 11635 -7411
rect 11669 -7445 11893 -7411
rect 11927 -7445 12151 -7411
rect 12185 -7445 12409 -7411
rect 12443 -7445 12828 -7411
rect 10218 -7519 12828 -7445
rect 10218 -7553 10603 -7519
rect 10637 -7553 10861 -7519
rect 10895 -7553 11119 -7519
rect 11153 -7553 11377 -7519
rect 11411 -7553 11635 -7519
rect 11669 -7553 11893 -7519
rect 11927 -7553 12151 -7519
rect 12185 -7553 12409 -7519
rect 12443 -7553 12828 -7519
rect 10218 -7571 12828 -7553
rect 10218 -7801 10378 -7571
rect 12668 -7801 12828 -7571
rect 10218 -7829 12828 -7801
rect 10218 -7863 10603 -7829
rect 10637 -7863 10861 -7829
rect 10895 -7863 11119 -7829
rect 11153 -7863 11377 -7829
rect 11411 -7863 11635 -7829
rect 11669 -7863 11893 -7829
rect 11927 -7863 12151 -7829
rect 12185 -7863 12409 -7829
rect 12443 -7863 12828 -7829
rect 10218 -7931 12828 -7863
rect 13150 -6860 13526 -6848
rect 13150 -7094 13230 -6860
rect 13454 -7094 13526 -6860
rect 6135 -8172 6245 -7932
rect 6135 -8198 6165 -8172
rect 6134 -8212 6165 -8198
rect 6215 -8212 6245 -8172
rect 6134 -8481 6245 -8212
rect 6134 -8517 6166 -8481
rect 6206 -8517 6245 -8481
rect 6134 -8536 6245 -8517
rect 8805 -8172 8915 -7932
rect 8805 -8212 8835 -8172
rect 8885 -8212 8915 -8172
rect 8805 -8478 8915 -8212
rect 8805 -8521 8836 -8478
rect 8880 -8521 8915 -8478
rect 8805 -8536 8915 -8521
rect 11468 -8171 11578 -7931
rect 11468 -8211 11498 -8171
rect 11548 -8211 11578 -8171
rect 11468 -8477 11578 -8211
rect 11468 -8519 11498 -8477
rect 11542 -8519 11578 -8477
rect 11468 -8543 11578 -8519
rect 5970 -8608 6124 -8587
rect 5970 -8702 6000 -8608
rect 6092 -8702 6124 -8608
rect 5970 -8714 6124 -8702
rect 8644 -8608 8791 -8592
rect 8644 -8702 8670 -8608
rect 8762 -8702 8791 -8608
rect 8644 -8715 8791 -8702
rect 11312 -8608 11459 -8594
rect 11312 -8702 11336 -8608
rect 11428 -8702 11459 -8608
rect 11312 -8717 11459 -8702
rect 4014 -8978 4518 -8856
rect 13150 -8978 13526 -7094
rect 4014 -9240 4114 -8978
rect 4408 -9080 13526 -8978
rect 4408 -9240 13524 -9080
rect 4014 -9284 13524 -9240
rect 4014 -9390 4518 -9284
rect 3861 -9641 3900 -9635
rect 244 -9675 3900 -9641
rect 13862 -9591 13903 8655
rect 13938 8539 17447 8655
rect 13938 7163 14018 8539
rect 14052 7163 15676 8539
rect 15710 7163 17334 8539
rect 17368 7163 17447 8539
rect 13938 7029 17447 7163
rect 13938 5653 14018 7029
rect 14052 5653 15676 7029
rect 15710 5653 17334 7029
rect 17368 5653 17447 7029
rect 13938 5519 17447 5653
rect 13938 4143 14018 5519
rect 14052 4143 15676 5519
rect 15710 4143 17334 5519
rect 17368 4143 17447 5519
rect 13938 4009 17447 4143
rect 13938 2633 14018 4009
rect 14052 2782 15676 4009
rect 15710 2782 17334 4009
rect 14052 2633 15200 2782
rect 16200 2633 17334 2782
rect 17368 2633 17447 4009
rect 13938 2499 15200 2633
rect 16200 2499 17447 2633
rect 13938 1123 14018 2499
rect 14052 2186 15200 2499
rect 16200 2186 17334 2499
rect 14052 1123 15676 2186
rect 15710 1123 17334 2186
rect 17368 1123 17447 2499
rect 13938 989 17447 1123
rect 13938 -387 14018 989
rect 14052 -387 15676 989
rect 15710 -387 17334 989
rect 17368 -387 17447 989
rect 13938 -521 17447 -387
rect 13938 -1897 14018 -521
rect 14052 -1897 15676 -521
rect 15710 -1897 17334 -521
rect 17368 -1897 17447 -521
rect 13938 -2031 17447 -1897
rect 13938 -3407 14018 -2031
rect 14052 -3407 15676 -2031
rect 15710 -3407 17334 -2031
rect 17368 -3407 17447 -2031
rect 13938 -3541 17447 -3407
rect 13938 -4917 14018 -3541
rect 14052 -4917 15676 -3541
rect 15710 -4917 17334 -3541
rect 17368 -4917 17447 -3541
rect 13938 -5051 17447 -4917
rect 13938 -6427 14018 -5051
rect 14052 -6427 15676 -5051
rect 15710 -6427 17334 -5051
rect 17368 -6427 17447 -5051
rect 13938 -6561 17447 -6427
rect 13938 -7937 14018 -6561
rect 14052 -7937 15676 -6561
rect 15710 -7937 17334 -6561
rect 17368 -7937 17447 -6561
rect 13938 -8071 17447 -7937
rect 13938 -9447 14018 -8071
rect 14052 -9447 15676 -8071
rect 15710 -9447 17334 -8071
rect 17368 -9447 17447 -8071
rect 13938 -9591 17447 -9447
rect 17482 -9591 17519 8655
rect 13862 -9636 13902 -9591
rect 17487 -9636 17519 -9591
rect 13862 -9671 17519 -9636
<< via1 >>
rect 1441 2706 2055 3196
rect 2055 2706 2089 3196
rect 2089 2706 2738 3196
rect 5925 8323 5988 8484
rect 6051 8324 6131 8483
rect 6202 8324 6282 8483
rect 6314 8325 6394 8484
rect 8924 8291 10483 8517
rect 10369 8289 10482 8291
rect 5030 7516 5269 7519
rect 5030 7214 5064 7516
rect 5064 7214 5237 7516
rect 5237 7214 5269 7516
rect 5030 7206 5269 7214
rect 4070 5342 4316 5560
rect 12461 7503 12683 7504
rect 12461 7184 12464 7503
rect 12464 7184 12679 7503
rect 12679 7184 12683 7503
rect 12461 7183 12683 7184
rect 13352 6744 13514 6920
rect 13352 5818 13514 5994
rect 5998 2906 6104 3012
rect 8662 2906 8768 3012
rect 11324 2906 11430 3012
rect 5019 1648 5202 1953
rect 13352 1936 13514 2112
rect 4098 938 4260 1114
rect 13352 1010 13514 1186
rect 4098 12 4260 188
rect 5992 -2813 6098 -2707
rect 8668 -2806 8760 -2712
rect 11334 -2806 11426 -2712
rect 12270 -3719 12275 -3405
rect 12275 -3719 12477 -3405
rect 12477 -3719 12486 -3405
rect 12270 -3722 12486 -3719
rect 4098 -4044 4260 -3868
rect 12915 -3646 12986 -3574
rect 4991 -3950 5147 -3946
rect 4991 -4214 4998 -3950
rect 4998 -4214 5141 -3950
rect 5141 -4214 5147 -3950
rect 4991 -4218 5147 -4214
rect 4098 -4892 4260 -4716
rect 12551 -4315 12607 -4242
rect 12940 -4315 12943 -4242
rect 12943 -4315 12989 -4242
rect 12989 -4315 12996 -4242
rect 13192 -4860 13442 -4570
rect 13442 -4860 13444 -4570
rect 13192 -4866 13444 -4860
rect 13230 -7094 13454 -6860
rect 6000 -8702 6092 -8608
rect 8670 -8702 8762 -8608
rect 11336 -8702 11428 -8608
rect 4114 -9240 4408 -8978
rect 15200 2633 15676 2782
rect 15676 2633 15710 2782
rect 15710 2633 16200 2782
rect 15200 2499 16200 2633
rect 15200 2186 15676 2499
rect 15676 2186 15710 2499
rect 15710 2186 16200 2499
<< metal2 >>
rect 8856 8544 10450 8546
rect 8856 8517 13552 8544
rect 4110 8484 6417 8511
rect 4110 8323 5925 8484
rect 5988 8483 6314 8484
rect 5988 8324 6051 8483
rect 6131 8324 6202 8483
rect 6282 8325 6314 8483
rect 6394 8325 6417 8484
rect 6282 8324 6417 8325
rect 5988 8323 6417 8324
rect 4110 8286 6417 8323
rect 8856 8291 8924 8517
rect 10483 8291 13552 8517
rect 8856 8289 10369 8291
rect 10482 8289 13552 8291
rect 8856 8267 13552 8289
rect 8856 8266 10450 8267
rect 5012 7519 5290 7538
rect 5012 7206 5030 7519
rect 5269 7206 5290 7519
rect 5012 7187 5290 7206
rect 12426 7517 12727 7528
rect 12426 7167 12440 7517
rect 12713 7167 12727 7517
rect 12426 7157 12727 7167
rect 13320 6920 13550 6962
rect 13320 6744 13352 6920
rect 13514 6744 13550 6920
rect 13320 5994 13550 6744
rect 13320 5818 13352 5994
rect 13514 5818 13550 5994
rect 13320 5802 13550 5818
rect 4014 5560 4406 5616
rect 4014 5342 4070 5560
rect 4316 5342 4406 5560
rect 4014 4848 4406 5342
rect 4014 4624 4104 4848
rect 4352 4624 4406 4848
rect 4014 4586 4406 4624
rect 1218 3253 3130 3434
rect 1218 2612 1420 3253
rect 2932 2612 3130 3253
rect 5978 3012 6122 3020
rect 5978 2906 5998 3012
rect 6104 2906 6122 3012
rect 5978 2896 6122 2906
rect 8644 3012 8788 3020
rect 8644 2906 8662 3012
rect 8768 2906 8788 3012
rect 8644 2896 8788 2906
rect 11305 3012 11451 3020
rect 11305 2906 11324 3012
rect 11430 2906 11451 3012
rect 11305 2895 11451 2906
rect 1218 2401 3130 2612
rect 14888 2811 16695 3008
rect 13320 2112 13550 2154
rect 4979 1953 5257 1967
rect 4979 1648 5019 1953
rect 5202 1648 5257 1953
rect 4979 1616 5257 1648
rect 13320 1936 13352 2112
rect 13514 1936 13550 2112
rect 13320 1186 13550 1936
rect 14888 2109 15147 2811
rect 16349 2109 16695 2811
rect 14888 1859 16695 2109
rect 4066 1114 4296 1156
rect 4066 938 4098 1114
rect 4260 938 4296 1114
rect 13320 1010 13352 1186
rect 13514 1010 13550 1186
rect 13320 994 13550 1010
rect 4066 188 4296 938
rect 4066 12 4098 188
rect 4260 12 4296 188
rect 4066 -4 4296 12
rect 5970 -2707 6124 -2697
rect 5970 -2813 5992 -2707
rect 6098 -2813 6124 -2707
rect 5970 -2824 6124 -2813
rect 8654 -2712 8779 -2696
rect 8654 -2806 8668 -2712
rect 8760 -2806 8779 -2712
rect 8654 -2818 8779 -2806
rect 11318 -2712 11443 -2692
rect 11318 -2806 11334 -2712
rect 11426 -2806 11443 -2712
rect 11318 -2818 11443 -2806
rect 12223 -3389 12539 -3369
rect 12223 -3738 12258 -3389
rect 12504 -3738 12539 -3389
rect 12879 -3555 13023 -3541
rect 12879 -3666 12898 -3555
rect 13002 -3666 13023 -3555
rect 12879 -3680 13023 -3666
rect 12223 -3749 12539 -3738
rect 4068 -3868 4296 -3826
rect 4068 -4044 4098 -3868
rect 4260 -4044 4296 -3868
rect 4068 -4716 4296 -4044
rect 4960 -3946 5193 -3926
rect 4960 -3956 4991 -3946
rect 5147 -3956 5193 -3946
rect 4960 -4212 4980 -3956
rect 5161 -4212 5193 -3956
rect 4960 -4218 4991 -4212
rect 5147 -4218 5193 -4212
rect 4960 -4251 5193 -4218
rect 12528 -4226 12631 -4216
rect 12528 -4330 12538 -4226
rect 12617 -4330 12631 -4226
rect 12528 -4342 12631 -4330
rect 12915 -4227 13018 -4214
rect 12915 -4330 12928 -4227
rect 13002 -4330 13018 -4227
rect 12915 -4340 13018 -4330
rect 4068 -4892 4098 -4716
rect 4260 -4892 4296 -4716
rect 4068 -4908 4296 -4892
rect 13150 -4570 13526 -4520
rect 13150 -4866 13192 -4570
rect 13444 -4866 13526 -4570
rect 13150 -6860 13526 -4866
rect 13150 -7094 13230 -6860
rect 13454 -7094 13526 -6860
rect 13150 -7126 13526 -7094
rect 5970 -8608 6124 -8587
rect 5970 -8702 6000 -8608
rect 6092 -8702 6124 -8608
rect 5970 -8714 6124 -8702
rect 8644 -8608 8791 -8592
rect 8644 -8702 8670 -8608
rect 8762 -8702 8791 -8608
rect 8644 -8715 8791 -8702
rect 11312 -8608 11459 -8594
rect 11312 -8702 11336 -8608
rect 11428 -8702 11459 -8608
rect 11312 -8717 11459 -8702
rect 4014 -8978 4526 -8860
rect 4014 -9240 4114 -8978
rect 4408 -9240 4526 -8978
rect 4014 -9400 4526 -9240
<< via2 >>
rect 5030 7206 5269 7519
rect 12440 7504 12713 7517
rect 12440 7183 12461 7504
rect 12461 7183 12683 7504
rect 12683 7183 12713 7504
rect 12440 7167 12713 7183
rect 4104 4624 4352 4848
rect 1420 3196 2932 3253
rect 1420 2706 1441 3196
rect 1441 2706 2738 3196
rect 2738 2706 2932 3196
rect 1420 2612 2932 2706
rect 5998 2906 6104 3012
rect 8662 2906 8768 3012
rect 11324 2906 11430 3012
rect 5019 1648 5202 1953
rect 15147 2782 16349 2811
rect 15147 2186 15200 2782
rect 15200 2186 16200 2782
rect 16200 2186 16349 2782
rect 15147 2109 16349 2186
rect 5992 -2813 6098 -2707
rect 8668 -2806 8760 -2712
rect 11334 -2806 11426 -2712
rect 12258 -3405 12504 -3389
rect 12258 -3722 12270 -3405
rect 12270 -3722 12486 -3405
rect 12486 -3722 12504 -3405
rect 12258 -3738 12504 -3722
rect 12898 -3574 13002 -3555
rect 12898 -3646 12915 -3574
rect 12915 -3646 12986 -3574
rect 12986 -3646 13002 -3574
rect 12898 -3666 13002 -3646
rect 4980 -4212 4991 -3956
rect 4991 -4212 5147 -3956
rect 5147 -4212 5161 -3956
rect 12538 -4242 12617 -4226
rect 12538 -4315 12551 -4242
rect 12551 -4315 12607 -4242
rect 12607 -4315 12617 -4242
rect 12538 -4330 12617 -4315
rect 12928 -4242 13002 -4227
rect 12928 -4315 12940 -4242
rect 12940 -4315 12996 -4242
rect 12996 -4315 13002 -4242
rect 12928 -4330 13002 -4315
rect 6000 -8702 6092 -8608
rect 8670 -8702 8762 -8608
rect 11336 -8702 11428 -8608
rect 4114 -9240 4408 -8978
<< metal3 >>
rect 5012 7519 5290 7538
rect 5012 7206 5030 7519
rect 5269 7206 5290 7519
rect 5012 7187 5290 7206
rect 12422 7517 12728 7532
rect 12422 7167 12440 7517
rect 12713 7167 12728 7517
rect 12422 7155 12728 7167
rect 4014 4848 4528 4926
rect 4014 4624 4104 4848
rect 4352 4624 4528 4848
rect 1218 3404 3138 3430
rect 1218 2431 1265 3404
rect 3065 2431 3138 3404
rect 4014 -8978 4528 4624
rect 5978 3012 6122 3020
rect 5978 2906 5998 3012
rect 6104 2906 6122 3012
rect 5978 2896 6122 2906
rect 8644 3012 8788 3020
rect 8644 2906 8662 3012
rect 8768 2906 8788 3012
rect 8644 2896 8788 2906
rect 11305 3012 11451 3020
rect 11305 2906 11324 3012
rect 11430 2906 11451 3012
rect 11305 2895 11451 2906
rect 14917 2868 16661 2969
rect 14917 2075 15027 2868
rect 16426 2075 16661 2868
rect 4979 1953 5257 1967
rect 4979 1648 5019 1953
rect 5202 1648 5257 1953
rect 14917 1926 16661 2075
rect 4979 1616 5257 1648
rect 5970 -2707 6124 -2697
rect 5970 -2813 5992 -2707
rect 6098 -2813 6124 -2707
rect 5970 -2824 6124 -2813
rect 8654 -2712 8779 -2696
rect 8654 -2806 8668 -2712
rect 8760 -2806 8779 -2712
rect 8654 -2818 8779 -2806
rect 11318 -2712 11443 -2692
rect 11318 -2806 11334 -2712
rect 11426 -2806 11443 -2712
rect 11318 -2818 11443 -2806
rect 12219 -3389 12548 -3365
rect 12219 -3738 12258 -3389
rect 12504 -3738 12548 -3389
rect 12879 -3555 13023 -3541
rect 12879 -3666 12898 -3555
rect 13002 -3666 13023 -3555
rect 12879 -3680 13023 -3666
rect 12219 -3758 12548 -3738
rect 4950 -3956 5194 -3925
rect 4950 -4212 4980 -3956
rect 5161 -4212 5194 -3956
rect 4950 -4251 5194 -4212
rect 12526 -4226 12627 -4217
rect 12526 -4330 12538 -4226
rect 12617 -4330 12627 -4226
rect 12526 -4340 12627 -4330
rect 12914 -4227 13016 -4214
rect 12914 -4330 12928 -4227
rect 13002 -4330 13016 -4227
rect 12914 -4342 13016 -4330
rect 5970 -8608 6124 -8587
rect 5970 -8702 6000 -8608
rect 6092 -8702 6124 -8608
rect 5970 -8714 6124 -8702
rect 8644 -8608 8791 -8592
rect 8644 -8702 8670 -8608
rect 8762 -8702 8791 -8608
rect 8644 -8715 8791 -8702
rect 11312 -8608 11459 -8594
rect 11312 -8702 11336 -8608
rect 11428 -8702 11459 -8608
rect 11312 -8717 11459 -8702
rect 4014 -9240 4114 -8978
rect 4408 -9240 4528 -8978
rect 4014 -9394 4528 -9240
<< via3 >>
rect 5030 7206 5269 7519
rect 12440 7167 12713 7517
rect 1265 3253 3065 3404
rect 1265 2612 1420 3253
rect 1420 2612 2932 3253
rect 2932 2612 3065 3253
rect 1265 2431 3065 2612
rect 5998 2906 6104 3012
rect 8662 2906 8768 3012
rect 11324 2906 11430 3012
rect 15027 2811 16426 2868
rect 15027 2109 15147 2811
rect 15147 2109 16349 2811
rect 16349 2109 16426 2811
rect 15027 2075 16426 2109
rect 5019 1648 5202 1953
rect 5992 -2813 6098 -2707
rect 8668 -2806 8760 -2712
rect 11334 -2806 11426 -2712
rect 12258 -3738 12504 -3389
rect 12898 -3666 13002 -3555
rect 4980 -4212 5161 -3956
rect 12538 -4330 12617 -4226
rect 12928 -4330 13002 -4227
rect 6000 -8702 6092 -8608
rect 8670 -8702 8762 -8608
rect 11336 -8702 11428 -8608
<< metal4 >>
rect 5012 7519 5290 7538
rect 5012 7206 5030 7519
rect 5269 7206 5290 7519
rect 5012 7187 5290 7206
rect 12422 7517 12728 7532
rect 12422 7167 12440 7517
rect 12713 7167 12728 7517
rect 12422 7155 12728 7167
rect 1201 3404 6152 3443
rect 1201 2431 1265 3404
rect 3065 3064 6152 3404
rect 3065 3033 6480 3064
rect 11163 3033 16820 3037
rect 3065 3012 16820 3033
rect 3065 2906 5998 3012
rect 6104 2906 8662 3012
rect 8768 2906 11324 3012
rect 11430 2906 16820 3012
rect 3065 2868 16820 2906
rect 3065 2846 15027 2868
rect 3065 2840 6480 2846
rect 3065 2431 6152 2840
rect 8644 2621 8788 2846
rect 1201 2298 6152 2431
rect 1201 2293 6157 2298
rect 4963 1953 5287 1983
rect 4963 1648 5019 1953
rect 5255 1648 5287 1953
rect 4963 1623 5287 1648
rect 4979 1616 5257 1623
rect 5970 1133 6157 2293
rect 8639 1153 8793 2621
rect 11163 2075 15027 2846
rect 16426 2075 16820 2868
rect 11163 1995 16820 2075
rect 11165 1806 16820 1995
rect 11165 1722 12273 1806
rect 11165 1157 12171 1722
rect 5970 -2679 6124 1133
rect 8644 -2679 8788 1153
rect 11313 -1197 11457 1157
rect 11313 -1445 11458 -1197
rect 11313 -2679 11457 -1445
rect 5904 -2707 11459 -2679
rect 5904 -2813 5992 -2707
rect 6098 -2712 11459 -2707
rect 6098 -2806 8668 -2712
rect 8760 -2806 11334 -2712
rect 11426 -2806 11459 -2712
rect 6098 -2813 11459 -2806
rect 5904 -2866 11459 -2813
rect 4941 -3956 5239 -3923
rect 4941 -3959 4980 -3956
rect 5161 -3959 5239 -3956
rect 4941 -4233 4975 -3959
rect 5211 -4233 5239 -3959
rect 4941 -4263 5239 -4233
rect 5970 -8571 6124 -2866
rect 8644 -8571 8788 -2866
rect 11313 -4214 11457 -2866
rect 12219 -3385 12548 -3365
rect 12219 -3743 12248 -3385
rect 12512 -3743 12548 -3385
rect 12219 -3758 12548 -3743
rect 11313 -4226 13023 -4214
rect 11313 -4330 12538 -4226
rect 12617 -4227 13023 -4226
rect 12617 -4330 12928 -4227
rect 13002 -4330 13023 -4227
rect 11313 -4347 13023 -4330
rect 11313 -8571 11457 -4347
rect 5916 -8608 11471 -8571
rect 5916 -8702 6000 -8608
rect 6092 -8702 8670 -8608
rect 8762 -8702 11336 -8608
rect 11428 -8702 11471 -8608
rect 5916 -8758 11471 -8702
rect 5970 -8760 6124 -8758
<< via4 >>
rect 5030 7206 5269 7519
rect 12440 7167 12713 7517
rect 5019 1648 5202 1953
rect 5202 1648 5255 1953
rect 4975 -4212 4980 -3959
rect 4980 -4212 5161 -3959
rect 5161 -4212 5211 -3959
rect 4975 -4233 5211 -4212
rect 12248 -3389 12512 -3385
rect 12248 -3738 12258 -3389
rect 12258 -3738 12504 -3389
rect 12504 -3738 12512 -3389
rect 12248 -3743 12512 -3738
rect 12874 -3555 13111 -3451
rect 12874 -3666 12898 -3555
rect 12898 -3666 13002 -3555
rect 13002 -3666 13111 -3555
rect 12874 -3689 13111 -3666
<< metal5 >>
rect 4971 7519 5338 7554
rect 4971 7206 5030 7519
rect 5269 7206 5338 7519
rect 4971 1974 5338 7206
rect 4966 1953 5338 1974
rect 12388 7517 12788 7562
rect 12388 7167 12440 7517
rect 12713 7167 12788 7517
rect 12388 5118 12788 7167
rect 12388 4798 14256 5118
rect 12388 1962 12788 4798
rect 4966 1648 5019 1953
rect 5255 1648 5338 1953
rect 4966 1646 5338 1648
rect 4966 -3136 5340 1646
rect 12236 1547 12788 1962
rect 4769 -3138 5348 -3136
rect 12236 -3138 12786 1547
rect 4769 -3208 12786 -3138
rect 4769 -3385 13426 -3208
rect 4769 -3743 12248 -3385
rect 12512 -3451 13426 -3385
rect 12512 -3689 12874 -3451
rect 13111 -3689 13426 -3451
rect 12512 -3743 13426 -3689
rect 4769 -3817 13426 -3743
rect 4769 -3818 12786 -3817
rect 4769 -3825 12541 -3818
rect 13106 -3819 13426 -3817
rect 4769 -3924 5348 -3825
rect 4766 -3952 5348 -3924
rect 4766 -3959 5341 -3952
rect 4766 -4233 4975 -3959
rect 5211 -4233 5341 -3959
rect 4766 -4345 5341 -4233
rect 4966 -4346 5340 -4345
<< labels >>
flabel metal4 13704 2468 13704 2468 0 FreeSans 1600 0 0 0 GND
flabel metal5 13726 4948 13726 4948 0 FreeSans 1600 0 0 0 VDD
flabel metal2 13406 8408 13406 8408 0 FreeSans 1600 0 0 0 Vinit
flabel metal2 4254 8400 4254 8400 0 FreeSans 1600 0 0 0 Vctrl
flabel metal1 13592 -4022 13592 -4022 0 FreeSans 1600 0 0 0 FvcoBUF
flabel metal1 13012 -4654 13012 -4654 0 FreeSans 1600 0 0 0 Fvco
flabel locali 7474 6756 7474 6756 0 FreeSans 1600 0 0 0 Vso1
flabel locali 10392 6756 10392 6756 0 FreeSans 1600 0 0 0 Vso2
flabel locali 12174 6762 12174 6762 0 FreeSans 1600 0 0 0 Vso3
flabel locali 6972 -4850 6972 -4850 0 FreeSans 1600 0 0 0 Vso7
flabel locali 10092 -4862 10092 -4862 0 FreeSans 1600 0 0 0 Vso8
flabel locali 8644 9054 8644 9054 0 FreeSans 1600 0 0 0 Vst
flabel locali 10726 1058 10726 1058 0 FreeSans 1600 0 0 0 Vso4
flabel locali 8194 1032 8194 1032 0 FreeSans 1600 0 0 0 Vso5
flabel locali 5608 1072 5608 1072 0 FreeSans 1600 0 0 0 Vso6
<< end >>
